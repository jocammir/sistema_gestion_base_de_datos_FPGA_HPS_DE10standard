��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�(H��$���x�`�4V��_.]�-!�`D��I��L)]��姛��V:z�e�۹�I��+*Ny�Kk��H%��% �A
�k���������������=J����u����Ā���d>�g+��M˳وdM��R�
��=�kd�[Y#&���0���cм?a��m������d�h�����Ϳ�*�x�����3r��rOogi#+��)�*�&dC`��r�tȠ��英mT�St��)�=��	��i����=�GMI��5�?��55g<�7�����9� ɳ��.��Z�8���
�O�J�<�K1^���M�o?�x�zBb���Vݗ�J]�n>���F�xi�`5lXFpF��Z�L�	�����yV�Tg�oM�\�� �^6V>�:�h����L�h�hYu�F����Py8�m���$_��Z�W��	b� ��L�����#f�n'���	�=Z�S+�ї o�����h&F~�$@HD�Y�rӉD���Hu�G:���� 'ǜ���9`Y�� p�:��u��,\�1G"����a稨�4�s��6��M{W|�1�'�b�:�^v����2�#|ЪQ��|C��L擄-��|M��H�����d s�r��L�w���8b���`�FU��>��wӣs�')u�h#YTYNAz�M=�e��6�7o������/�������_M\�1')������a˲
7�p��巻��8�2�ѥw�����2�!G�(�~hv�N��6���Z/��+7���T��b�Q�S�����s��A��6
���q^E&2ۆH�ͼ��
��/C��ɲh��uW"R�<�5}]<��ҥ�{�n�9ځ���:��I�^[|8�K�7��|�g��r�/8����¼��\k��a�&\f�vѳ�����\���Ae�5{l��	^r��4��rpe46 �n�<�~�huP�Z�(GR�oKJ����BX�gJ�xӈ�7���60fBܗ�<u�8�sC��*ے�ΠrF�V��E�����3)�rgfp���ʋ�d��>�+so�1�%�vk�5m^�Y%r�'d�A�>��>��]�H�X��5"$~��?�\a>�,��/ʯ��!�P�1��ZH1�"������/ ��C؀���F�:�Lߗ�L�x�	+�WxQu��<��H:���v��{'z��ߜ��,3m$5B��`Q�.�D�uN4��F��=�f]��U�F���}e�5/Ʊ��4���[BGy��aFG�����f����9 �t!n2�V>��MO�.���] �J�8L��}�K��/޸�E_��	&[����n(��^���&��a�5�l��s&I��3��@�H��%�?J�U�hl�W�K��β&W�P�\w,�d��s*��)�	���wI��d��C!��%�l�[�WF&X�+Z��:�È��,�7>�|�8��$Z�O�KWč�cA��׭u����)���zCH�-ʺ�����yS&�H�[�5�OX�h�}ݗӓ��1A�G�dy�l���d0`fwo:�}zYTT���0<%�=r��kJ���Y� �N�K�ۗt��:� ���%B3�,����g��}�����h���@v�S]��@���8j0��~��m�$�L���B4��j�DK]YHp���$<ߐpJs��K���&�
=e����;�(2���/����KT����H�ⷔUB�u恿hU�b2lbD���M����Y}i�A�t]+|��s
`UƷ[������k� !�|���ү�P'��Rէ�[\y&���q�����Ȕ+�S�H�^�ts����|#�����1�J��������旱zu�@��=N!�f������H�3����5��{�s��f�>����UB�\ӝ�V)�B��Hi~�-�J��&׋�47��%R ���)�%f�`�h�th�+�':-��N.>A=;�LR�|���om��/WST�̫�=/��6�9�1R�����$��cIt{�M�舾�x��Ბ�!0<��R��uY��������3p&�� W~�i��FH\����s��󜃈�w�P�A)�"e��0	6� ���s0$W��� ��n��V/*#���O���Q'�Z�������Ә>/!}�2^��L=�E '�s�)��2���Mg���<t��k����Gv�۲������d��ø��>� ���j�6��Y��m@}�Dш��rޕ�YlUh�Dlܳ�$�i���lKP��0��Qr`�����p��Ҡƽ#�ܩu~瑙7*�9�"�ƒX ��E�-�\�qU����$H��x��j�E���?��5DdڬX�6�6�t��J�k�����W�79V��a�x��h��z�s��mZ�#�U��>t��#��O|��ʸ�C�:��N���S���-����z��:��ƥ*"-aJ0��6�]��58�߹˩�s�L��=��/E&]�H�,���a��H����;�i;��S����D)ǃyKc>&�p�C���>w��5qRS��7W�J��nN�2A@���V$��e�Փ���!<U���[3-<�c�s iq[���Q�s��k..d-J]��uQ4���0���ah�L>����b`��ˤN�����̯�U��;kڣ��l��0<�;�S�F�����[`��pI�G�_k� ~��mv=Y��ɥ\�l}���(5&.��8J	�d-���M#�S$��Գ���9�*'3&P�a�zZu�u�g߀�d��(6�����Ŧ���M%?B�ǆF��بk�4I�L�=ݶ�R�=��dZ�SW7�M�aUc�e��-"�V/�k��fmk��J$�3�q��r�b�Fv���1>H������Nb���Z��aax!�e����H��D���>�+H�h�ޮ�Yl���?�3B*��`"b�Oߞ�I��{���Q�����J�8�2��{_I$pXAW��bCKQ�?����#g�%?�y�'�F?O�n�&]�|e���fL�1�m/\1<��
xW>硃!RB�@�F�K�Q{�_��8ƙή�G?IW^Ǭ��S�p����B#�9� r��
��6�_�W�y&̽�9|��)�����trr7�v�`���MA���k����-f�@��:	������&W�$@��L�XQ�ǡُD+���d����ۉU��f!zǮU:bF�Br���,?���R�X�|[%�)5i��4�j
*Wa�UՖ�������Y{$̙}�Y�������	�>QO�c�*���F*�~��*���%Mȋ��0���TPq�DQ�u����O�e=v�F���MTW2��=���IZ�U׼F�	�G$Mfi�y�#��j)c�G��'���7f.�B�z�GZB����?U-���:�'1+���z��fq�Y�"�C�T�.y W��۴��YT�X	}9�w�IbD\_�_m���>�y�Y��������s�{��}0�f>OpΝ`O�7�6<v��h������sԢ�O��@ L��F�:	*g)7 �fC�i+U#�|.�#����l� ��+%����%Z����&����>�1X�X9~��*��*�NυN��e��D���@Ѯ#%�1׿J�_ d�V�f��"��y+��EQ���|���f�u�����q�$����+#��yA��eʻdę/����]L#��~QPS+].*c���r���W�7BI��j6��t�P
�l�v�UOF!S���*>ز\L����LU��ñiSNt8p��W��h鮻Jh|z'4'$oZ��}hj�lv�����mb�Ǘ��Pb�xó��p�5mc�-O�}�i��~��㥴C���'��ǹ�4��k�����d���a�	|ku�c�τR>�?~�j���~�|�L饮��=����'bs�s�����DV���A/�g^Q��	zd�9���]VHUó�	�s�p@��K�1U �A@R�-R��@|���t���xY܌]�i��?�Jō�O��Z�pC(�5��7F�f[�x�����U�\B#6J������8S��ˌ��Jq�w@ۋp��C�=u;��8k��Pj��dO��сC�Q��B�(�hp���i���#yˍ�Mǎ�3O��m��8�u�N�SG_�K'�6>�H�vV�KT�#�oi2�}	���V�_�nL���kH	D͠ݣ�$��Ӊ���FXE�R&�3��[�Tf�Ԅ��9^Y�I��<q��A].�3(�o���6%]��Ȗ�B��Gv�-�o�
�) ��J 44�����_�e�.Ɠ6J��d�_+�.��E���rx��n^�z��{ݨ�O�yG8�38j]#@rY�rC�
@Lm�%�F=X�;1g�%j�,�/6�0�Ν/�r&��k���&��	�O@��ev)~M-�W{�i�z<ꇩ�*�OX�Dғ[Ry��]Z��8��|q媹����:˨*&b�s���+$�(��ჟ��l�xS���ݵ��ߣ�<��>�՝D��'4���@u�X��d�]ZQߠQ�.Z��ᤕ��)@�"<�g�R]}�3�J��$���v���ܮG�c������E@��R��Ɓ�B�w	���{�$3��e�,�Wԇ��NV�e�����Bl���M�Dc����ߥ&�@�6
\D�lt ���e��y$H5���{~T�=���?�t=���L�3��W"���tLr<���������wI�^az5��it>?�?n�(%�����'���^@wW�-�+���H���bJp\ͤ�SQ��ת�B��P�F�/�I{ɿʭQpΨ�a87�N�ͦu����mp�w�f��!,|����Ma�ZM�_ ~�t���	��m�iG,#(�/���w�r��@{�<�~��=vY���+�
R%H��ԜK�g���
L4���A@_VI���
�m�Ə�ݛ���%��8�C�pN1OI�\M8��Z��uYS2���{��R
̌()
�^!���>��'�qΡ�6x�Ĳ���3�>�=�:I̜�7 [�_DE
nJ���K�G�Ź��g2̼{�Y����PDAJ(��'�Z?iu�2����.<����9���N3��8?��$��ne,ΫO3?7h���C���!	 txG3���n��A�R	9[��K1�w�)��F��UW#B�1F�g���+�rR:I�u���=Fs/�����")��#�@�	r:yʎNB���oq��׷%�EUeyRA�U��*j��6�n���P�h�z����\x����ƚ�T}��A]�gSI/�hL��7r�g$��V6a���9�����>��־ᰆ�Λ6�F4B��Tb�+h�Q�B%$#���	�wYy�x�I!��2$V#0����������q��|�
s���ن4:�X��1�:�:t{��e2��0�n#���g��ٿ3҇���6E�.���yC�1��=G���^İ�gy�*`�HC�mԢKG���,P17�ɯ�F�Gʱ�f*.���`^�08:!�[�r+a��/��9D�)������@�$_�c��O�r�1�?��ǫ�0|����Z->F���E���w2�.�.�I{���.����>��,�gg�m�J]=jt�ɔ��Oy��J���zEэ�Ȩ�%G!�TN����b^�?Ox�z�:�6��%��� ����ͥ�m�o�T,b�GW~x;?�k�<�Pq�v�9q��B�!�	Q>�^
��+�_�0�Q�L���D`��궏���Hv#taj)mvsg	%a��RF�����Ջ$���6�@�NU�%?�����o� ��2 �C������C,a�g?��S�5��*ճ��������3τ#.�*S�F�ܨ3�DB�e�ܢ��E2~��dy�%��9�gU-��V�Y�q�l�����D>���@�������8름q��@g�k0�3tg��9
W-��X�']��j��b&�*$���J�Hf��v��w�K��/�����|��RXB�%4