��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0���
����wC��s�;B��h�o��1@i�M��9.�y��mu��d�ZaV�=xˉ?�fǯ(u����l���*ƛ�շ6D�J��5�#�:v��IIN�w��'���=�\��ZA?A1#�hq)foP�lM���S%����g8���
^�?���&��ßw��9����eB���`u�Pn�x�����p<������8����Q��+)D;5h)��	�r�%��f���W�kf�!U����?��xu��[kc Q-��%bW����Y �9_�ªg�oR���ns����F��Ip�s*f�����M|�c�]2Z�%!
�Ixz�������0He�E��d�㌂O�D���}T�;1��"]���cjφ�4_h=.Yo�c�Y��]��+�-����+SCH����7u�@�CZ��_/z�lm 
�!h�7h������2�K����U��{���0�@���dR�g$ҦR��x��|pZ&0>q�eG��]�b�\�>�����L_V��^ُ�fԊG�6��{PKa2�&@S��dl_�i�aU�%>M!V�4yn_7q�M}���&4n�ĉ�m�}���6;���X�������|�I�3t(3��T����s��Tn�o6�R�vO��X���u� �))�j����:��H����<G혬}�����L��B�ĥp�G5�~�CO����Հd���n�.J�3��~?۵V/��
W�:���~�7�('8����8�%��?�w ����c5{�W��ݹ�5\�& �S��t��
NÒe,B��JJ�L��雳�%?6J���S�$��^�'��"O5l�^�Av���
�mg0�'�!�k��}��E1l�:!j7�rt#9�l���+V ?x���n%b��l�e:zg���V�����������VP�U��3qrh���B�&-aPr�����y���)�N��ܷ�@�YR8��vk��/\>ΰ�#��g�w��?2���*�kU��FI�K���N��nY�ɟJ��X7� 6j�ߝ�jO.0�q�s����g��h��G�}R|E��-����Yb�͆/�t�H�:��:���X��6�9N�B΅�B�X
��_�c�7P��	�bya�\p�xJnU�e���������qKUz{5�ל�Չ���9��S��p$QMK޶୓A�=R��ѤDf�=�uSL��-�3ȡ�\n
W���Q�d{��)+P�G��@	�C�D��G4�cx��K���|�ײ\)�FFZ�3��ӌ,F��U0թٵZu�OM563�-�պe��Wsɸ�B#Z�y�иC��'a�ˤ�V ͡NK�U��Z<�2�}T���r(Ŏ��c	c��U"\N��N�Ya+�:�V�߄��y�/��Y��T�`N)�v�k�O����ߦ;��#���0¤�s���3���Q�/�m;k�ۙ^Gvy��G������o�_�#�*p������'`Ď�c�_PU�m��;O�����@�墖|�g��t�
(����Vh�"�q���6���_y5��H���x֣��U+�5�ve"� ��B&ش�p�8���fs-`rߖ �������>�k�wU�ן���J�D���@e`{��vAp�[�~�!&D,��>�A�dͦ+���4�՚�O�� ����]��ߵ�1�S�J���]u�L�[�O̭w�aX�[��o�t�&3�-����.����(��!�QC7�ݎ���^�&W7�]�t`%�po��]�XTˢ��<*�% A�LgtH��O$���*]yy�
�M嗙2���E��_3��Sl���`�ҍYP�:�#&x�Ӛ��+�#X��\��)�ĄS�]؃1��������K�^��ޖ����V�5��T��`� �}�'�/�G�����6�����WH��6��䉀�Xq|�d�LU��$�W�'_��Dkc7�[��x�v����S�=��`C4f>�9�L!��r�b�
�#?a�O�$(�0��T3�^�^�W�%�~������.]y9�pT��*���:�? �l�T�X���r<�&j}��;my���]��qߐ*5��8����w�u��=`�d�{��*0a��50rnP���t�Q��l0�h�ׂ&��mP/����-nZ0ǟ�w����3ue���	2�YtG�Ģ��"GB�k�-Kq�����S$����j.������3Uu�lJ��bB��<�����3Ǚ	�;�f&A#��?!m�r�u�sO��� �72�ҷ���G�i���L�P���-��0�j���M|�*W���5�KB���Gv}$B�J$[�Èo����VW�LRM9X�����m,\�]����B�&N�Y��������#
�a���@cc	t5����q�?ZN/��4.r3^	�+���(���qg�䖝H�h�C����z�8h&�^��\�76��� L�N=L�FxKl���_ ��j���Vԡ������ee�H��:e�fn�K�)*�-f�_��v5�U�e�Eޘ*����2Iv0��7��e�DJ�%n��v� PI0oJƹ�zQ%ʫ]ԣN,g�i�\\i1ʁo�L��\H�)�$�Y�#oAss)�)�8������N_���.�j�n3W�" x=���٢��-䵈u���M�55x(�� uR���!�4�8O��j����'� uB[w���;ů�����M����_���R�����Y���4@T�R���s6%XH
�C3���NU �.U9�(���>�[���t!#M���+~^mB�_b5t]t�A�B��$BJ@m��~�G������D��ϝ��D�xYj���G`�?`��%��ym
�=���]��#i��b�QY� ǅ]�T+[�R���]���K�@� �i��! y8hvV��vߩ�n3w}����<a�������|�@���T�Uhْ�\�rQ)�DS��nJ��̚|d*����/ⷣ�����U���'�����Q��ȧ�к�3�yU)�ƾR"��)S}w�V��{]l{5I���Ư�d���N����[��y��� ��w�v ��>�����o����H���O�mm4^�}�O��-A"���Q�n�>�茋r%? W���ӸQ��fT
��Ml��l1�f1�&�h��7��5���ͯ�f*�^�O/��Hd.���{]���A��&�t*�����'s����$u�Ґ;�i���s�́��T�6ܝ������5U�AmD!y:M��s�7�E���VY��Nԅ��j�l튋谍��y���0�t�/vh<̠͡A�$�hǘ��v��k�_�V�^"��Z���gŋ����_���ҳc�OM��L��N��$�:��?e�߆3��*�o�Z������o�(Y����*H�qY�K�|AN��Q�K��Q���C�+��j!�&����c`)a}���d$:���k�a��E��oQ=�֋���
$�!u�::T�|�a��Ko��w�28�) ��(TI��$!�J�@/���E&!�<����O3��
�"Nb��NwJq �}�i�N�ٻj)/���%�c�c^oi2Sz�*�r�y�D�t
؀)n�Z�֑����-�,W2Y(�WO���r�m=�mX�=�A�`F�#^�NWM�7Ⴊ��K�ѧ$+x�&�Ũ��䔟ixm �(i��u�����ۥ�F��(f���@b-@hs�ƅ�������A��`n�� H'M�2���|A�r�UE���+�wʨ�y�1w�?=N�����i�BՕ.�tp��w�h�[%0�x���C[}�bX�y?}�U~a+V�!9o�]\2,ٶ��I��pFh���Gc�:��p	(OIZv�P���C���1�t���s�wTBty�!!՘F$)�<���N �rq�R��^��kq	���Ҫ�D��������b<����Da����m