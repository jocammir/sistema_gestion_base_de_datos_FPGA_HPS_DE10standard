��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0���C	�i��EM'XGi���ozmo��L@��i�ʉ�f�wkmrsuڟ�6A3��ؐ����#�#ߺ��,�^#�+M3��a����?�@���jK�£�_��"kbN�J�/� q�h!�Fm� �,+���)�~��$o����.t�C�Y�C�Q��7�8�p2s�쵿�׎�㏨=����ҵD.����O"�p� @Z�0��ļ"H�H��ӽ���rm�O�L�A��u)���F���'�ý=4��X3�:��
I7�tȱ�%�7���aV��J�)b�piy�gT�f_@�G�rAR��7B���X�Y"^�#�S�Uw�ר`�s�P���U�;e�����Sd�ݾŖi��9)�f97$���t���j���?4�!�7�rM��>����+�>�B y|.iq�L�j�P\� )�w̌���lr�p����fK �p��9-�M,F�ܲҖRb��a/K���R/].��_R�{e����8�?;�9����-�<ꪉA^��1��6�4��p�e歋T-��`����c$ΈR��"�O�y�}����O���%�	���]d��x.Hf��)AǪ��r�ύ����]mF�����<��ֶ�_����E)��q�}��`1�&/g͖��h&I�-E;Ф��'��y��:$���B��{/М*�z$��{�xu��SU���j�����f� ����x��6�b�S{$�#J�Ƅ�WS�&���K�ٻ[\�YB��K��;����s��]1X���>�N�8��� Ry��1�;�� �D��#�����[H���S�Qp�q;�Q�E�D�[����5��m���]�1-����p�o&��)�=�$K�eY��:�#ld=�ށ�^��$������y�\2����i<Yc�L#�a�ߟ��C��#��JqR7�aSp�>�R8AC�/v��ze�<з���P���G�����P�e�Q��+����2�E+�6Ih�Y��Fs`�Yar�*�.��L�bu����>�<@�3t�����L�`�\oq\��I'��	��h��(9#��YOs0�:�u,�k��&q��66d�8�{��?��%����_�V?; �$ȇ}F����h��ex���ם����rl(��i���E48�?k�N�G����<d��|���ņ��ڬ+{�>�������(R���5�$R]Yn*,ǊD0�A��u+D`p�JtiY�Jĥ�'�ώ鲯y��Y���Gƙ��t��ќ�.���_�?��A<�z�`��* 9�&E��7i�#��%��ǧ~��i΁t?}`mu�Y�s�B%���~��**����e @!�&��N;�
��]@�ߛ���Q^��R8[Sf+��s��w�A��?<?Y��H��Ԉ������cn�g/i��_U�	\}%�� ��o��vP��w͇�<Z\�%�U\,[��5��	��>�[��P������ ��{�6u�����܃%)1C⥍/$rAT$&Ұ[�y���%�{�>əcU�b��\e(�Y�<5�q��.�Y�@u�~V@�����3��<�֟ ��qx����J��E���.��R��j+>̿T�v�*�<2�s�Q"��1Dš4v�f�kg�G4:HU�v+-�CꄢqǼ�����+lT����nZ�h�E�Z0����/�a�?��q�h	�t���6\.�y(j4�3�����)=�!%�ퟦ��/4��{��[˽5�F�.�:���5]������_u��V��p�0��Y�x�@ZO�>�v��[�6إY��7۬�E�Z��Q��3y�N��+Q)O�5�O�&�gb�
�Wef'wE0�"���"�ͽۆ��R�p��BV.y�d��ܶ��r�̺4����ऌ}-p��qpM$��2�Gdo�_7Zs��D��Q^3�y͛vv1ו�VK�m6Y %��p7R�n��=^(�-u�w���wi�dM� ������ �D},˸�:��S�3��J{'�"{s*�y��<aZ���ۇ��?�z��l�fQt�����Gׅ�s>�eG{C��}�{2����ei}I���o��{��ny���}���	�og��+p�Y�:���Mrn=���E�IS��77�"����>z�psG�[M��ͯ��U�QXZ&������V)��-��,c!�������lg�v����y����Ї�U��4B�o��� �˔�93��x�C��