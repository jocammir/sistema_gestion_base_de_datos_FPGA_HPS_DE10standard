��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0���C	�i��E�>>�S=��}�,���o3u���F�[L	��\�d,�(N҄,������6�C��z�(���!����]�A��N>�R8��b��ꗕ��Q |���J�����E�E���!ZR�k%�{t��@��L$�>x� :K�P
��~/�4.��P������Ӎ�2R'�l�K)��&�c_f	U��bM��a߉U4w�J������oE�i�k����+�|=�C�)z��W� e��uJ��td��Bq�����fq։f��}���m�?�Y�p<(�7��A�����XҮ䉋�zp����v���^,��U�\Q߽� /���6���z�ހ��i�aTB��&�<��_�����/��rس��[И�e(�ɂ����ue��@zBV}ɩv�� ��+���
�yG��;�jrl���5�kh�´v|�� �k�`xgׇ�i����O��	�#��b]r8@��P�
��f��C�5��vfG��n���5�&��N��I�'?��NVߚ�Ѻ��,�k3��2tfV�{F�u"�� �☛=k8��^��h�v>IX�+_�!�t�+-���G.�h0�� L��%t��
Een�2z,_�M�t��?a��O���5q�rO�LM,��nL7z[�C�y���!)s�~���B�m�29��6n֢\�2W;��G�ڛvxFp2?c<*M�T���"�Rn��@Ɩܵ��)�����[�Y��?Ү���;�K�R���,���`%�'����Xh���ø� �Hɇ�4W�{LM�C�O�@HV_��P�[�r�di V�yq��R-�݆&V<215�+�r-)��lS���������nntj8��]��~��YVu�_�}�+p�"�1���G��D<�]�C��S�I�>��P��(NN�ߨ|pѬ�9ש|�\�t
9ˍU\���m�fSa$�Z�DX7�L;|\�{ �+A*
C����nš�Td5
&��o�hLnД�ơ�(�F���]�}�<ׄ;6��n�������<��9G��m{�l;.�%���eT<rf���C�1�0s�2�a{N-X��xK-fbi���gD�>��[ ��&�j	*�`gF,>J�Z�a�E���.h����J�_o�����E��Ƕ��Ի�]j���&|4!�h#�PU4g��Fm,I�
���+c��C{�v��&������[4