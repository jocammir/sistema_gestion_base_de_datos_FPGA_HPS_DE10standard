��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0���o���*)?]�<��gA���4���5N���W�w
�cfF�sP��@|����礙���Sʼ��F"Z��/�n!���͐'��"wnq�~1��,��m"t5'Y�_�����w��!��Vz^��S�#P��P_@�M4-P����B��Y���HdSW��%���`��E�J�"$�����ɋ���	���H�9���5��m`e&�F�N0�/�T��9�a�R�~򸂘V�p�T��xw#��s@n�h�l�4��_�*���sw9�����M*[]'HԮ��M0��Н�ô��Y�_�E�gnP��B�J�s�پu�r0���)`�25ki��#�֠I�a��_�-�����\)b�l�F�Pc�M��l:.c���������dP��@� �(+����m��[�0=�}����v-\<�K=}Ǆ�t�3��ς�L��^�x�f��N�f� Σ[��0��8I�UR�!I�u�_��CImk{�����3�It�uW��N�1�_������U�����'c��x��R���i;FW�K���?�Sj����]����>����@��y�I4�;?9�}j��v�%���Ez��1�h���t�vhU�:���z�n�A�/S�;C�%��+�@�B���؇Li�Bx= ����
���;#�b�k�Y4�U�Q����T�17�����F�O��GC#]ҼK�#�hXPڮ�i��Ҷ�N�F}1ɴ��L.l�W:3����.�9�|0r�X�hz��q&��@�03�"H8C�Ӧ# � �9`� S�1Z��5+�Eo��8*�ן�L�E㶎' �������H�:I-ZLW�Ҹu��\Ԯ�rM��j�j�Kd�@��-�o[�H�B���l�Z��� ��,��[�v�u�Ӄ	r�kӎ@�/�l���}�y'w2���{�r�g�p����ye(<�eC/J��0�0.�PX5Y�ۤC�r�X�� ��Dyʼ������cu�FZ�������_�k�V"�zXX�=Qp��W,y~��.�����ŋT��F`�tx�oـ��@�����Y�������-��(������9������b��5 ��j��$"1�,ѓx�U�@1s�M=���@3o� 4�wnM ��b}�$tL�ɦ�D5
v~��EO ��Qg h�����2�����+�d,67ADo*ɿM�8Xz	N�XIޣ��<,�7P���~�׈�ۉE���-.�Pcl��d ��x.l��Z��<)���EP�.|x��W��l"K�70v-����a��j��D:8"8��������ګE�]�&��hﺢ~�nz]����,Û���D���u��m�~�7�����F5�"�BWx��������_�Ψ�^�=?����p�خ����X4j�`��Ϳ��>�n�:M�b�[���rN+Lk��Gȁ��?"t����?�9�t�p4���|Ðc�k�P˙�Bcs�R������O
��Fnq��ş;�6^*��7| �[�.�<G 4�pl5H$1�LÊ��+8�leZ!4H�.y8zJw[D�h>�]$`'Y���T,x�壯s�[=�-�ٻ������ݜB!�2��3ֿ,����
,�Bѷ5d��DIxj�艁�l�������-�n���6[{�$MĮ�nz�/bRǕ<�p�����q�e�d�.u,s�����r�'�6�Z�q&�H��4��!���/�J��Nqif�VS[d����!�������ߨ>�)O`����⇫5cj�ڈ����o��/%����
�C��Z|U�/��
�c�m��Jk����?8���,y��D|��Ë8��Fv*aH���Ө%?܃r����#���b����L(�za�LJ�� ����+����_'ʇ,��va�>�A��N�P?�6���:�`f��S�xs�0��lqt�_%9�C/�0�;�ߖܳ"�]�or6��'��h�֘���M��V�Q[6{O5䢻�3��(�F�;�do.-�T�:��rЭ<+���l���yNFĄ>n{?k+�y	��V�����N{N�*>���v�~���i�q\Hr�Vs�!J����~E�����78���ı�!�'(�#'߸:�i#� �����f�ufZ/��[oO�N&����pp�ŖxZ٘��ud���}�y�@�	��[n�fۍ��pf�ـ�vʹ|<Y
��q��,������|�`r���I�)�)dK.���K�����	��������a������JΨ��G�����.V����1��	���<A�,��D��L�$k�_ه��bO�W�(%��6��E���	؇����$�
nE�Z���,R���`xš�ty��iP�ARqI^Z��ra6be����惘N�eD���r��� ��ļa��GC"�r�<Ω�k���7�o�s~̽;T��I��]�ԏ@�Z����6�P��m�����P�&�s��!Ƙ���!�AB�J] ��^*�>���XA�K���&��%��f��$>6��w�WgM�x�fl��X"�_�sr�,5N��F���{ǣ!	��s"�S8�x���f!W�LYԫ�A����v��/t��(4�=Ι�Jo��.����*�ZC�N�.��R����4�/�����NM�T'7xݑ/͜����V��Ow�<���-me'���N[I�2��y��'{뉍���qPS�e��vQ�n��/�Ӣ�N�s�>��e���M�'��̣a��X�X��ɓn�nӘX���3HYB����U��EL��F-:���ĕ���L;`��΋�ٝ�ZNξgwwt���!L޵����|CSyH��Ԑd_ �����$#������o�_���%;�"�Ϻ+=T}r���s/�����9�|��"��ٚ+
̛x��:�r1�q�r�1}����T��s�l墹���`-��Ѿ;����з	s=/��ҔJ�;�M��� #����X�eXE�:���6���c�ob��N���e����
y���z�ݙ#��\n�C��ix��!�Y�F6��z:6[�����$�8�iecf`<�}?���\`�I�C;�[	G�Y� �h�{­��6^��_��/kY��/��F�8�2���Џ��*�;����;W�%t���tSFRVGɅK,����ȁ�����w���w<�� )��_5S�T�������y��Eu4(Bx�B�"�0y�D�J[��@r�f-��iu�0eǭW�핅3��E��
��$���0��scM�
�TYO"O��C�@F��'��x�]�����p]�ǭ��I�*�ݜĆ��}ʒ՜�ݎ�
��b{����: n^NXFv�0�~誗6� R	Y�� ����b~��*�$�?�OО�$�f}	6	�[�G8|�(T��Qr�<	V��mk��ٟɬq�$ɥ%Qj�<�g|���)�,��߻�����Q{�!�7��Q��Ҽ>{��^o�5�A�l{t�Y���P"g ׮d�A#z�r�����+�;���^(�d�����2�������x82���	y,����XRBr�f�7O�����p����=}� �s��6m����`7?�	 aA�un�c"m&�`�PFQ&[@�`b����-���Wԏ���!���a�.P��d�88��"��/=.�}F
g�������!^y*ﵨ�_^��7��Y���T�����YU���2Tf����%j��$�&�շk�4�w�=C^���g`���d��5�RhT@�Q03���F�y�*�x���4J��:"ȄA@Q�z|���=m�p3��ʺ��=BB�_������[E6Z�<?Q'��C���9ȸ%��+��0ɳ���KJf�����Y>��PM��� H2XT���V�H�p+O�R����w˧'������+���4������"��3A�OII�%˪�����%â�z�C�x�
Rk�zsH���a��i���@ɿ����C=%�餠��_Uv;IU�0"�����`2G)��9�g�[	�
'i�	\�����k��?��ӷ5��Zlw6L���?�\u��
����h6$Z��Ǌdkx�Kzy���#���>(:r~���*X4I#�ڲ��|,��f��E$��Ns�x���M�7��]�Hs8W��2�YW��L5����f����'��2�k�p7|�>��=h.t�~ ��輎��Lc�\���kK0וө���!�NȺ�m�@Ȕzt�o��o�cO��?x;�-=:��jN����t`��@I�@��;��AK�T�c��2��e���nN<����P�A���꜔c��qp-��_�L�1@��6M������4��7�1�i���#��ӓm���&N�R �l/@<ch_׮GhѼ�d�����~��d�k���:u��{�/�%��n0�#�(ZI3��r|�����F�V�a ��P�OH��HPU���_���4|�w�9���.�Z�	R�N�W[Vf����ߋ��}7Mͱu��>�n�iȵIv:/�m'�w��I�M wpx?�32e�;c�Wk�S=�RH�>�=�Տ�O�Δq���t�hI��X���y�^0巵�<���:bq]����T!2f��"��>}�-c�`�
?q��M���1ׁ�	T��@&
����\{O1�s�(��9�l["�q�({��)s��%i���\���zR������I��~�w����񙳁�y�E6ȓ�z�n�U�]�3��`����(�^N���x�Bx��A ���,kŎx�"d=l&��x~vx �	�2�G�^ ��R��m}�ڡO6�)*�W�H:��:�LG��^CŦ�3mON���Xg>!�xM�Ɵ������/z��F��0IR��ݞY.ܮ�iH�sY�%ť�&g"k=������禋eF�q*,��I�?۔�2a�TX�<g��$no��6��IL�)H�M�I�B�W�9f^i��/��鞒\��m����=T̩�#�Q)��g��.�iAE���]�2���oNX;y�l���X�1^�'���<Z/w({�x�I�7Z�=#�� �8޲��w1�����J�+�~��E��\M$��x�k�lC�-,7C��0PR+f��џ�ţ����G�D8f�7np;�ԊN�����w�wyRզf
���{�>Oo�S,:<k}�"���s�s9p�k���ú�ʎ��Y�B`Ld����L�/HBYc`��V��&\��P���<��>Uho�|���+��qv1�L��`���/�<DG�����XD�uDI���Y��%�_s����qMג8,�p�j.t�4�D�j��	"¶ԕ<Y��ݺ9^�[ټkHV�M�y�מJ$��� �}�Ԇ� ְ���*ٍD��-+lե�%�ح��%+�d�����������7�y��Q7�q�u��u���>�P�3�;��Zc/QC*uFS� �o%?�>�Okˀ����H�Y"���O��Ak�\<4�I�߫"_�ǭL��)���ib-^Iac��@8�.�K7�պ4�M�]��I��d�:���A���Lk�-?�W���ᾧ���R��f��ݡEΒ���Tj�trr+O)�3y�Q&��C[ɐ�r��A��n����U��YF��E_ϖ_4�%�<�_L�+��0�ٴ��+a��w=+Q��T(WI�3He6K�:����B�G�<c���S�E��%MQ�I�8.��+k,h�2�*��#��ĭ�G1��C3��9�(HX��[���!1)2�Z:�������'Z�Ԯ&��{5���r-���N�եU�ئ[�ּ�}l�C�Q�}�*c,�0�z�0?�v�f�(����C���e�V�U�A�c�/��<�E"��k��V���8�֕@��P��,�������~��V/┰�t����s(��{W�9�t������c�֊V��]�����2]pb��W8t�n�n�R�(�E��o ���ՏG��0�?�@�QҰ#3�"@�exz�d�a4 �,���Mz�3`��B�fj/L���MP�H�l	��F�\8IѴ	������h���&L#h^ca*�3�K%	��!S�p*�͡%R1^-��1ó|��;ga?9�ⱌO�ߦk9r�K����^^�9t���>�������w��S��\
O��6���� z<W�s��æ��+�6�����!��8��D�㢹@����V�m�T����'ڋ+�
�{(�������vo�:�7�~��;�
kP��d��zp��	3�5���i=e�Λ�d�a�$
>�ki|@m\����A�IU�����[�����J>�<���1��)�l�&��c�b���e�y�=v��M ���I�=��g4�u��v{4�._��PSyq+ @�&�Œ�˳�E��/�y����	�J�'�I䭓�Ν��S�6��cAY�	�hSE����a}���;y��ιB�v X���z��g�(�t� TÆf-��-<�c�fm��(h��hi��J�2
�k�2�@Ƈ�� ��U��0w�� !�۪�'Fv�;Qni��!j�VQ{%�_�6���Dn���N��q�l�O0��	�;�џ����j`&�Un{7O0!ĕtf���%��,C+ �*r�ܮ��ao�v$��Q3��0�3�l�������9�Ԏl�B�İl\ǋ��`pm�C36j�
�L#����	�r{����ӄΎW���G�>�twJ�W�.Mק!���׿�i��y����n�iEc[�;1k-�k7��(�D��	�7���4~A>T��������Lal(q'�������֏��W$xƈZZ4GU�Ѭ��;� �c%���Se�� U�Z�t*KLfJJ���Ԅ��20i��f���ϥ�;���{�'fuH�S.X��`'�%@���Ȧ�[-���:v9�7��:�3򎷞<�>�wI�)��_WQ�	Fm�����AL�I���y�2!��S�:2Ԧ�g3B�tE`�ݞ�d�^��~m��Rٷ���n�+�Z�XfP�$�X�F݁丫��E0���� :���6����ǥϺ]������>��0'{@���Ѵ�+�j��Im�evH�x
e8w�^qv�ׇ�Ʃ�w�	���7d���؃��-X�0�n~����*�_q@����N�ڿ�J�����_
�ۥ���،����:�C�a��+N��r >������������7B��b�E�%�o�M9�x���v^��}ma��Q^ۨ��O�!y�?D��t������r��fLPu�����EZ��}0���Y��dX2���T�l�$/�J��D~	��}��۪g�yR�Qy |�/��qKp����E�L��3�N)�oS企=���a�k����.�T\`�,�\O*[F)�>�=��E�J�5�e�jƓ]9�?�t݈��U����5d���=�X�O��s�*Id��r>i�9���<:*���9B����6=G,�L�##��Ȍ^DP�I���M��Ui�Pz�CZ�y^~��1c��oT����鞪�8��I�`���#�_���F]�;K1��Kv�aѬ�̓� �v�7���tێw/)��Fq�;���t� �[Σϭ��5�4���q	tl5�x\�����C�_�Q�H i�dD������Ȕ���*��U�Qz�w�彏]�R��j��̡o�V��ve� 1�\i=ڵ�٬f�mV��1����`�;��F��s�����O�V�V�8��{p�u9���X��ʕu�=��U��*)>{e��P ��^vg?�L,	(��%�E��<{O�z��@�̂YB	����m�њ^�h�.#'�C��/U+j!l����q����t�	�|KK\��]��3�#w&E"�u0#��?b��V���
���/��#��؎_��qC��*'�S�RA���������J�	B�_lk�R��cv�+�'��ۙ�{=��
g?Oɸ�a��$��I$ګ�DA�~ �e�'�Wf4�.�(�l�A@�2��
����/��%�BI�2����Oa�Vs��/�ͬ��%YJ��B�Ki�����?P0Sq���z]�/�p�v	a��pjr��\����M2�t�g6��]�t3X|6�y�,���.Q��)�fg��D�� q�ke���3�q��f�4�i�,�5\�tΒ��;�1 ���%�8m���u]��Nw!�6JRoI�܃�{H4%���5��lh����A����B!e\G�Ԏ����nHP�n�<e���Lj���W>�x��F�u� �۷�Ň{�@�hf��?<�����Q� �&	l������*�׃�&=OK�sу��h��]�/�;3����K`�I	4K~�>O.a`=�k���j��P�ʫ�����Ȋ��u���$�I2i�DF��m!��Y2�Tb�C7�;��ȕ�Ң*"@���ky<�_�Fw�˗�zu����5�r5�=�$N���{�G�q�("�ҡ=�L�/Ǘi��!]����f�~�o��.Wh2T��rJ������I�$�� ��D��y#|�B���3�m� #�9�R��z������$z-Vޤ�]�r!&���&�d����\�T��>p����V!½^I2��Jz��Z�.!T�K�kv��#?C+a��*�G������8wF|s��Z�;?�����,���F4�/`��_��8S�F�G5_4��?X�3 ~$��fH�s����'i4�6�_�zu�5Q�Èr�F������bBbj7�o��'����d~��m3dg�٦B������\�w���������Ǽ���FL]��7[D�E¦@Ɵmd�Q�v���� ��BIӗ�[��(�e�EPR㢁ao�X붸�m�h�����y"�:��7k�\QAOq~���1�.�V�|�>Q� ����qC��1��kr}g#�=,��t�8�Sz}2�X��|�A�T\�� ���dC�G:�A�u}qL���$�	�/&�\?���d��T+ѳ�A���G\�>�!&�Aĕ=��fK�k��I#|!���G�� ��}��b� ��s�Њh�� UE�$��z��t"M�E&��c4��N�\��:Ǹ�xZ���uA�Ze��7S�a͑�EIC��7�h�Μ�6��b�)�0�
�r���oɖQ��eD�	G�P,|��q X�uv��ŖâJF΄����W/d����@7�f#�T�����:d妷�$+ �������P-�i�2��ݯ�l�b��\�}l�k���Ҡ�D��k�>��mc-6���&�lr��2C\�I����G�.#G#�g�šg~�g��dl�l�;��r#���T:8;u���J����=/��b6^zu>�s{J��2����,�7����k�x��lZ�EG���_Hk�]p�l�ͅ\q4�P�|ZT.N�����n
3��8ͳ���TT��{��͹?^�!> L��f�xb#+��	T�����e��$�1�\�j���f�ӈ|m�'���y޿g�X�v��,c�~�^I1Y]?�G�N�~U���eʾ���$��J\�0�D����s�3x-o8���	������CM� �]1s">tϼZEX��q�ؙ��U0b(��-�^)�e����5���@3Ȃv� 4�RkSm�B�i�.S�QpD�T��M�hA����}�@8v~a�����hߗR�J����Z���:��l'FE�0UȔY&�B�
J�r���w����~�oŰ*�h�I@Z~:�x�_��d@���%]/�;<�)���4{�I\c �wLf�҈���z�����iK<���f����0,�غ|�4��e�DC�0�\��-ɣZz��Z�I �C��ca"�(����
����Ef\7��T��Vwx[_�_�|���Y����)K�%o����v��Y��F����e�pF�����GL��r%Fb<t�� ��Ԥ�f��ja�]��擞%���x]>� �ϵG��!�<a��} �h����
Jy�w�&[��~�Ga����Z�_��jl�^[�̶�@Sr�����u�Kz���R󼷚���zR�������3>��e�N=�������Y���l.$k��W�ˠ�;9Q��yZ�C��	Q���z�fs�� ��7z�Grwt?}�`I�uyL����c�ǰ�Qq!�[�`e��6(�}�L@�w���f�/orR��X��d���/�xT�I�J����
��Q�!ȼz|��@�B��~޳�a%0�D	r����z�)*_��bJ����{���h�R�����JEhjE�"�3��7$F.ʢ�?'O��M6u=�Qh`�#��i��o�-��*v�Ү�����ԭJʑ�l=Bw�䥠ɳfd�eH1��bD@l��j\`�A��"�Ad���IK�t�+����N	)	�p�4�f�q6���(�~4�2�5�Ώ��*q_E��q۵�R*I�e!y��=I��'ƞ�_�b}	�L�8�O@�vCZ��'%�/�	���3CN٠�Z��^i�WpʶQ�з�?�PjA��⹂u�����MȞ/��S�]D�~��4���o����[^ t?V��J�����>�Y�b'B�b>|Ө��,������{����1�����Vq/r�R�%�#�~���8K��ylrW��n���䛇�Ә�ۈ�/,�Ӆ�S*�>� �S�T��r_�3og��׵@VT���?;`xx���W�0��0��52qs?��1Wj.��6��~�>
a8��H��;�*�:7�켨ە7�hi��C�*�!�ҌNT�_�H���Y�ba�����U��5���`s�5��Ik�`b�\j˩A��HWj�w0���%����Ç�F�N.�_?�"�?��u��ʍ�u������r����c��h=S�!q 5v��c��v�w����	��8����sC�-���99����>�G��@{P��H��K/W�}ʻ��i�	��&2����xgn���|J��.	:��ԩ��JE��OV�"�r��a�z�ė<����d�^���a3�&vڅ/�s��tP�/�(�2*(�gF^��d=JWKX��.C��y�Y;�ut��k_�
��tYa5�`�T�*��J������]��C�p(4ē�7�-�|2�����u�5-Q��ڲ;0,�'V�8y/u�wa�6�ó�w��Wo���˧y�T]�{Ҫ��㶈�DC�����C�8U���l}�j��k�~+)b��y�p����B�k����^��[Rx�v(�L�Ѳ76�gFM��+l;��EŬL�x<��8�r	�8�w��\(��
m#/ĎP����eڴ�� u�{_�_��NP�d%�OdZpي.T�7��C.LĔ���Y�%zy�p�:_���c�}� �֣��Ҭ �_ �!9hɣ�tNe�+�"�	MN�ۈ���m,�� z3�8)>�T�m�gs12���z8��̉k;dgXn��V1xX��=��{��yt�J�x�%�wwb��׹��=�,Û:�9W�Ưfd׶�t�Ce��E��}8��� �z���"dO�e�/]������� Nh���Xߧ���� B|�}��dy �a$ �X;���"��.�9���-��y��<Q"��	B	����I؛z��M�n���J��o�>���	��#�:�,+������c(Eoq��ړ1z�P@)��`������'2[���MEh�D��U�3�9p�r&�=��n��3mt:���U���p?�?8��W���E��IIE�_פ	v����[�f�Źq�I _\_�727i��K�e,�J?���]��q��fl�M��D���/]iP6���`�w-���X�t?����9�e�rL�n�wg�']�QU���8�r.�>(W-�炬���'�h3oDW��uʋn��s���?p�3 ϱ������;�����!@��a
^���#�O��r�3?�d
� Ɂ�1"��O���2`#�-i4O٫��籽(�S)%"��n헭�	�Iw����cA�B�t;T�%�x~�]��Fy!��ԈcE�xe��U�j6�V�b8�2��������Ѓ���=�%9��[p7��<hR�w`5C���ʬi���t�5	m�U4���cx,?��lH�x��\��?�3�i�cT�/uG����(<a��]�$4�x�B?�ۻ�`-x����>噢T���Ǩ��> �M�I7�BD�_D�RW$J�B~PJ/��(d9}�H16vi��"��J%�0�H6"�n�XM��g�J�<��EK,C3}fi�����E�	�A���0�9������̗��G�-��C� �FG-[�ю1d���39�N#H����Á,=�|���d5����f���ܞ���eŌ�vSEX��Uv"�Ʒ ��*#n��u5�ǵ��@�(j�O���(.t�؆^I������=vBy���zi9>yrkD�l��Sׂ:��[���+G�y�hjnQ]�����EH�P.��W�L\���:�X�YJw����Y����0u	ҎY�1�(�s,����t�6�v=Z �Z3�O5�v},�����4�Ʊ)�6�Ԍ;"?��A��ך��U�%l�P�R!ߧ�˒$���[���~cO�(`����E-ii*���&��gRy��\s�9r����V�2���r@oұZ,�wC��D���~_������`�,,�n�uac�%*�=�{к:1������6���o���{;_XW+�p��ɷØ'����1��c�"���cZ���r۩f�^_ ��(^� h�{��$����f����x.Y�������	�N��0�_��UL�zy<���=���7��Cf����[J�t��jWb��j�%�3�]�䓧����C���M��%����ߩ���DI� v0�����,W��2$�&�c�Z��n�����(ɮ�+xs�;�������`�7nxr�y�z��ڈu���p>Ju�N����(Q���M��q<0:B�ϊׅ#i��n��wHmת��1;,��~y�@�^�fQ�<��i�_�.�M�x��47t]A��Pn��<8}���?Z�CĮ��&%�@ܮ���8����r��RX��zU��i
�<���_K�H|{\w��9E{��6�$���e���5h+nV� �l$��m��\{"�Ab��Y�7 ��I-.C���.��#T�I�����	����3�w!5�g�-,dbx�]P�MMrWAdB�ɀf!��o�pc��Ǯ-��h �a�>fn�:���?Lsg���<�L�R�mpYۿ�[�zӦ���k�
)�-�M��Z1�/|��T�F�f��g���Zt
3�V����O�à%�X�=�^@*;]�XiP���@�W�5 r��D�L��и��H����w�|���<�6�ǻR�Y�В�g����:�E� z1����F�����"^O=�!����B�iX�έ���@FW߷DC<,��m� �� "���_�m2�r�#�E̸�0|����-�+��7'�J4|ҧ۫H=��F̑��F��̂�\�O��I ���3g������ Gf=�۹�f��Y��^�x�y'�Tc��ۉ�nz�y��hTخW�v���A��o��9��sO��zm@����u�����3�DV�ho��J �� ��r�.�l)/:�RT�V�w�ai���M��K���7��qj�E��osʟͿ�-x�;?\�t��.�s~`�H�<qx>�(	5|ԧ�ls�iJP=�Y� �,G���P����l��s�o��k;@~�����<��84J87a{b2z��E
?O� 5iL������L���C=��w].��%��,���H�ǿ�a���#�@Y��e������B*�T�����"N� G�r �v�p+{Is�X���s�W�Y۟�(��?>�n�!�������="��d!��bR;ó ��^@�����L\�؁�δɭ�n1"��c����?u���3z/E�b��#NUl�s�Vc{9+��-Q"�����_�x������!V����4�9�f<�Q�H7X�"�������qX�ӿАn���t�)a�YR|���j��W!%�f��X����FK�B�Lam���0nd�q3v��~���r��hZ��G�@���/e+�˾D�M�]��)AR���6�?�9��lF{U<������?�ϧP�H̊g��p�F��6���ǂ<5�0.�C���}�H��{_u_�zK�86�IX���="���пc�	��8��d� ��d����Fuk�J�ӄ�wn�T��%�,(�-Vm�H��&݌��2���xF���?��V�V���I�O�jh"��-��&�j��&,ҟ���ݸ��??�71��$<+I�N�x��5�$B�Q������v��Q�^��',����H]���m�����H�ig�Ь��'��	$*�N�=�g{��H(����A�'cg^?�fX�߾�>��
�8Q��Y�g��)��0�|:d��@�D%���%�ƿ�tr����9Ev��DQE���4=C6FQ�GJ�ZW�1�!�TA�f��;���ГDO�i�������A��:!��^�0Ի)��R{(\�7�%j�A{�8�hE�z��+tڛ����闚n����� l�(�ؕr��o0����9����=���F`2��,?��$��n>�p_�vG{[V��?���X��*��ֳ9��9��OZ�X�z(��X~�֛��}���֤���3m�J|f���}ɗI�|R<M�1YOwX��&6{v�OS��V�����~���^;��Ѹ|��24����
���[��oW�+�J�3�4��0	�����p8%�+�Վ�|5<Q����g8�a 6|!�/H�o�����xe:8Z0���� ��E�-a��f���o�Xn��6)l'�����f���(F���RBt���1y��T����6k�E�~~�5��D�E�q��nH2D}1���U�n��zB~����f�F�{��@�������A���;9C�sr`�q0�Us�זa暈��n�~����]�0J?��v��97���6�Iv��T2l}���N�.J��w�
���$�ZI�����X)Շ���D[ـ�����0K���ؠ���X�8���j����m值D&�i­�!ySi)x��V�Y���~��wz|���ȅ�n�� �I�/�ʦ�8���WC7;(o�����j$��4X L�[n[3ȹ*��n4���*�Q���u+��
H�H�p��]�_�daj2���`q�L�a�E<���9�*-Y�bwEt�b�L��ka?����#��;�`w�� �u�0Q6��^s���
���p��cH���g��׸_�tऎ+��iyࡰ�-�x��j��c��h�6���K��յ���ؓE4W���-��?�$��.O����HR�p���|�m�%�5"��-�%�%��g�b�e� ��򙷄�'�D���K(�O����I�u��#g���0U��I�7L�&t��˂�@��Ed��jd��0p����>bZ�7qj驜�1kV�,�5}���� �)�d�ߖ	W�-@�Zr�S�}7�k�Q8��%�H�sה!�ܠE�Z�m���@\P�㗣�F�� ��C�1�Pn&#�-yAb������S�Zq?�����.��sLƪ����m�k�Z��]�� T��gD��4;/s��e��1���,|���ȤH�K�U��Sƻ���cќN+*̪�?�\,1�S,
:Ǖ}	��9�%�o�o��"y��}�)=Y��<xx���\'�i�pX�r̀���Y��j��u�"Y�a��0d��[S����	>�
7V|t���kD]2���x��p��V��`)�Y�#���9�o��@9Fl9V���[�{FS9@1N��z���a��
�
��J��sb+�T \�0�9u�3yV�5�U���O����Q@m�3�$Y�E�N+_�>`-��r!�s�17ԚK���������啘A����2�z�)��ЛxG�\�����׎�P��vC��]�Y�/��E�i��%Q{���*�Gr$-�Y�(�gy��f1���P�/B#��$B�ly�O^�zd��*��˲Rѳ�=ƟO#"���=�Z�3�})`[���X��4��iL�/oM��!oE]�<6S����]� m�,vW��R
~f����t���!4������+����.I�cƦw8�w.[��hQ����Mu�"�t�+s���s��<��9;�V?��(���i#NWX��qu�@=;7ϯ�_+EM�8o�'�����Ef���s��K�'w䎈hD�q�Ke��9�2��:�xτ��D�dj2VQ@�thR����Y�u�1{�h.�!_��k��$�7�q�3��&W���TD*��LO��}pu�}��^���4�ӡ&�R�D��U�����(#����NI)>)%� ��;�7��W����5��c�c׷}��~��[���!#$
�;��R)��"�-
�γ��F��?��n�R���+�+��\�;^;�����9{O�h�r� ��J��?)\h� ��^�?��� .�ɶ��ݺ��	v/����NX9�fF��2�����a8��5T�l�K��݈sEW�"2� H5�R"���eǫ1�o�E�P�K��*��s��� )ޓ�ȕzU�ɻ�'[��CT�H
�I�p�^!��>&[�Q#�֧�$������W�q�FAAY������Ƥ��`��uX�4�_�։���ҩ�]q�]���E�֌��JN;���y�6�+�A�^�^[��J��r�l$]͍��;{���x�}ߥ�i�ܐ��jV��V��i$8p%E�u�!�_ 3j0�����\�5��i����+�Nv⤻?�/�W-�B�+�C��%2dsݛ�=���b8�-齇+8,R}~&��I�8�/L����H�	 (��p+�m�M�t�,ѹ@kۉ������@I3`���{W�k˂Tc^��U$�������"�Orä�������f�S?7�\ �@���`�M�:(:/�(�̺"�'e�u��B$ش�_��w4�ZDQ�3e�>���JI�z8kIh�_����k%';��Vl�������\ၩ{������Ug��1����i� sn�t�4A�P��A��I��c���o������3��-��D�vLeǼx �x��(p����D�"�$�媷�Ǌ�N�&�Y�+��� �E�/�N@�ck�71h&�iP`��Ud���%� �y��*�<@0Գ�h,�I����\�;�����"�w�(�n�� �u�Th+\eGO��h�C)���$��V�!}pJ3_�&A�4mbV�޼V�!mn�p5[_�lӿZ��������#lGP�4�o@�0dY'��g>�J��d���݁�?��LZ�o&�\vlVlH��n����6)费2
d�{ɁJ��pđ'�� ���M�?�J^��N�����B�v�b���/��l6���1�#\�C�|`�	�����>BH���}�U��9g|�Ø�Cc�5��	���[_�l
�7��g�P~��S�׳�����-~��lN��F&+�B�S���bSjS�.��Y�|�9��;�v�����$��pY4
�]��'Ci� �~m����z�A�W�ʘ�g����d�W�����rKfB�Ʈ�jw��4Z���+�n�pC�4��3��tKOKe��/�威�3h�Ȕҷ�S۞��EZ�t�G��&����h8�W�:M�C�nfɩ�:��� "y�]{S��%]c*q�T��ϩ���S'�eAw�
�2.����P�p�i�K�=�N� �i���
S�U� �`_Z�+�n�0�3�A���g'+�6�n��"�e�~uCO<�B�>�B����N�$�	;��J�I�VBy{�x�`EG�5"9_L�	�hb8����j��NdN�Zr$+�m϶4��'W�&��L�OI������N*U���_�������$�(�ᇡ���
��_�N��O6)D���`>4��gE�����|p�i�g$.~�aC
�dQ0OS�{%���0��§�JB�s�L��^�,�k��ݮ�Ԭ�pb��Y`iO:ρ�#UZ�߰��?����q��}����q�yl�MG0�8.h_w�vp��#�K"�@�Q)�� [Ӵ�4l�$ �l��c�5CR�J�U�ˁ��5�*�*��
u�*��#�<|&��&j3���T�Vd���Eq�%Zk��U; ���o�}%�4^Mt��nJ^�����#J�id*��ծ3i��`L�~0o�R�7h)|0��6���
��+��j����O�ٞ�y�l�ȓ�>��e�*��=/J�1�>��c��v��f:�(��,��Qȁ��gXB1���Q�Z���~Z��핷rO�>g�
L({����Sh� m3=���J��_c����ʾlA)Iݕx��4Cn@��ď�H��U�ܕ~
�F�p�=�g�_XH�g���_�E���F�)��o�L�����%�'X��w�����	rHR��0�x��Yj�:��Z��>{ޟ�aI���p�_nx�I~��(�9V/���ra_��-�,:�o�K�+>*����k�)�t-	���)���V����1O2�dF�*�k�tp�Xnꎲ���ڊ�Ri��8QaN�"�a�Z��}>h#�<
�A!
Z��+����wȵ/j�*�!̡R�ղ('�6~�q_B�'g��l<��4OًT
$�~���Od3&R���/*}���Ly"����T�3뀎F����Yvf`e��i�	טFp\މ.�6�O��q�Yh�G�D��Ɉn3���\GHWP[���a��ar�>�G0o|�(�i ��V՞ǀh�g�OV�@���G�	V���R��&)"�y��V�8�\Y�<�������
ϙQ�K�b�?U<�b&y�4��y�W�?"�ZtZB��R�i�}b�g\E�_����}N��03��L
��b�1o��zj�Ѱ]͠�9k�<]�b�;q��.ĩ�JI�^�V�Q�Ɂ�O�u�Zu1�Z�0[�|�kZ���^U�
�bd6��%a�I��2zv���Y�H���L!l����Y>�%���Sbچ��(��~0z�������MG;�ϟ���j��t#�U�í`��G�d!��<��Z�� ��0� �y%���M�6�³W\
��;�b���+�A\Cf�V�Ҥ{�)�cV+�2,�.ъ�쒘�1��@���2^�#m�׶ب���N��H{��r�U-k�~��Uʍ�!�&Ez��5�1_k+6�@^������x����w�Xޅ�bO�05[c���R(�.�Mԓ�p��`m��fW���պ+��x�qC� +��!�J6ޛ��|��v����b�7z���`��J�k)��T;�L�k�C,���ps$c�h���,,Z�ݶ귊9�р�ٕ� y��!�R#�Z�&K��͞j���e�;�����Ψ)��\$λc�����ý\�#o��KT�T�d=[<�x40�x�B����-�Js ���0�ݧ��	�Va|��H�7.��T�9tά��%����I_L���*�H�ھ��TO?�w#�O���=Hʔ	GٗS�Q��O ��epf�w��;�z�:ۇ�dKE VE��*ݹ
��O�0�Mf�R�����v�au�1�q'x�1N@��'МUO�r�����7��s��K'e�?rp��&���{��R3�U�w�M��F�u���{�0��u��B�1�m��r�\y3�c`|�^13w��[Vu��؛۹0 ��~�se�q�=V��qs]�5���)t7c�9�Mo*�*eJ��S'z+}b8�V�lK>�O�g�n�#UqJ�/ʿd摖�H�o%3��A�����N\��zJ��"�Գa�J�|~ٲ!9#�����^mJ�ؗ١�=֯@_"g�{3��R$�P�ku|���5¹�T��C�BLE��W���v�D�F���� <׶Z��BS��,���0��3�`�j�=* &����E���*��s�ھ��g��<r3�.Z�6VBk�=��4��(��E6\-��tM�?V�l�,еTw3Q% �[�N�k���"I�!�Kc�])��q88\i@� qm��4m��.��,�۶���SN�uZ&���<V����i�8h����CAo
t����Y���"�����N�ҧ5��v�`l��}<w�ѣ�Y���Ҭ�� ԕαLc�}��tDO�j�p�y1L����!�� ㋞n����=�Q��6z}U&����K��A���^8�g�������2ڝ��tJ�W��5�<���s{�!�bA�� 88�h�������i�����j�F���td��0k���Uyp��T�C����ύ\ae�H�ۺ��,�;x��V��vע6s�@��Ɠ���0|��(e~��\��5[��f��Z�i���LϊoԽ!�z��sj��NP[K#�snk�~�ĘgC�K`��`>�=D�����9˼���}�aq	�t��P+	0V�6R����#�y��(��{oIt
�]3xX��`��E~1X�%=kv�~���%�z�.M|t��*@�O�#:�j[����<�!�����8Y%*Ĕ	R<������A�X �bSxp����y�FzS�y ����i_G-0Z�!>V��sN��h0��0�'p�[gp����!�]O�ŏ}�>�t7�x;CԤ`����W�St�Y�)�ճ+[&5��h�Se%ڪB�~V�Oڲh���H�� tBztb�FP�%C�N��
~�ǯ%{�ӛ�s��,���Y�yr�N�.��
�XL;0jd����&�Exq���C0A3�+�-�g���&и<��M��zs��f�$�vZ@�4���-��ƊQ8���l�|s����>���-�R��t3m#As��͊k�!6ÑoFl��U����`���ٸ��K�ġhb�w��D(9Q�Y�)���0�x�wT��Խ4ԥ�W\��,NA�d�K ��y�d�.:�����Q���%H��(B��G����M�EO�<�4�[��;%گ6��G��/�ab�f�0CV/��s �3�r;3��p���x��E&�k?F��MO���[@r��V�GGn�� i
K����L��Q#�(ۊ�:�E���L�J � 9�/-�UҌ/�)`{T���Z��ԫ�$EjS���U��#��D�硈F@�@���0�p#&E���d��0�Fg�V1t,��"y#��l�9U؀qikr��>�y[!#һ�5˚��#��]unW�Li�����GR���t������%�	>�f
s8}������5������Ҵm��@a���~�QL���̜O�"_93/(]�خO�r����� [4�~�XF����<�"��t�]��m�;��<��5�>�ň*���z�ٱ^UpV��]����S�^�p��H����Ri�쮍u�J�7ٔ_�@�s��ol{4����G����%��$;0:�%?���:�:�mɢp����_�!6u^Uv�)�Nu�?]0�u�LG�c����BgS�� ���C�o�z�*pϣ'7��lW���'���Y��}��V�i�#��6g�M��Wj�\�?��"G�>2��ktL8KǇ(�B+��~�V��xj-����e%+uOb�f��$��nU�>u�.�e�v�h�X�<���	u��P��[��l�C,TK�ʁ�A�S# G%��6W]�� ��C��X4��`B���dn�P�=�!
�@��D�纰��a�n�1�vr�]X�[XyA.�{ɡ��FT�m]f����+l�!Ĥ�}LYiXBS�1kB@�v��\t>�����h)�����y_v�'@OL����o0z1���B�&����2�*�}�p<_���<ُ�ӑ�k0�{�7����j�8�̈́s�f^p��[xV�����1�>�
���KC�0ȃ���}L�d���h)GQՏ�[���\�L.�Qw��lD=�_a�9�[���)�(4b�Kc]6S*�gz�<�M���[Dh��M�w)�v��Y
] �Q�a@l�Mn��RPC�r��
�P���Ы�4x�fq�:�f��H�	s��7�~+�]�ٕ>c��v}��jg�;��i<Q�;ي�=���� ���-�OrUy�I6�R�ΜO42H�G&�ښ��_�a
���[q_]+X6/��=�?�p�1���2���LēmyU�q�Z᫪�@c1�Lbz��c�c�����m�+�I�ql��")�h�}��y�p~�%{��B���W�Q�׃/�ޭ1a.p�w�윘�1Ȧ�%��E�� i�ho�	xͦUrd���Qkd� ]=8�3�3&��B��Z r����R#a��jt0��S�<��"K�o6�k9�\���.����F�"`Z�>p��0êc�K%x��ǣS�l��c����q��!՟;��x�	��Q���������*�MX��:��4�0�G9:Q���m��䰤\f�X�I�vԊV�Zib��<�� 3�qD)YhAW*E�U^�$�����NzUډa�X��UurT�_"ڎ-�t�le�����L'uX��
��n��	l;u��~mH۔ ���5�+HC�qf�g�92�����8��:�5 ����ܛ�[1z} �,���Z�u��%�)u��2��4�+"uvؕb|�5�&��SQ�Z�B7?�z�Y�v>�cr1�M�u�V������d�_���wN3�I�&�ؖ\�d��4�OhZI�ӫ�OU�h⌯8r��Gt��?f��9H^k��J�����WG`�����=���*ͪv���pS��~�Ϝ��&�ƙ[�AH�U��)`2n#�N7<j T��d�׍�xo �c�Q�fv|��C6~�G���k�z�_�=�\�F`�K�4^[JW���ֲ�B��2��-�p6<~�"Q�����|;�/ �Z�a�����j1�x�G�P m4�=����}fX��|�y%�9 ��2��v'Xd{d]��_Rw���\.=8�"��x�B{�z\Ƨ=	C{�}T�7�`&�j��D��$�>3;D�vd~�~-�1���jo���C���+����$K�R ��8��Aj���]��b�+΀xB*��˻R)���Ҹ@�g��6�N������h
!�y��]}�Fr�J�	��VJ�d�i#��2۔��jyُ6Co��h���-�Nrll�� �܈��E�Ո�|?Q3𦕥��>g��e�Z�+dT�}���i˩	��Oܜ�X���=~#v�d���t����(4�V�嚡��O�s�>Ŏ� �?�J�SܠQ�[���錵��v��q�j��~�#b��,`m�i�tJR��M�M�14FY�
�c��W��-�M, ۗ
��~��oĢ"�e�Sa�pT'>��[5R3�i�1�q�ܸ;�b� _��r�X��"W��l�X7eٰ����Ӡ
x�%��鹬�Y��@d�X�E���k	?f Q��}`k|mb�^V�YL�cV?�
��:�Vx��1�ScX�<Fk��-D��*��L9+�c�8���)>�5�M��t�)����)qO��c�Q����4Ze8��U@�2���M�C��D�VNq�<ڹX�vnm�z�D�>���i`h���m��c�I:mS�o�;1tV���M��|���{�'2���L��h.���8u�ʌ��e�uu'k��M�w�SV�A��:��^|7jc]9<"R7wAD沆���/����*��8��@�'6������?��#:�%W�����<�����渗rn�r��I3�`�����x��E҈4��d2��d�E�̹��*�{x&��d�4��p��P���g^��`N��̽@�C�s(U	7�?ꈹ�nз
�I8�]}^���,s2�[���J��7��,�dD�x|����@�ci���Qةz���l8�!�ʽ��(BS�� �GT����R���i*Bӥ��W���J�d~g-�.H,9�փ���n���nsfx�:����<<h�P��%��,p?rW:9�w5�7y;x��!|��[�K6W.jpQ�r?
9VE&2�5h��O�6���dI󀔵�芶|�6�ǐz�6����gHb��p��:_��뾤��P��E�Y�{�­'�y�pTr��(�����~y��.(�Q��)�GRۉ�I�)�����9N������E���nUִ:8 Ms����g��Z���g�z�P��R�w���t�#r�AY�f	u�J�����{z��dX�]�q���N/	K�CQ��0T�4���Ym�?tL��?@]|�ރ��{�0E�S��e�ĸͅ��7�����~���ܳ���4�4���(����ȏPW����%�$�~3�k��4��>�:�t�����q��s����Jo�F�uŵ5}�C�V9�]Ѥ���E:XV5IS��I��dl})q��`�2(��pt��|ˑ�0��j�i�"�-.����v�V1����%����~�4�̲Ut�]c�᪓D��v�h��N�O\b)鲳X�[=���S�!v�(�����.�׎�Gh�ҙmټ�RfG�99.�`���;�TґK��_����J�PD��dHN�bL0E�}���q�+�4���%���JlD��Tx0I�/������瓀���p�-˃������;�ݞ������Hy�����5{��YTK�q����Oәѫ�q�W���0����9s�����j2*�\�0{��x�,p�^O�T�I�ҩ�e���~����'i/W�-�,��xk�g.`��@x�
_���`���<�=5R�f� ]ȕ�0b���&����a�;Uo�ouT�����Lo��|C*gݵb���N�����L�}�=NJ6~q@{�&<��s��W���8-�Q�s��okLw�6�������U'�7Sz�>�p@(�ZW�Y���Fn4#?��g�D��Z�;�e+�w�,�%��Na�~����x<���z�~�u���d?�(�jc��8��U�E��|��t��z�/��AG�YJ>|s>#W��ڳQHx�uƈqM�UYߚY�>S [�d�j-d�3-J������1���^u�Z��r�����wYF�7�N��g���QOc~��XȢ`H��5�
}�?_���d�a�q�+d����}�N�P�&���^�J��|k�N�z`+��p\8�J(���6�p1���F��\�v+��ȫ0֜	G%�e���[��@*I
��ȉH�T�裓E�牘뫱�wk�E�:C�U�iG�CP��Y	��L^���P$��8�1X��e.�����R����vDi�R�;H⢪\���5Ex��$6!�����14Kit=p��9ҁ�B��Õ*_�:��s*�m�1�[&�n�F��8�[�T6&Y�����x��r���'�i�"/�Z2�n��� �u���d�=�]�B*t��<�ё��إi̤�K?�H���O��Gm���כf\�,}��d;G ��jS��(C��R���m�{k���M��T='�4J%�V����U�TPu�elǏ6��3Ej�X�� �$ϯ��ԯ�*�N���I8����F�&���	����|�HԵ��^��j�R�E�2����y�ԭ�T ��M�^P�.�Z]���&��H�F	��"���`)�ROM|���2�E��̜��-�N�k���O+bS��C��W\�B@|��@�E��9\H��+��h ��xF�$�E��
��3>z��^�D5������}���Q���f��}�y�,�� 2�=��!�(�=1�k��䬏�d��t�	[�A[ �� f$w�f��y������/i����:�7�S���0G3��*Ѡ_h��F̉Rm�d9io�]��Į���o�<��.��/A�������b���~�*�@���Z��]�	�@�;��j�#a�lln_p�C��.}T�� ���4������Z����^��J�DY+d�ZlI��+�ס���ÐR.����V��}Hx����f�\ ��S���ϔ����������~��ژ����k��i��d�2	i���2{HBެ'ܚ��it<_!A��(	;��+���E^n&� UJL�*)ɰg}}���群�ɪ��ǔ�#�-�"7�.��i�J|�j�Z#ቜ���ӗ�$���=b�xY�/}�,Z"��8_i��f�#ߏf��A���F��_źQ����'��E�����
�P����s>�3�3�DnEx����J�L�}��؁�đ�Y����������W�*7�LǠ(�?�G��c񱔰U�8	�b�Up��}����H���!�VQۿe\��b��,ܯ5ǹ��{o�L�#�P(}L&�5�$��qz�[�:Dr{��#����?YͲ��.k����)�
��Pq��u�!�ON�+�e�
	O��QHQo��k���1��LG��7ݗ�%�s���4�;�����?�Qo�v�$�^w)δgD�ʦ&ڻPQ�2�Y:�^G.��3���� ~�A6�w����Q^?��_ �U|n
��I����
X����_h���I#�D�ء�p�$"�:/D�)�-n�26�P-D4�+�bh�n\�j�]R>�%�3� ~��~G��T0B����z�8/un��طs�5̐�'Zc�`k7�O�z'��O�١��>��͗���S
Z�V�d��ܥBVvi:u�nL�-{�;T�YX��Zw��K�4-U43��}����k1���c�,R�R�9�R�����,d=�>������+b]��_�u�p<�UyE0�]���w�/������s|ˠގ=Bx��f����%LN:<�GlO������vl�&����G�L$-4�U�D��N�V�بQw|�����Z��@"n?oRs<f ,��NB��8��с�4��L~dye㙦he@��e�+F�D;��\�����~WO�#)����[hL�a�����sP}d��;�1�r��9k��v6���d?^�"k#P�!�d�̇���*�h�!�������խv���{�+4�3�O�b��7;+3��Lr��M�=!(U��Bsp	v��9`̴���k�ŠZ.�8@�
�����ERշam��19