��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��Nڭ�	�����B�#Z���?�4�j��0�ΐz�A�y�[��I4�fB���_Ɛ���-����B���M'~��k,���'zf���]A�� -̭���ҧ���D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T��P�]��h�� �x��ɻ/�akB�����L%��s�A�ۆ�)�a7�$�HID	���� �դ���ᑧ4(6t��	x�ō�Kh�/h�}��>�|a���r��>]zu���f@-<�.2�]ޓm�D��_�!���Us�e��Fl���F@��.�zn�^!�rY�qE:$�Ĝ�l��8D�V6�!�)$D��������u�Zp�u؂E���7<�Qaۊ�.�� *�Î)�$4��K�B屎	�,�֯��S0�"��M�����Ҝ��Xq>ڠk*P]�N�S�`Ѹ�qZc\��J���0U�[���C�|��/�pQ�y�6��e�5 d���7���bh�Eu>�[�[s�an�uAJSS�'H�h�n��@���8ʬ(��'�W�j"o��seQ"�V�4�!�-I����k�y��t;��5��ĺ?��{n����J�d|�������z�ϔ�3�v(�&N-��Ro�]�&���gL�LUF�gT���\�^��}��pN��'zP/0+t\��zag)d���ǈ�� ��H&�s�G'uC^]���`ڏrA���`�����\�!��E� JC��o�lƎP�0���Y�>5�3�7�j�b�e�F���Ӭ�@Bth�hXe����k��� �?�'�Y�d�V�%�T�߾���H�*�M����=7w���=z �#����Y{��I�a�t�=���ñG<�.8���tT�$o�ԣ�p�;K4�Q�|�8�uGZ�����BÁ���&�~H�x����Vi�����a�P'R!ұ�TB�)\�������$��j�&w�"�6t& )3tu�S��m�+�[-���@��|ۜ�l@Nؽ0e ��N�_tweG��y� e"w���ᖩo!h� K��ɽ���Y������`����w뀠�^��'��� �ִ�g�P~z�)+�U9
9��g�i�ξ�h<XO����C,"Fp�"����x�l8`x
�0��[�:	=������e�$�_���k��������	_���'X�;M��*�����=�Z\��#����j���	X2f-�����x��j%[ᦙ�;_:����p%�X,��`(/�T����#�1d�;�y~���!�e:7�xF\&).��?5���il^1cIrY��Y+����$X��A�+7 �c���S�������=]�'��}m��qS��a�'��,��t�v����q�KDcŻ����O�qe�V.�T#my��nE7R������#������׌��Θ�f�K�"�3yVa[NI��k�yɫc�Pby�]�i]!n�M�D���,��U��pk�(w�H���*L�i�3�a��i_j��=.���Z��1�9�<q3���YK.�Y;-�)w`[�?�+]��	E��k{#����u7�z��]b��B3$��������7�6�65�$�h5�J><PEa�t�u�W���ː�z�0���A��˕�ck�3z�](���|�g@(��}	�]�2��M���nJg;h�C�1�vgumG�w�i�6ɘ�|}��z�<���c��-��ȷ/o��bG~���E� hd���V���Q�=��?T��1��'$��ʲ��A�h���
��y$�g�n7��k���u�s��v�$��B��lHT{��њ���ol��?�a�u�;��g�w'|zyq�Y�x;���vbz}~��f�!Бf汁���M�KO!	\rۺ<������ j��i*߿���H�d렐�k�3H�ʙ/�+cy-�h)��j�byP�����!&�Y-Py��oܑ�L83̓�i�s�l��t���Թ8�X�-���<��u�ck�u�T��<h�lA��Is\��RÁ���<� �P��|�g��Ow\5���+������Zξz���!T/����׍
�²��q3s�	�Qꬥ�{'@L�g//���^��+�J���[�E*/�Ar��u�Z�~���Z��h��LT/��s���aN�r6�^Ɵ�g��9�ri���A$h�Jc0ѥ��lY���E��;o`�v���M�Ӊ�x�)�vpv'W���� K8�o`��5N�X^Fm����ZG.�▁'����Q"23z�Y�n�$�e}�i�e.Xҟ���D��y�)���z `�k����,U&����F.^����Ƒ>�^��^nJ�����2O����u=�]PM���8>�:[�A�Ȍ���q��D�.��Uxӂ������,:܋�,�\|���w�:�m��q�M��Iј�e�&�N��[Ì)��HLoBlK�����Rq*��#�9����/s�5�=G����ǖC=�a�4[�e��Xt�em���~����[O�WLmE��]DTFo�J�A��rN�ŕ�Lx9&��n��ַ�7�(�s��(>ľ�2%��7@A}�{�Ab��n�]s��~��:+��ok���L���p^��0��1ӣ�D:{B(�b�����Wו1�me�Q'���}g9�dIԈ4��"q0��{�W�[L!i.^���̚pֲ��&R3�{���.,)+sk/	 32T]@�F�7[D���� p7X���wE}U+Uv;��B��p_�\,��L���'Z���М7��u43	 /yq�(��ߋs���f�2ӄT\�6�%�I� ��w��ɰQh� ������!��a=Ey^���f�aF'��B[6�N�y�2�7w�4{��[����҉�rTN9ʰ#Q��DՉ{�n�=��h3m�u�>Ҧ�����ծ�C��.'kz"�~E����g]m+�����.wĀ�uΊư���mq�&�giN���t���15]ټ�e����w:�:w�a�@��ꘈ'c4��s;�6+
��&K�|=v��� bh����)�����^���0a�ݿ�#�[�#��B����R�aގ��p�	�pM�k»_x�-������59 �b��?	V�U_BN�|��X�Z8�TJ&0;{XC�q`q�1�����A�ad��/���q�jL�sO;-����nhV��
�"9]a�=܃@d2b�b�31lZ�b ^�R���	٩��Bad�L�#���<|�������!�I^��1��Xvq�We!�eV���k߰jv@���*[����8����ꣲ� Ը[����D&X�Ts�5(������	̿��㨂U�6s*Aq=;6,�#�����`J8MY�%)Y�����k��RPz��7���,E�F��пE����}�$�0�z����nk�o*��k�Kx�$�`�ZFU���ω�\M�#?��(��)z:c5�UK$�wT����n��C���=
]�$�Qro��+�S|l�X�-�O�t>�)�a�;��}���e��J��k~���� H��#U׾�����8�B����շ4��
(U�s��1(�쐃��1�K����m���l~�UGE6�ڼ}�v�f��T�#���n,�s���Wq%^G��_��)��*q	���>.�*���rً�y�d���i��j/vÏw����Ȯ7�5�z�I:
�]K���(�q5�&v�O��o�����,���7�B�,�R��ش����Т�YK��-��k�J��nG�+��;{!GW[*�{W��d[�>��1n4�[��{9o�j�É��?Er6"���4�7)3rH$�ʓ=l���=a�f�mwݪ}���h�	���i��=&//�o��x""
ནw+BO��i�,L�r�F�A��%�,�,�� �\r��?N��C����2���$X�y�m�xnk7/�����^;$U�a_Ԛ�-�&g[+o�Ip[/�|U������^��{�w��{x�|e���X�1���+�Jb��q��V۸�8l~�G{�F3���r�~J̄����#G��).�ۧL����Z�}��w��=�o!��$��r�Eo�}� �9�$W�W8�w�`a��,B2S8�s!E۾b��8 v'�oG<��KI5���Q���'T�����~Jc�i`"��7��'��M�K���XT��^��ɹ���$���	~��˄�XA��Ɯ������C<��"D+bP� ��oS����������=�,��� Y)��@�/�׎b�A�/w�b�wf�3�cyB�IY�.� ����*e�<g���Wd�̗�@z��'�N��a�ۚs׵��)P#ݟ���{�W��1��.��MH��t~k�d�U�b�RƱ��فq�z�[�_'q^sCJZ��;Ox�	���)FG��{�����"7(�yDA��d)���]�}l(�|�浌GOn�!#�v�R������El\~n�P�L+�J:�y@Uה��(��ubQ�������(�s�S����=�êh�)Z�A�]x�4��x�~�h��G9%�5�,Y�5�A���W����E�jgܲP���B��9P�<�4PM3揆l(�I�K�_�����Ն��22V�Q���b�L.��4�n(���w��^��B��	�p㈼�x�M�N�X|k_n�;u�H�u�k����T/������h��[~=ӅXh�y��_�A�r�AeP� �~^�ucx��P��$*;�0[D���JҚ�"��e������=l��H?���+w��'X�4���^�����Y�c#/�;Y>�y��
|p��E�a�`R�T�Z7�l�o�#������T���I0�^�X`��f��/�<�";��, &Zp�I�mvb郾�3�R@(���
�z�n?q��h&��z2$��!�1e��gGJ�G�z&Ǝ���h�ϭ7�D� b�ַ�zjϕ��	�e(���
�	��s|q��u5�����|��{���.pX���h	��*�mVY�B��p=�7h����¼	£�,��b�4�_.��y�VT{o�8{Wh�q��|6f��t݌d������8��f���uFa�c~���E�x!��v��8�6;��_�O�=/�By�����%�3������V�6�8kF|����lϟ~����Zw��Su���&�<��p���G��n��R�����Q�a?z��X�/��p�+?aB���0�b�U7ñ�[��4H{ВT#N���,RP]�7����g׌]H�:h����`���`��>�x�K�QǄt_���<�z��3�#�Im�ot�}IڿJ�H��/� j+;2�� #�4f�|Fa؛��X�͕\ң�f8�ׁYӓН�ƾbv>���x^`bd��&����l�5 h-Oh�j�����J�s6*0�����6w��U+n����R6!�s�<��K����q����,�Q��y���Q*�6&�]m���e:��#��ɓ-�=/�#1�K��X��H(�6)�kj�ҋ��R7ˮg� ~�Bb�Lx�v��T�s� ?�U�.0���IOz7`�?�zF�&`��/�RD��lS��.�ַ��L�ה��X� .�.j�Z8|�����l�kj��1�V����Lc�E���n�dQ�����kP���`��*p�q	�����cV|�(E�H����qO{e�O{>�����Mw���'�3��B���4˹�X?�@/H�_���F���\���st��9i�|R�tИT%�T{-��=~���V�,r���,�Sq�!��Ȧ�z3�Ⱦ��@ԯ<	6/��3~Y����#����rh;�B:�&�^���
���<+h����G�醗�,e�Z[��4m�{P�wy���5߲(8�y#?�cd�w82��g3H)��خ?8i��{� 2��3�9���GU�݂�;�@�������>�N��v4}X^ߴe�iJ� ��Ԋ��03g���;͔6�p�軬4+{Z�^���H�ԛ"S=y��_Y۬b%���倆aõ�ygG�s�Ʀ�2W&�*�&�^�2�q��?���F�*qWb�\���(C �tA����!c%g8�T_��/�#d���+�G�]H��i�z���>H��ƈ�(-c��]l5�_�z}u^�8�o�E���V��rـd�,U=���q�_�{-�0�)�����o�q��w*��v:G�0@�K�Mʃ��j1$�E�T�K<��KM~���wd�_����+����hI�k!Dfϕ'���G�.JM~���"��������6H!���%�9�6u۠�h����≣� ;Yt�_fv�Li�	�z�� ���;L��4�K��ݹ��<3�7LIGAM����E��EI���S�rS�D���ү�M���(* �({S<��kAc&����a������q�s;�"��Il֏N7�,{!��E/���h&I����
�kka�����n��n�>�������v�"�mM�u�k�j��[xz��ºXRC��m����I�-�����>��<![s90���ˇN1J-�B/~M�����f��.3r"�� $��J�[�K�4��CbdD�zi�C��z����{q0�E��mr��Oo��ԔC\D�4��q^�Lm�]3����_m�B*�C��Rk�\��@,ҮC�m��%��<p�Q*��� 	S�ف��po��8OaЭ�X�48h����;�ø�ږ�YmɎfꕑ��+Ft�y�+ V�����zo���4�$5u<ɹ�;��m8�m��|�v)e�v0�;B晧�P��w�ϐ�@�6M��E����ڶf�U���(QO\�͗P�&%�v=�iy��d�)e��؏4���3��_�+�s���wubdX=(�5��o����뗭.=m;3�����dH����]��/��W|
�yl
��v��f�2��p�8T]q\,x�@2�K��]F�|NSAt�e�!@���O�N7GbZM^��O�"L!L��¤�oi�MS��0Ҽ�	f�5�w�g(�����4N�2Z	�pK �w�%�QI����z�6Μ��� �"��7�{\�e"�Pcpy[����Y-1`�L��ț8ђ��}5�b�����; ��K���5���и�w��h���؄�0:��f@@
��aL��I���f]�6�tR|R0e��?��̚{�f���z8@��+4��4a�
��K�D]9�0!a�����ps!5�/�ٙ�}�tC�VGO������	�b�$;6wЂ�rV�����	͖�K�5r�hl�J�#JT�b@N��ӻc�^ G�wQ����\#[�[�̒}��܍�� Z�[�.��i�)��6��n�H���{ˆS��q��/QaK��=�IX�߾>׌h�՛B���y�.U�Xr,>ʂ��k�纏:Q�����x86�r�&=_ܼxp����Gd�j㪔<or��6C/M~�K~���v���+i���˵�:?0L�k�=X,�t~I, Wb���z��k�C�D�`��e̸��I=}GsV�s��㦪|��6: ~��	���KZB?;��G����K������a���t��\�y�}�z�ئ� �0x j��6i��|��X.N��kFY�jeGdiO28�L�v���W�j:�_���YGq�YDZ�JK��:=窊����{N��]5 �SB�����U��������t�No����b�� �_�=���*|���ˑ�b'u��]�BZ�-���'z2� �
BsI�
CW�w�Y���N?�B��x���|]��4D��̀Gq��f�e�4l�+BiN�D�b:�`3���F&�i,�����i�3�g�>хB���P�,I(Ψ�S�J0���j���d�A"؄*��c����d{8�-��f�i��B����MA@��s�O�TD�k��zVv֦�D&��	FF��?x���\jwrQ�t�8����U 1p8�F�O��ϣ3BFiH9��0t7�����y�i����_�l,׮�A!�#�.aD�{Z$�V�ƩJP?��l�w���l�p;��:�3�9D���-�"����<�bo��#�a��� o`��_��q]*H)-�OR\ξ�nP�p��<��:f���m��e�������E+auQM�"d����%uKez���d�sݥ��}���B����`����nq�7I��	i�Y��`+�<�͏P/&ѕ�.$�C9�!�k��# �4�6۶=���:�[u-�Hʬr��u�[��P�L�,\7�3�f�<�/�:��]�),n����ivi��v���Η#/�����
��6�Ϗ�0�/tCԻo���(�؈��啿��a
ȴ����_K���ܮ�7������GmY��R��<5�_�|�x�!��](�	�?�/�'q<�Xb�;�DVB�|S�������_�K�W�p.�k��9R�J�Y����k�/���vFwߍ0�|Y��e�[�
�W��1-���7p��+�7��2��Jޮ��\�BS��ީ8H�z�eH�b�����@�@)B�ƝT�q��2)!���;#�/��&"*�_�_$���.�ՙ%5)t�袾��;XjO2Ds�[{���(w���c%��=�	�������D{$��pa�Ms�N�����4�E�I2��6n�g�ǣm]>d��㯲wn��?l��?$�&I~(	��>��bQ�WI�d��5�y����i�ExQ�˰`�nO*}U���|?��ﾃk`��3��)���k�����/pl�'��#�>�����&F���%U��d���J��'�B?�/�Xc[�~�T4劫71���
��n�Y�".&
�x�Ug�4B�P�4�a�7B�n}�^;�MšV��{J����N���������o�|:U�_\�,[� ���L���E{���n�kD8*�Q�܈�D�.B9��<4�X��\���V\�r&'@�����k�AVåJˣ�W�h�R�+�{,S��e�6�D-�G����� �X������Qݬ�-׳�~���������{��.`$I�,��D�4ٹ�U�¶�.�/,��2����,H⥵���١1�����|�H0	�o�H��ҵ.�b�6�-����o3/C�Տ���Gn�HJ>�x�[!48���%�*����cCɯ����q������,C��J� q�P�7n�i��TB�4�/p��w�u�>e�B$\�)	����6[�u1��F���	a�ש�t��+��v�p���r���<]�H⒒҈�+B�ڭ�/ g�BG�l�7dP~e@s_�=6�S�Ĥ��@!��)���n>-�|�0��o�� ۨ���C��1Q�`a�U)vY6��ѬF��:]�fA"�{l�/��z�1��&��T`�ː�7(�^+V��0�Z�nX�n��@�g�\^�1��k�E��LY`�2�H�C\|�pG�I��;�K�:�r}�,���L*)~�n`�Ùx�`�f��Ѫ�U��󦨦:�+���ڴ�Iˮ@Ȋ-�r�^�^���8�Cr��/r�kק�)�m"��9�����w�@N-�����4.���~Dݚ�u��m�`C��o\ `;�i�Q���W�����,���c܁0�I�f�:ްH]{�G�>sA�ɜ����0�D��u~���������b-*�p�Hْ{=�6٥�^��3�d�����5>�A	#ƨ��(!l�x1�Ɲ�̔S��\�?�m*u7�4�`` �G�|�DUon�����������qL�����p��&� (4
k,�ZI/3�Sq_y�Dc=���k̢FPl�N����c_~��^y�^���0�֒K�h����{�0��.b�����9�^p]��[N��O�ĭf�<~k�������ڐg��>P[Q(�)̳�x��������,����� ��`P`��U���g��_��J�n��d+�0f��W��>PyL���F�'�𜝚R�{�S�:����ř-�Bl��bH.���;-�׫�X#�qb������[�>�=Z��ET�v��^wR��֣��	��7�B;n��d�+e9+	��'���3O�p�uo�4��_]��jp�#�r,��@A���|P"�� .����R���Z,n����\��9�c[���bo�8��_�6������W���ȋ�� �(R�|?�z�᭭��w;A�R�U,]-�)���*�]�$��S���[?Ry)�en��PZtj�gz�O��
�.P���	�I��2���-��n�������$c�-�Rq$}��[;8��贠F��Q`6Mw�7�M�%(i���z�D��1�&=O���ѫd�?�$�#SE-NJ[R�֎4+�\���Le�ld\�?�u=R�ҭ(��'��.���r��0Ӝ���xd�
O��d�X`��q+��aL?n70��ݖ�J��_�NgUZU�F����uc�D8�o���Q��-�oU�" ք`h��Ͱ3����L�����|w%:}����.+�Q�e�f�������8�
��D��[&hIf3{���XܽM��k�f'#��/�0�I�(߼,�25���*Yv�c$	J6���
Y�=�U͏�~�u�wj�\�U�a-��zɜGYzu���O蛜����ԋF!0�olv�8KʈE���h���^�L��f"h��pnLoY�G?\�h~V�!�d3�.�U۬'מ��:�x_+y��"�5�l&��>f����d&j�@�\5�0u��i�gD�/���q�϶i��Wpd���j�%�qj:�0,�9Ya{�.$�m���3x�M�^r�F�{�wZ)�(D��Z��Yz���������*��&��J��D��`�L�����V��xwQ�v$�R.?�r7��Q��4ℊ���C`������+7d�.ܾ������Eg~RD����ZΖ����6����x�^��T�YX��퍛��R��"�X�h��e�2��A����䍛�W��o���QP��t��2i�,��;	l1��&�ݣ���i%�y����tI��`�S�x���I�_I=Ci;s{	x��8�L�>H����Vc�_df�𵻋~ zc�xq�i[���
��k�P�=�I�{����61Ӆ�?�G��̏.7�>��3�{O�H��g��C�w���""{�Kf^Jk��6~W����ʦf?c�2��#>�<<�-�~2Dm�i�U�Ǉ�ޔ���D��O��j�x�x�e{+t��sE9��|M��he�H�=%f�j�J���`��7!r�]\�����?G���C�Iy!th�6���p#3&:��-s�A|EFw� �M(�qK~�S�����OK�g1Z��E;u͠A�YsuԂ �'�>1Ok���)��f6Zp5m�����)�(�ڷd��O�Q胈I3��*��[}9%m�r�.��n��d^#3��L��o��ѐ��;�b"�@[1��<�[�u������Pbg��r�ݚ榾��oZ5J끮&��	��}��>�}�ۑ+�N�_S���AtlW�8��'ϙ�U����x��l��Ь�!��f93�-���+���_��`�Ԫ�E�6^�����d�^�0�6�y���OD��Td�4���.˕�N�fe������p3~6������̓�������6o��~�"��t�v�i'wq�l�);�p�m	�R?Gp	gq����+Oz������G�Y빖�)0~&-���*��h��.eKC���ʭ8
���6�|v��x����؟�7N�1������������Z$���U�u�"���+(�M	8Z�I�T����:.i,8W�=$�
;������)�V w�yƊ��{��L
�E�=�OK�T�c�ٍ�ی/������$ȏԡ�1 ��u��nt�u.@���,�N�S��R�>M;���2m�@�:��ʆ쌗�M�*�b��hÕ����Je���N@;�>������>���O&��[�)��K����5`� $��c�y�&��n������G�����Ǎ9zl�j��4h�zh3�hG�Y�-4�x�#�..VM���ġʞ@��^�fW�-ߗ�hE��~)�V������n�CKB�+U�q���c�pd�h��B8J9�Z�c2�����c��&�� ��i���+�uv���ϡ��_Ϲ81&�沔0؛ZG�""Ի��:oM�B����k���Tt��+�^����t��ƴ�n����J�Y�ֿ�����|�N1���u�>y_AL�kcOeI�a'�f4>�A棹|������#�X�8D�K����wZ���B
!8[����h�5e�ll9�B�RP�����=��~"�����>W֕s<�Jת6�F�2��Ɓ����b0[}jgb�|ק��`�e�0�~���x��ǩ�P?�����*I��Ǖ�$���UD{=���ʴI�aN�G����V�&s���_W��լ��Ft?LV�.�}	�3�q=��x�H�35����/ ��q�Ȇ�^^��>�A�s�4�7,��E#]���@�D�?��<+�����`��+x�`r]x�u� 
ej�lc���Yc8-%�O jt���W2{bB���Ty���������q����@�D\lc��=J����l��?�N�v��+�T�z�m8Xط���N�?!j��1Л�$���H��{�&��]`���r�}�ʓm�p��-�ʱ[�M��\��[�f����X ���'���A(`����NU���
o��~)���s��Z=:�łoB#!Rǡ*~{?p�'��B�xk]5:�)/�����?��|��,h�#�Ē)��7;<��'��evȬ�'Sp�2����O�I0Z���)�W�շI�HFz	aY|�1\��B���%*�`�0Li퍀����2�P�E����RP�"���2Qr(�+�w��`�X�`�5��ĩ_{���L
�U�N2�� T�ݑ�,\v������kU5���ɾ8uI��r���Z��Ҡٽb��hj_a��>"9jM�TQq/H��Fpr���N/ܴ+�!�w�"4Ej���'�v75��!p*c�4y�Uy$&:�e卑�!~PٗD�rp�$RL���K�'|���n%�6�h��a�0":�9W���d��w���o3�ޗR��>�sm���R�WW'X\�BW�	����JD�DW�dx�VӾ��=���Q�x���e��4�Y�nn��/�!3���}p�N��.{[�^�o�|�j��_�*f@�`��ŗG�P
�RF���Ϭ�Z6:��� ��Ɋ٦����w���G>ȯJU��l��̊�!���9�s�[��-�$.� ]�Qn>����l�����y�t0�^���qY��_��u�����c4�|jW�:0�N$7`CeԂ�Bf��q��)��aj�GC�|�ROl�>i���?�L�^�n�;(4��o(#U��]����y4UN[\
�`s7|�?���X�	�R�&���짓��	>^�y�}��]Y��X�f&�y��YZ8ؼ��SM�:T�D2؈��C|��Fssĉ���*�=� ���#t�Ω��u�߮��Oۦ��/��T�����oa[�}�\�$b��9ӻ�3%�gS]��mcsg�0�L	�2+c��'�~��g���C��'��Ѓ������&�ޗ3B#�����ppHX<K�ˤ�O��'�ځ�G��O��k�X�����|I*C����s�v�>�_�uW�b�/r�t�9�\��]���<��*���+5�4$���m5L���`E��ށ4D�'���;$ޜ�Q�]���T���z���9�ˇ�j]��$��a&*9pU�N����<,��6�ޢ�pm�א�aց�|���@y�S�|�{�G����)�������1�*^�B��*@E��=��\��ӊ
�i��>��5�7�f#&��ɟ@�*X��b��!y<�5��j ��F�"�΂Y�C;�Pxk̦5�̦��^�^�ٌc���������w�ϫg�{����%o���x߮|�K�nM��xj]f�旴�3�;r�-�J��4x�(7r�5裡�q�h�!+��Ʋ֊_`��Xf�WK�-ƶ]C�F~�t\�v���f+�z�\�5^M��ޑ�:P�
:��,$�0�^���ȓ��L,B!=�JXl��b���2��`�a�d�t�E7^�������x��"iZ�-UO)��iND�r��y��Ͻr�׵�^��?D���� �#k�6p��`ʞH��a�P���_n���/��?.uDP+����묵mI��	O ���aY���^RK\d�G6mP����(�������U�^>ߙ��ą �b_mx@�8T��ԫ`50�C��`���@���άG�#.�޴1(�����{��@RR�_��b�7	쿦E����g�{(m�JMWi�ʚc�����uIt��z%ܟ{
����/��	m���~�i�E�ǉ���"��x9:�w^?�KłOV9�P���H�Gi11C�o�)�?p��d�="c;t�O����e`�=T���=��9$�F��s�L�.r2���,�Ջ�C�J�m1ْX`Sy̘��c��R�B��V+*��o��%!5�*k:tQA� *�u�G���kb��� ʼ8�|�	p:���l�c��$����\�ݡO]z@IM�Z��O�=C���D)!�u�a���o�2�jD/�XRwհ�UU�z^���ɜI�[D�X8i�h�y�F��Se���d'_6��tB�3iǺo��-�� ��l�`[��J��`��>`�y��5\�<6 X��1+?L�Ƭ�f����l3���_�#Sj���B��0/8C�H�!�!��x�7�>�|j�.��"n�'��f��6����iG�j��\3׬@k}o�&,q/Ed�i�Q���Q��8&3�X������v�2��g�W�V���gCt!�m�ؖ�P!�j��X�b�	3�ւ�Z�s.Y� sYk�,'TI[nV�"���߬�2Xj��]��C��xm�wC�y��5r�	k�U�����0�xoޝ_�(&}�YK7#ٹnO�����zj 5��xQ�a�����A^P�5Y>O,�ͼa�C�����-�%i]A(q�_B~K#'�Qf;*ǌUC =��W�Bu�%r�Wn���D�:PTď	���箑>��$�����7&e~�қ7%PZ��2hW�瑭���Дx}Yl@�0d�L���-�}0�5��F+�G�cq%O���
���[W���D���s���z-1ώT��uV�SGs*C!��k��aG1)?#MZ$�[���"�t�#�|y��V��M�bu��*��B0�5�3+TAK	��.7��6Io^�v��n��M��T�����VO��H9�;�}�B)]&{��kW�K��g��t��0�Mi[`�L�㬇x�����0�s���>�?�g�l""�^7ֱßr������3[e�b A��rq�Ӽ{DT/��Aǡ�`kt�g�3�~7OVr��Y�I^hi݂��:X��;g��r�J�;�d|��?��M�M�<Ih-m�7Ȱ��9�,�Gu�M �����-���/���Ny�B�ܽ�E&#�]��$�q"9��s;���Sa�2[}��R��,D��v9��4r	�9CV:����J����2?��m�:y�i<X�O��I��aF'��X�@��ѣS��L��-�ț��}�?qN5�idW�_D�zN���yִG��;=��
�a-iÜW��>P��[�N�z(F�Fe��[����?��c�<�����?��#���7�fG��W��k\e=��7��H��,��>�X�&���f���1Fu�#ِ���b0R���URIĜ�����j&7��J��l�f������2�цf��Su61��Я��B�Kb4s�zT��( Ij�����`�8���K��Q�?��Sm���1tC"p\9I*A�?nC���ηb���!V�l����^��
�h8��.5���''B&Y�Y�,R�G.���F��w2D���`/����0~q�X��a'G�Y��<��x_����f@L�h�:m	ƲJ�@C/�2gu	L�l��g�J�����8EI��)e��̕E焬�����R�'��2�2B��v�mhԍv�y~��ÕtP� eDN�U[�ͻ+<�s���ڤEt�~���CW�mm_�ޙ��(���C����i����c��|'~r�<�H�AX�t��b� �::P�.�cC�/<B�|��h�7�Cz|�Q<���R"Due��ܑ�����"l�u��#Q����Rk����K���R������q�M~��s�t���A��!.�4��:Z�6Q��{s�d쌇q���=	W3��$�=l_� "��j�3�d����ϷՃs��hs0�g�3���#(�!��r��oD�p0G�#O	V�Q��76s� ���B����R/�?���]�CA�2�|�l�g��oN�P(F�se������$��I��ͰLnn�$Ź��ύ�&�V�MUc&�%'��3�[菌��f�~��䤆:���$6M�)WU�mA����u��k�FИK��߄��h�Գe�;��ȗ���)5!4$�Y����#.=��ў�Hp����P�������c
��ч:�aOc(�xڧ��$q������`X��H��k*}�eu��i�ym�(R�t[���1z�'����T���"��^��,V�'×�Nw��*>*5���y��~JW�z�ų�s"�_�m�_`�\P���m����\i>d�  �ðr�՛���z��~dP`�=�`Mu��*�գ5��>I�!Bn�~6��a�B=���]ZT3������?S+S~3b�:?d���/�{pN�H�3������黤��6�U���+���U�sظ:�%޻�T�q���3�z�JX�y�O3��a�mV,9a7�X�r7��'.�}���#ʫ5�zdX��A@�' <�9e9lOW��b�K.i0�R.#p�E��6�u���I�>�)	X�_�@9<jz]Me���m��k����N-��� J���o������ �f�"}ލ,�&����֡|
�E$=�RZUT��9hQ�X�=�sc������������_s��5p��c����a��|g���=��9cl�H$qO Z	���q�VƑ\y��f���{�|��:va&O��"]�Aw\ϝ�����|�;)$�\T3��j/@S3����H�lB�ETw���:o�:;9���=�r���h�0�T�'y��4WI(ב��6o��}����uaڮ���\g9�iR��N��2���:yM�{�t�(�١ފ=���؊!���2�mz�*��~Xԧ��N�ݟ�Y�M�_���s�h��7�e��U�L��Hg��lC����j�*4�߳�V�1<��r5Y�-J���D���e��H%��-��W��lDg��^�F��uwM�񲥨��B� t�ٛ���:�j4*��7ϋ p�X��~$Fe4"��|�7���1d������>Ő|> 	�x��%���ޮ��6�� pV�I(�
a�|�Аr �t�s����n����x��qg�b'S�eC��5�yc�ءAj��n�ɉ��sF�Sn9Jη
�*��.�Jc�6�`V��ݨC�nǘ*��S���\ֈ�a�y!2?x���Q��C�$s�T�K�� ��MU	�y��^��!�����z���r��~],��D|�j��#IfxZ��e�P�?�^'�p�iL�a�-\F	,{���?[4�����w\슯�����R6�J�Nw9�$w������/��	�J8�e/ֶY��P"]-���Ne3)R4�1��+$�O�2���6R��^�Q/�TJ�-�<�r��?}]%D�V��y*�Q����?�L&a#���(�����I��g�^�����"O�Ct���}�ZX�˺@�%Љx�+V�I���(�.�O�a�IUs/Nc���:Ę&[�#�z���y���`�%�[�\���BC�����~(�T"׳�S.0#ꯧD�s�����i2?�9]�ܡ�#Y�����!�Z�pW��U�7�E��w&�_��vq��)ib7t?����?0v�rqW��97�%�3L������l�l^A�L0�AO�� ��y�Kvt��W�5}��W��LZ:��D��$��컞��u�Tkx���o��z����=����5��5��8����r��Gxs:��:�NӴ��-���.��wbL����nS�\G�x�A�q|.~f.��/sq��$�(�� ��h�Z�L��<S��GU`�jZ�D�lnҒ�%�^�8��'ea{�7@�̟eηѐ6%//����LyM���A<`/�����*/��
W� ����O�gBc3�����ԙ{)V�T/F������v,$g|��)�4����Nl�J)οr��g�?�}�ާSZ(v@bz)�i�*H�jO���/E-��/B"�ە�����<�n���%G��j}T:�q��g'W��b�-o����mN	Ǒ/��V{�7)�T�����I�`,@X����e?�z4����	�tq�C��h�R��@��3�#h�d|��A�rX�k�����/�$Z�B��M&�e(����.��fWf����e���q��)!y{�F�]�2RPϤd�bznڛ�T��48-Z�SXȽug�c�ӎ{���g�. 7 ��o�"�%�R)d3���qU+[b����#)Q�	��Ʋԝ�+�:�'����Tq����M�F�X��ӶA��M#0qQu�z�E�zd�R�?�;�5�Z4�s+E�D���D��ɠSD��_A�v�X��&+��e^:�:&-;9z[�vэC!V��XF��йP�:;����g�H1��;�߾�$i��L��Eeg�Cu�m��nՕ���1�N�Ŋ��P��9CJz$51{��̐��:�~����ow`AVڌ�ƙ�Y����bߏ��Q�.U����n���g}�rq�9V������6������Ry� �ȥ��VU��J[ ��O��ւW��:�� ���f�.�o����K�cL�����α�.-R&J�Oѣ�J����I��㐫B6���12�iQaۗ5n��ɲ ��SS��l#<��Wl��j�$��a��W�8��D�\�����"�����)�Nzb��x�p>�AӪ���_���=����3�(��V㱠p,��������h�'�Bq;[0Υ-7�}�c��%�v=���LB�P|�Es�ͳ@�^9zG���x&o]�{\�������֋�)G��t�D̞��W��}Ƴ�08,(�w����ڸ�jal�LF4���Q0b-��9�݌T�Y<��B����A�}��c�)�;����,&��_��x	�l��o�A.�2�%7��c����o�������ǉ��:�|)�������c��q�������W�f;��Uw�\��Ke;��P:x�s�F]��6�:�Cȃ<�*���\� ]R! �v.lz�P�����{���M3?�%�GoƼd�|j�s�-�h�UVw��V����������0B��RЄ�y�
�t�	�6Qv-<�N=��|�P�C��%�܈^�E����!�"fW�ׇ�a|���ˈ�1)J :$�s��Cz����eP���4�}��}e�Ghw�z�7�̆~I�G��FA�����R�ʃvy�0Fk�(Fwc�o�#���ƒ;��d����?㇈p���a�I�l�l}K~��� !�N�,}H
@�M�ۢf "��k�i�M�s!�/ʜ���-�l�r�l �`N!S��E��i ��4.��2�TwJ}�"7���;��d׼+��yΕ�*:���{���]so?�nп�X&Ā#R��	4l{��5fz�������S��u��=Ѳުp�,���4�
������en��+<���
 >��$�/5�(����3o�;N�Bue�F���	7F�A(��@*�n�է�"����қkV�
�j�9S\����m��B�Ue߶�.��rCtӮ�G�~H�D�ń��ݽ��J�l`Ѕ0_�Jvv��W��W9��8)P�Ó	��H	�{�����4�0�=�N�:Y��ʩ��d�8xA1��6c�ez�^�6�f2�����RG��gsۑSHklS�.�V�T�9��s�F�hǊl����q]�iI��Y�9M֙T���E������ɏ��T!����T����#��.�y����u|����0/{h� d4�gg���Ô>R&W���&�VB��C��U�A"!�T�nMӔ��T��/"�n��L�ѿ"�ʠ̯�Uv8�5JMH���M�cB�s�P�d���W�#�:��@�