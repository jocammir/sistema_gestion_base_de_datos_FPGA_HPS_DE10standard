��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0����_���3���eĭ)|u��XXp���,�* 9w�����r��웺���#��e�jk£���^�\_$!�  ej�)���s������qҎ&���>��f�UɖD(�ee�,��� �M�cNG���d%���j����y��_�m3�[1;q�o:W�C�-���ih�48 ��#1{p���{�=Yl��B�	�K��������s7Oia�"�U�3�C�!Z��Y�V��˼��
W^���~K�)9H6m�+@4|� �N{������7�&���v�{9�$Nôi��m����?�|T��B��i����c�B����.���朙K��t�E����V\ѯH�S���z����
g��qM|#�G9ڭ�vOѷ)N�{ჹ���T�Hg������rP��6�j���*� ([`��!_�@����N��g��a��7���P���������1TE�)�)�_�%OO���G�{���9���Ø�2�*	�pg���;T2!�9�n�ڣ�*�Qɓ��<Nه�Gͽ�OW��`]��O��:���8�#����͐������Pz�UEs�ý`�����q�;5ֹ����]�T�x�x��Zx
؜x@ �"��Ie��;�YT6����ۚ�>�U��=�c�m�quF���BB|�m�.J�"�vP4璻qEߊjk!p��s�˷WFP�"�wWA�#�bS#�&K�DMዊ�����Y
�fiھ�'7S�ď�x�Z�k��'�~�����~�R����lʐ�Ȍ:�R��IlFc2V5ȕ�-t�2����m�R���J�H�)��%�����ò;�7��Q�ǣ ߢ6zg+�ȭQ�-���1�FFv�J�A-x4��l�X�6 RR;HnBh�Z�﷡�x�	�5�C�%��'���X�>v;@���qX���n[����kRؑ�S���T���h��,����W��C;�p�%��9J�K;�ДU����^�e��v��}�	��,�+Lk�������]�S�1nf#[^�'Jd�T����R�&4����B���K� �J3�7�t�J- �m]u>M�����c;�͇V&�I� ��r6<�Y �RQ�J�~�=W&|���,��|���9_���77��Kk\N�5wdM]_3R���� �<��[VW�q�Ŗ<h24��#��Д��h�h3��4?���T���>VQ�Q��| 1�D	�(CǵT�Y�G&@�"�_�Z��	���e�0 ��!�hI��(��6Jw��v����Tzp���z���%�tʜj4w��瞲QKuJ�B�5���l�m���l�#�3��xL�#�%�'�D+����.!Q�{�#�+���v������3J�����F0)����n�_')s���[�a�x;��N�ci��6b%�b5�q%�!ÿ������/���y|�����5���UOK[Q\�%��p�kIs�Q�ؖ�J�ҫH�|mO�ga�D<��.l�RWdߴ:�c�8r�j�P�Xa�ظ��g�Ix��NT܆��6s�?(X�|N�L��@���bmy�H����%�u�ާ���״�E�4�!�o�=��C�p�?�i���ZگCӬE���ۦ?�r�t�vGc"�dDE�G�ͽ��;��eM��%l�y;=��dm���<P�������!���D�]�?�$AN��fj�,�Gmp�xƃq��|��j��N��:��n�q�'q!E��eav.x�Vn.GI_v�K�� 
���BN�2�Z	�3�L �G���/a�C�ǈ��s�4��!��7"���Xl��T����D�D]ݐ��ɜ������-Oi~j�q��aÚ�U�]R2ѩ�gE���;�U�$��\��t�Ω�N�`A�靴�حV�W{^Ȇ����#R��K;�C����| L���@UÔ3y�����+c���3����T_h�
�Rq�r�[L��[y�<N��2D�cK�� i�5P��F�E��%I����}(GF;��B����Lbρ�,:���1��4[�kmd�ơG$AR߸F��PY�ޜD}���� )-�� sٯ�@$��"129CCaS]��3K�P�G^n|#
!{��e���?�@����փ��C���� �i��a7�<(Ld�g���5)@>2�e��9"�ZXB��f��tWXn�K�dH��z2��M��8#� ���]X�D��2�up%x2"B��7���N���M�;���Ȉ=tt��1|JO�W�5����̴�+������	JY!ї����XIA��Gyp������ɬ0�u�0�%�R��_i{��Z����0��9n�\�/����&L����=!�YH�D�d�Yߜ WA�e�N�e��X �Q@C�V��.nF��o�ց�[��a!^W-�t9p�g�}�4�:�U���N07D�b�ɿĜ=�9a��0����>WIml�0	�[]{<�>��y3�ףפ�p�M;T�e��^�_������/#Ʊ�ah���V�-)2��^W�xb&A ��py;<�%1����O��d�<�ӽ�4����k�Up�Z�9�@�K���e��7���F��7����p�to��C/���}�6�<W�]�R]Iok#8_��F3��;���\B�\Y+KR��"pXU]�
��է������h�V�5!�J|��s��]��I�r�3�:m��8���8�'D0�-�5`�� ��L,�����q�$e��l�	,RטL�u�X����o�g��u����R}��;,|�􋻏c�� �]k��W�K��ڭB~�c�ʷK��B���$г�b��ܕ=T��ح�1��%����Eׅ��;r���%&)k���x�y��:X��,��X��)�&�}��6�z�"��C
N��c��m,�-��ӤZgiS�� z��t����x~�McQ���'=���k��s�N���dK���b�D�[�E�fPff��=A�<u�{�r�S����n���9��.�"�Vk�1�����7At���& ]E,����[[��� !H@,�%�I>�i\�S�j�O����b�'a1r��#%<O[�Ͳ�?u�$�\"=ʬ��+�����<FVQ�c�d��N�5��j����4@>�s��k��׎�!0��І5�B��ާ��-7����=��� ఼BH��S����NU��&�29o
z�f���jZ0z����=@Ɨ«-�0�=;�{Fv^P����X�:ʮ�"�B<s�e�xj��&��F�a*�4�~���b�],�;�����b;��W}]2O@�H=�W�鸃��k��&[�����"!�=��r���~��'�?�Q�ݞb��Vl1���~��X��j
u�����;5�E`��C�sm$�5h@���Mγ{��7[a{\�l Bץ��UA]�Nv�OaU���)�>$�%��XE(ЗK��^Fw�4��xYq �J�pb��4�l��:Ǹ�O�ʭ��aN��#��갿�����Z��-��_b:�t��V���@���.�pE���6�^���d�ߔ��B �pK�鮥�����-�W��Z�QE�������,MN��5��x�`����
�Y��_�����kB=i���E)R,\n���=!\-Vco9 W��k��_��+�=�+s��{�J�4���'�Gdϔ!��ycAx�v�iQǥ�_�j)��:t�m̲��J�T,�`����~YBǠ>Lcd�w�Av�~b�л�����D?C��[��A�i`v͚���Z��T.���6(:AMp��")�?��0��DѴФ�ޡ�^;�.�w�Ԉ	�����F�ݠ�3Z_���h.�`��Cx+�C���T��������ȉ0"���s�us79��A.���M�o��'P�Ȧ2b�����WP�U�&�!]I)gd#�ґO��)x`+H:=6��+g�wc��G�l{�!JB�� ��\��x,|}�^N3���@�*^K��fS���ݪ�!�wmo��Q�3��l���>�6� �����Ο�OO;���<�5v�	�Zv�+�ݖ��;3D =�.'��Jk�ʽGz|���I>�����gČA�ո%���m���7+��[}Z8�/���8�5�20��R�f�s;y?+�!��vM.3Q�Bk�f��ג���\wCllHQ�Z#�D/�DND}}�=M���������h�*�ױʵ����l�3$�vf���Ngz+9�\Ț�V�֙&3Ù��e�����e�9�@����$(4R��Mv�ͯ;�$`l��i��j�K)���*��¾f˺�#�����Ç/^�푑�z<׃9�6�d-tX��nx�15�%7ͼ�i�,�ƅw�ϡ���]�$��'C�'���8�x�x���T���p?�%��S�g�>�4xT^,�!^M|���"trhR%����cw�R�UʛR7���A�$��5��������	��%�� U���D�"µ�yp�'T�	�7�g��0���j��a���$-��3*�^�tق}���	���#/����B��Nl�D��
�^ų2����8�j�����t���2\��^ S�/�?�����;1VK��3
ֺY�E��T�7� �c(4K���gWv��e1cWL7p��[��W��3!T�jY��.f���{M��6:��
׋^�x�j%��J������S�F��b����F�'X�c<	�jȬ�|D�4M(b�-Dy�̗,u~O!�D����j���j�:v�oZ1Q���R�t�jx�c�������� ��v`{Z&B0`)�Ɲ8V���-Le��Vd� ̾9PMPb��_ 0��(�5����U��%|�zO�7LD���Z�*�|Ul7��h?^5D  ۯ�P�E����i��N�7���v����&� ��F��f�I0����V4��g����fD _Cr�#�-�ٽF�8�ￛ4)W@��:n�о�Λ�O��]�+g�.���������z��$HT	�9�
K��>�^d�"���mp;4b0��UCf��Wv����)�L=�̋��[�����z�z�$���'p�Z�6�H�X?�d�5��u�.s�(b�ѡ(\'yE�$���؅ѡ���u����.��oY잒2=W�|+�M0Q�hy�G���ԉ,�6�~��K����\���'�n�n�!~?��cK�Sϧ���h�1�g�+��F.o+��kkӶ���1�.���b�3 �H�H�Y:k���`Y�ƴ[~=(������t�۟`���\��!xNzU\U��ک�9���y�w	}���z�ʸg�;��c����_�:��q�L׊��>���ދZ�:�J�.:��UX���G�#|����[S���Y(@��X7�8�Q��0]�3���r�lA �;
.Q�<�U��1���3@Ϥj,�e���;��J�����<{O�w,A��)���1��`������#|�9��n�o^��cgU�;����ᷧ+}���J�W;�RC7���M����О�'�@��̣�pF�w-��w�IW�o�{��w��r�or�Cn����j�~G_@�~���%$qI�Db�X�=��뤔/<i[�,�h��u⏔L}��^�ɠa��m���� �=�������yh��>r�L5쿴�7��=	Z��  P���>���/z��O�Q_���;h(�H�4������U�鶒����@�����>�$��[���*+s/�3w�o x����JzWt���`�l\�>r�I���V��پ�mcH�-i�D}��4�7%�\4nS0R�
�eC����w(7������0��*;�g.M������
���'�<�E4�E�d2&�Z7�bF�a˟�yf��vm��"���������]_W �( Uݓ="~�����g���T�J�����ԧ���N^����"����R�#Η�G��4��]���V	�P8��=ٟ4���E� K��T�Sx@��H���1,��t����_|]���18� ���~��O���ε���� �Wƥv�7��O&�(�T�~S�(��E�.���/�r��ħݻr�W)ױ�������-h(�*9f�	4[Se��4b�T��y�b�_��4��8����@���9�oQm5�1��]�ip
5�~��ԙ���5���6�Y^׹�`otV`+�Z����Xs��[2�7�y&k׻U��7�Kc*7�e+'������8A�eO ��haQ3^e���U�e���`?Tv�V�t�\��m^��d�����܂
AЫ�=l��q�0��h�W/::���D3�,����/���0�=Z7��Ъ�/��<Cˡs�c���$h���i�m��=��5�QD��4[ w�2���r<rj�"q�;��F,�t��M���狃����.�xH͒��<\����(�C[7N:(�7- ���ݮ8'Z�aC~{�~��L�(�h!o�\���e�XQ`m"){�\ő�ﯫ>װJ$�	�Q�g��M��IcXא�9�8�����bg��N��6+��dq�&�����m��&`n�A���8�P쮔�V�B9=�&!������-�b���X���]#_����o,��͢���3�1�u�k,7_��Av$��`q����|q�s�y���&$�l��Q���@�����*Ml
�icA?����,<⡱��树�ҝ��)��B�_S\6�!:ke@���A��ҁqTEj|s�`K��Vʀ
����(]zi���T�T�׽��- c� �H��K��!� ���70���:P���jċւ�L�/1����:0F�y��msRdW��7�m�{^��}֠�nX��i�<�v��r��vP��}�p��S�F f����Me�؄���0.��Ę��x��!w��5�j�`���9�!1�X����h�gr^wҧU�#N��u7�9�9:�@#(4}�e5B�Ǟ*G�(�b���?Day�x_nΣ�)}����G�zl�'��M`�3>�؃\��kZU�Hv�c�D�~�Inc)�����(6���A�$�Q<�7C�E�E�6+kON؎U�����σ������7�D����3^ �ώ�����o�g�~T ���&Nj��$�hE	 @U��U�9�V|��̩��c�6�&=���ek��Â���H"`��#���:.�`Bl�(E������+�	��m��,&i��*""���K����yn��\�@�Y�oצɛve�Y�7�۾�~��KηǴ'�N(��6���7ȇ%ٟ�7�9C�_u{ˈ�yB�ї��vi*K�;�H��L�s�1M+l�%����X��$'�W��uϻ�fap$ڵ�qN�29!�)T��7i�"}�>��昪
��~�o�*C.�^d	�"���=��p��iZ�|X�V�� �2���M�@���wK������Z�wt�۫P�������
��g�P
�Pa�)��00pv7P0?�Y-"8���	<��S ���,�Y}�U
XoY{���$��7䠭��0,L�$�uב�l����V��n@���.a=�|D $�{g?�|j��y8oGM �|���S�X�}3�ssO�ʻ�]�Cc���I���<��������M�є�;Jd2{��/0��Xq�2IGo�._���x���Av�5�?��SG'���� �J�J��O��������A���{�e	�c�:f&`L�p_ʉ�{:#0�`�ψ���̙f�Ibħ~�>y�wF%��D�l�1�Ǥ`Z���ǁ$4�|�ooZ�¦(�z���G���'W�s�+Xy�H7l	I���[�+f�C_�k|��e���4x`Wx[����!�W�%>&�$�d�(θ3�F�(il�'���&���)L��[A��p��!v��Z�m>zzN1ܲ�}7��
Zp��|�B����e��͆�áir���o���K��k�I�'����s�����r�5�eX]�$!�g�R�R��ņ�gt4d��)�S��%�8VS�,�&�9�+���T�U��f�>�|��y���� ��������`�SC��/����zp�����M����j�{@���,zC�eW���P*���([J.���!��J5��K�*t|�j�k���=4=�8�-�ǘA��v6��=��ȳo�R,�u4BT�-@'�#B�^g6����GK���
O>UD����]43�Ԟ!&��F�@����������|�����	�u�C��o1| 2��������5��?Jk
�su��
9^ZB� �0��.><�ѯ�%Cb�vPH�Sڗ�Ã((Ba-�6� p�q�����ٹUv���_�[��I��Yf��.4�ӏ��ĥ��{ʤ��\V�-�Ų&_��-<�}>'��ZS�"�hA<9�M��N>�2zLHy!z��G��k��H~!���Ids$�[.Rg�r�!��N��Ѹ�"n|��[�zy�-h�s��� ( �<�4��?�sZo�0'�܎�|�JeG�r0 ��g�{n��y[�u<W[6#���L��yd8��e�Rnt��;��v��dRB��~IMY�)�ép�����.�m�E��s��y�w���&�7+-�rN>W�è����낃�����T�����\:�� �)?7�h��yO��.���T �$I2g��T���Txk��Ǽ��i��VU���X�;?�l��=H^�f��&(�_��)V�mt�3o��!>�=�w8T]Z��/��S:åB�=�>Y��:��Y3�7�����0[��"��5��̄�e����[��YM4��&����La1)��J��e�'ZJ޲
E��p��O���E��(auNٔ)�N�P���:�(g���$�)عM�g�:��W��}͜d\u"}t��N�N��I�kDb���L�]��*�pGT �E�S�}�F1�%E
�﷍�D+�p���hc�����.��oƮ��E��j��E�:�v"^L�ݡ_��� n�_��uY|�y*`�{�M��h\,m�D���k���9a&-C7���:n���=UvbN/�`8�ڥ�����ׄ]�$Ò �3�s0��sO	m�+T�`�Y�ɤ�+m�r/�i¥F��w��%Lcf�˛� �%%+ �F.v􈢳P�vH�V���fL����r��v�cJ=kh�CN��n��<b�~����KP���m���$�R�.G��h_�����@����%���m+�<v<N�xЛ��+��#��Z�x��b(��A2|;am6"�m��}v3�Q�?0�3/?�A�1�8�����K���8�©��
����e@�u\����
iY?�<.�b�~����+qHp�iX��h�<�천`ظ��g���q�����P���$ǽ;�g|l�5X*ׅ.�7��^rO�m�̵|�1�c��l���Dُ}�VgMJ��1=8�G�nNm�q�A���ysB��)l�H��]O�j���P���h��8��s@�?O�/<,Fm��& ,�:�i�X2�����\�$kkȷ���	G�0D�H���t��e+��D��眭�WD6����*�eKT{��%���I�:�Q���R�h�Ke�����T2�v�~��ψ���H�~ݼ���;�
�y!L����:x��������-��~���5,��OYy��oe�JY�uG����=��R��V��c|h*�55���o�x��n�X����|���؟z�
ȍ�T�=�*1BP���t�A3������D`+�U�hE�Ϡ ]8S��<-L09'<��ȿ ��~<�!��iȪ-�e�z���с/�� ����\�O9�i���z�,ł5_��\�-�u�%��������_�8�!�L��:Q�ZA�ġU)\T�"6����M�>��93�j��Rj��U��e�jK� l)�DZހ\[�-��%(9D�_�nu��n�^�T/u�����f$0�,d�A<W2��yL�	̱UJ����=*WZ�Y_GgXi�v��`���b3M��H��!���hd��`���KR5" ����V#�M`<Xc%yq�G��w��m�����o�b) �ҳ����S x�b2�/���<Cc7B�^e�B�����߂=فW�O��h��FQ2�u���L?�|�_	\-@��^0���Q%KJ;H֪�m�	���
%G��dIU����]*P�i��� ���h�7���+rU�Vg!j�����>zc0��8x��"��\J�c�;=��V����#XB�[Ւ�-{&�� %�
a��Kng���5� �9�Y�2M���%�>]� �6jcD��1��C!�@��#
lm�D>I~ 3�]aUz3I�y�X#D$��L%�m���tAߐ+C<���+�xs���p�z�ah��)���%�Z@'�l��~ϛId������� z�+ 
h0�7ֹy@�(��y2؏�u�x��!�L�	>�Np=����z4sswC!0��z��q�db�� ��ʱ�z�uf��̐C� �q����s)gm���3����0��諰�m�y�y��*�M���� A��+��J���%��c�c����-ұ� ꪷ��n��P��pc�՟0-Mw�h��8�*�"�L�F��/l����]a�����\+����?!5�f��Պ�e�N#d;Ҭ��`� @7���� ���3Kr=ܱAw_�X{����z �|.�6#��\[h�Գ��&�p��.}�?�C���t�NzHk��D�� ��=�	�{>�pi��O"��A�L�8-6>W �]o��������!�ù_���e�����U�f��O�"��Wm@@J��kmIz�x*���D*T��J�'nOo�a���y����U�H8���E.������8jF�(.vG���Ǥ08��X��ǁ���M���S�!���J��*��f��E�J���x%��>�zY��7e p�RFܻIr�<z ��s�!8ّ�8 Y���0B=�x���gFX����ՐI�w�ӹ��c�ͺ�"XҐ�̝�;����۟�Eut��`"Y���0Hy,I�`z����Z]�`ri	
�MGŋ��������'��~u�a6���BP���Z��D�nM�l6��'��׼�r
�m�a{�$_2� �<� ��b�4Wj=�7��{%����ȏ����B��)�����t¬XF}w���懲�Wt��%�r1Z��`��G�fSw$)�uj��>f�h�ׯ�v[U����a=o���Y��A�����P2�8�W�@=Rk|P2��0k�&���y�mǝ�;��Z]h��E�~w
'U�S���V���m�d���;$%x��#A(8�W��Bw뙬���Z&�DjK��-<uC�`�'` Vl����:Ӕ����6���Y�k�,u\��j��)�˶�����R���<HK�j�����[��,elV��L���K���:��}b���<�rG} �~tnNZ�l��/p�)8D�O��9Kz�a��+�(��c�׋�Ec�e�d��G;n5��>[.�F�9�������j��q���pD�ѡ�=�7��4�Om$�!���ʟG���[D~\�,���Wqz��9�݇����g<�6<k^���C<��*����6��2��0+"!���vI؇���1�ڏ�I�R~~�ߵ�-uc�/����# 
�	�oD�bo�5v�(����7��r�t�ٺ�:�)�F�8�ds]���?�g������auʫ�������7�~r³��Ú��,ןz�+�k�?x7�pC5{�p�4qJ�	��Wn�JYu�NU:��=��c@�,�H0��8��ǘqd`6�?T�x�D�0��ns��*:?�S]QT^I�D�%�>�v�&�s��U��� ���x.�����d-߈b�
���p|Z`����0i��/1D���%_��عL����`d��a���W����0�ᵲ��1��p^�i��O�R�;,��<��F1n��7�>���@v̌~�xg�n�`�
`����n�beĉm;qi�Jc�*T�W� �b2EHٙ��Ւc�婁7L��RY�ֹi����2���f@��0�{���&�_�<磁�J�cu+�P~x�x�VX����m�wI9�I�_�89��Ҧ�GW�.��jyk��H$\e������Ú���a�`d�?V���&�r��l>��������Q{Q=��^�ʝ�[���>�k�"��=1F=����n�NFy 4�K8C^g����JdzJ��� �خ�������w�Z����\Q�_[IV�$����;��"V�r���S�����<���{��A3Л�j ����PW�[��A��J>�4=��� �1�c|�9-�uLJ�G�5�J5ܶO�C��yU{Eډ[���w�'ɋ�]0����ǹ8��7��[���=&{I�Ge�����L�B��:�>��L�(<�MI&ia�B%�*�M�3�}�p���sx�b�	:8z�*(!%�k:�&��m��[������!��Wo�C����k�!�c����C�'�[���
�Q��H�M�o^�ҏ���|u\�0(ꢹ��$���=h��7�U��������c�4�A���Q�����A�>^=�
BU�01���82�rOlj���gbe��68��)lZ��L��\$��P�,*�DIObU�+|6^���"��!�rqU��'�ֆw��9;[T���T��4�/�K9��гc��C���MWnWA�MV�
h&#�7����bz.Dc� #�v����0K��Ѕ� Pg�U`h-�?�⩑; hI�7����/���
���;��[O���bW⣤ԗ���v_}"�W�`Ez��`�t͘���iɓ�K�Q=$s�Γ�O��� �&�{<zw9bnt����֥c+Xk��j�^|H�V/�zn��억�� ���8h�iދz�P�GePs��r�/��nb� ��G�����'yۦ�|`����Ǫo?�7�4��o鲙����P���$�%���s���AK����K�>.R����յw�� !/�m���*��4�'��,�9���Mβ��eC��;(�D����JM~$q�G<����ˆ�,.���s�SR���1���U����;�@Hs�"nX�ӏ�T�oZU��R��d�-ͬl�w�|_3��K�|%Ȁ���HU�U'�����î*}۲���V�<� W��F�l�6��n�d0m$_�X[q����c��=_���R�3��E_V�ʧw�q+���38�r}�_��
���8_W�~�������ꉭ��@�t�T��N��B#Q�$nP��ug�@�
t��'�l;�a8}��TN$�lS����>��]ڶl3xC����毀��I[N�%��O��B$�:��?/����{La�Te�kw��}�o���y�Q�2x��8����R������Q��)�XG/nTGKQ�ი���kZ<�Ğ���>_��WL�W�>&^-�I����� ��a��IY���Ru�<J�7h�=)(_m�h�/1������ixcz8 ��b<�A�)�L����yZ$���Y~HƑ����;���צ�|d-�̿�U�}V�'�F���R|�7)	�C�W`����>"V��=\�k'M��\K�f�?�J�̶� �2����YHs�*���r���K�x ��[5]��A�%]�
]@��Uڃ#�ݿ'�4a��ks֎R/}4ޭr;郮55�Q*Μ�ޜ+�߬��/H6�ܤl�}��b�G�~s�c�
�&P�IuN3[�R����є&^���[��	�R>���,�-�����71���"ţ~g��X=�zP3���`�^l���V�G�� �#0�t'��$+xTt<*��G��W�vع��;Y�nh[	$p�2 T��؈8���7f�dq���d$�cAb�,yz��V��������<�)�l�Θ���1� ����<�R�Ӊ��q#�.hG�Ԇ@Ȣ�)�[-h��'�[��2H�u�h�<�,��&N���C�:�0l��G77X��}y����DN���{��1��^ܲwշn%��8�I�z���U��i���Fn�. ��Na'���Y�7�/�N�^O�R��,�x��E-��в��Gy��_O�YK�P����b��ر�~:Ѫ����R3CA�/ �!>�K��3��Z�I WYg�>!�'��ֹ�@h���pw����q9_E�+/oi]��D�Ze�6���>�rM7���g�h�i>P�%�����ta�% �I�Ni��͜vZ�"�Q����(�:�{��A6�k#�F�����M{<s�H��OV%~TY��?��)H6������if��t���)� ��=��aM�{�x����N����%������P�B��=�{��8@�E�E1޴�H\����Ɨ��]Z���<�KAa-��,r�폒��05s`ך�ܧ��݌���]�h������O�[�&���-�f�]
^����":�3
�L���g8[}�GM���.k[ۺ�s|H��� � )���f�RV�[�*p�MjF�: �������3忥��LJ��6�{��`Ye�zG���KK�_/g� Ҷ�j�A|��7y�3VҶx_C�wէ�Ҵ�T���G��j����s�?Ho^EQQ�AecU���aa\�q �߾�����|�Kq�y�r�-љ��"
�`���ǃ�++J�v8Bluj'���-V�'C��}Ԏ�,��A���d�V�c�ɯ!�!�&�Ƀj�sA`};��UAE��	ەX+_�K�J-���gY�U�ȻT�Q�tW�?�B\_�U��-�*��闌��H�۵v*o��f�HN��:�6��&-*��������-c:q7��e*��129����I�l���M�����7�&�`�h��r�ɸ�`�m�m�1���uo��l9�vٰY����vh�/1rʛ��#rR�]ސ���Lԙ�X��ֺ�kB�A�<A��q�tPz��a}�XJ��U([a�7�a8,����/��k�-� �7���4^����N�peF��)�B�o7(od�6��0���W����4O��&]ܪ;"=�T|f�h��r����&��t��d�|k,�W*UAeL�YJ�s��#����2aJ6ЬTT`�Q��.he1yARR\�n�k���#�ŵ��h���=`�z丽9�y�ל��v����b���Zt!��(*��|^��d����-��ń[EU��d�5��[��M���۸�45-��u-W3���_`[m���$8��Ĕ�U����x�x��o���E��bnm=��#���萹�Ѳ@����#}/��K��?��"����UC�{��7�۔5���p�q Ɠ֎=� MF��E�:�(3e�$�V�^F��vӊ�s���� � s*藘=O�0(5`�皶a��1#�nE���b�\d]�{}_9`����4�M6����s��Y�Qc�mJ�WP?#�&��E*��9P�ᯑ6�Y�=Fy�^�A�5�h��y���=rtDSu��W���1L�ڢ�-�>����)�`��/��\[�\`��݇Ҟ�ڙ+��;08F5�o2�0��7�0��S�lT(O<�`�����`��Ԝ@B\Fd�J$/FJ��]���ɭۜ�|M��.��-0��q�2�kX�؂��#Q����˻qNh�;��țs��2�~�t7*�|��,A-\�N3boƉx�^s���j��k3�Q��[�Pr����ݭ�d�4t�����1TI��Z�p�Ǽp�Wǋ3؈o�SWBgFP/X�����ϋ��-\=m��~��X'�lXi��F���&��3O��O\��`&�
8p �F��*�JC�^g!k%hHMv�������k�k�*��Q�z2���~>�̅D}�h��>S���݂b�d�g݂l��'�e�^�1~f����3�y��+�즽�b��օB�ӻ�BE�'W�'�ZTo�D�|$�dV��(��խ
�W��.�L���C�8�,�R�B�z�_�-~���tm@���j-̪��&�i>śX���e%<MgT��߁.0��W�G�F;�n�Ů���W��<Nݪx�K�%*��Z�_NB�����_��%���Vx�Õv�B<��[�B'ǣ�D0V���T�j����ܚ;f�˹�;�
��5����h�0��Q��e($��%D7Np��V�o��1�dG����lb�x9��Ϙ;���o�@�b�!8'wW�s#hm�sl/������h���Q=?�l4ĝ�"F��^	�KPB��(�ɿ�p�aۚe�w��8���b��f:J>͊�\?�䇿Df�*���P�(���)��~#���	��
��x�-B���?N"����2&yX�n��P*JE��Ԗ� "\uA}��o�q{����+\q�lԚ�|�>VNt)��/�LD�ˎ:��/�����GfG^
�j$EŹ��f���A��_cq}�	eg�I�@ {o��BE�<�0#fF��W,��DZ�m�/���2�6v�����+@	ܻ"��(R������]��O�2BҺ����Mf\�*%��P�:ʎQ
�o�e[�0E�?�M̒G�D���aNcC.M������%>R>'�ޭ�X���9IaS���O����bkau���9T3\	��2e�k^�\ț�洀��B�{�ff~_�h�zj%Ȯ�헣��AWp��A����������C�`^���W�	��q�z�8��ƞ�������:?�)r��κ5B�v�AQ��݂�]1ߞO]'�L�#�IΞ��������HYo��l�E?
�����ѓO�����S�w��?��t����� E�m}'�r�	B�����NGh� lx���Y>,a�6mi���f��4ՔS�[���ɒ��P�����!��H���+�GAr��������W����[k0�W�g�Vw�=�\L5����H%�چtz.�����}�9"
VTtܒ��P0Y�`�̀�����\��xd��(lHM1�H��`����?��脑E�h�pёQoU�+�l�G?�7���4�����FVK��ea� �R�]'��'�U�0a�*�UPZõ"��zҕt����֨p�_Q�x�
��%L�*2�a��-��Ch��\9�����ۦ�QM���.�71x���\��z�/I�(/�'�	fZ
�,��K���� ��c�x�^��v�$K���B>�ҁZ�vO�n�A�+vV0;z���Q1-f1�����iWqM'�\��7=0��$����C�6���1'"�ݍC���r1k�y�N��C�9ȥ��8�='�4޸+*&����ݟ�H�A9hpL��I,.��ړbc�d檻pS�8",�u���x�����䵻9T'2&8�mf���M&�<����C�"�B3G15�X��B��&<x�2#��ˌ�6UߠG��<����*d|X�!�e��;�ŝ������l�;z`�!w��]�s���se����s��W��E�?`0��J���`*��`�|�1o� ඙�����!��=plN݌�A*���V<�6a ��ސ�W�`�-\�ؑg���I���^���F�z��� �_�|Z��p��#��o�h@�w�`�ٌ�eY�N���".���x|.��+8�4T3=�[0���6E&�f��mB]o:Fa�jl�k�hM��]{�[����>\%6��O�R�B��^���6k�	Y��F�CJ'6�v�o͐�Rj�e=�|�;��	
�&���� bҗ��� �{2Qf��`�!��%�KvѴ��l.����=����@$|��G/��y�s�6�ـ���/!D�a�X��� ��i�^�sv(n9�M:��7��_B�'~� �L�.�e@,�hh��LI(���_��|^[ʧ؋/����,$�"Z ���pv����gP�j��No�1�!�1��m'	B���	�6B�0�I�����I�$FZ��H�0������N�헚��]^��ѕ��>�怳vf��D������~���1�ޗ
M�؍K��z���=LQy�����^5�ꑅ-}���H��Z �m��E��Y��zopS=��]`N�ow?��g���`<����Tw�&y���7&g���A=��D�;��#�����_\�z�
��k�͸g�1^`BU�O|��9r�z�oA�M�;��3����ȧ��􁏳�D5���u���vpy��9É��Y����ta2;��v�,��%�ɃV�j��%
/��¸��� �w8W��� ��i��JVn	�ԁrR�� ��j��sh�8���vFŻ�%&��d�8���8�G�O��d�b�2c�/8"��S�h���:�P3�hٱ�(��!a���
'o�`�uO�;����]��}6"
C�+}*i�jk'��A�!�RG[��Ŏ��#�� ��${tP��]\��zsgG�0���.��+w$�f�H���j��5��\��T@�"�l.7�������n*�_U���j�5[�����#��+�Gr��щ~�3��C ��|�jV��D�ӤX!�mQ�6E2d�����Ck�mY߸Q�rjH�j��¶׍�	G��:6�d��2��J�r�Q3J$p���BK<;F�-��~n�,ҙ���;�g6e����#v"�{��G�C���(�1Y�I�
�,�N`� ݢ�����C�C�7;O;��ɰ�1��ϷX�˻�a>�0���E�|E� ş�dt�=dKC���&�f_�2X���8a[�D��������d/�ݒ��YzmΪ�7I�d�S���v�`6Q�y�������b�b�D�(�`����|C�t�����[�E�l J��e ,WM�c�E��~*r���Gt���%Ŵ����u�㭬��V�F��:b	�o���ixoϜ�_�K[�C��b�NT%�I �lQ�#a��.�SY��o⇿�T��]+Q-��������
���μj�	Fϛ٫6�;��4�c�ҤŪi��&M��R�������6���I�:���[�r�#5�����@������/��]e���7K�����D��,�N��<�ߧ������F��v"��6�/	*|�d�U��c��ٳ�k59K�M49��L�~b�l_h���o�.ȁQ\yA��dWuՇެ����c������r��}��c.r�eF�*����Ie#���ƻ+~^ʡ���8m��N�?��הwՕ�s4R��Oi�b!�%n�� �����m�2��Z73���c88�X��k����l/G�������ЩLUŭ�mq+X�����>���P�Hr��Bf~����P��V$�������f�<�^�Y�xI;�kQ��rߎ�R�ON��t�0������uF�D��0<�ʱ�<¿�i.y�X(cФwY�O�F\�Q'h1'>���KeL��w����x������0���|:��@���A��}��㫩m��F>���:�ҞF"�B�Z�Q�z7��8r=jʘ}�C�GfnXL��=���l D�p��S��A�d��e�����F�pu߉W��:ǆ0�3;���'��~�9)�܊������T�p�W�ɳ�XH�U�<�/Ւ!]�.N�l�	P���L�q�ؔ.8�c}��H��8���26P��;�hQ���p��v)v�����?S��A�ri�]�40� �� VrW>c����@��g�_�:��9�˿�_� �S҄���)���ޤ�WhB�� 7�R��~=X	�z�_�"�?���kEZg��a�Qۘ}�M
��F�	,W�m�_�����jV����B��s䕱�:���*qX�AM�f���D�|N��f[0rT�� 'F❰����5g* }P�+J�d�
�&+��ex�A�ւ�����1R���̙IH�*���bF4��P�QE�v�(�iw' `g�/+��0VT8���r �R����dq�+��10@`fe�`1����%+m�c��������I���dM�nihj:��i+�OMQ�+��V������Q�uĩ���!/-��I�FG(T!t)n��͠�!�̨N���s~!�p�+��b��y���Ef��|m6?�T��f��w�����)�{Cj�����ɜ	��{�Vj����*�g4�6�3:�`W K�����>�?s�
�x�~��	�wY�g��j����@�����Ea��|wRk��AQ	Y�)��2��Q�4�t[1��p9���]U�lvM�`$\�$��U�\�
��������R���<�����u��K2��L�w����&]|���,�'�w4vcƜ�1�VO�3��+��#��؊��4�FP�n�0
�j�������I�,E��>D6�j�����<6�M�j�s������CT�wｩ���J�Ŭ� B���R�@r�!����[�&k"I[�v�44�IV�+ҳ�*��y���Yr��� ����]w��x�*o�p��	w��$-����ǐ��W`����ct�u�!�����@���A$жH�=0}YS�Q������S�G���:��j�{�&����*	�O���$��,�^��ҡ��Rl��~����,ԋÌf,;1�D�n��ih�~�9ГZہes^]T�('�#��7��R�e�>�c������Z��@����Iý�$H��.�f� �c���%C�c5eF�A�e�
�B��s��ҍ���̢���*
��i\�ӑg�2�d`Ƀ�֠*���;��\�
*�@t����+�z�����p�f��ة���^	fN�C�X'G�X}��q0�VG�-�h"�M�������Ţ^�� V8��Ჿ������
�����@��d�$bۡ�qQ�+Kur�����~_p�Rr���j�k@���*�CfDd��~�J"|�4M�������o�^� �d��`V����V���ˮ�����3\)׵ �HO��/Y�+���>�b-Q�}�!�Bg�+�K��v8f����9���Ux^kq��$6�M`���0�M=%���˧��xZ~7��X�
��w�a���� �
Pj�jJ���rI����V����=��3�:>Ҫө�K�43�,��iำHۮ��;��|��7�87�+X�9�Ã�>��w��F����h�x�*"MmG�KyB>u+�e�c�Kd�4�WV��c�l�kBGP�c�^į�7���M������\R^���}�	��nm� R?y*?�|Ul�2�����!� C�i���e*�%���	��#�Io�B�n��h�D���no�����٠Q��@���0�&I�^��	[`�"��[��<�~Tn\�Tg9��%�S�xiR�k
�
���r���Sk�s"�ZD�]����}r蔙!ż{��3ّ��Z�{����'H/S	���\/���L8����ʚi��]��ʍA���S�W�G�s
`�F�Q�hT:��p��p����$]�w���JI�L���@�<>���p��l��'��+m�9%�@�!)�2��u���.�����@."b�]��z��ҍ��ʀ���G�
f质��ʨ�*{O�8�˷������]UoS�2B1�] Q���x?%f)	�
F�Ň�?����~{Y������̓a[_*5�,�|�ߐD��O�I9p2L�m.z ��U��aJ�Ñ�	-@$�Զ&��}>I�B�uy�I�?�-n�wBd5��>/3'��A��3��4w��Sf����=��D#�F$(f�ӈa�IŴOL.�I=���I�(�����%
�R���]dt���"��~��E����Vy!-�U���mt�ۀ�-:�e�(�W7���������&N��lhNVT�RB�t��՚�x�$���-���R���S*Z��l�H���F"lH���à��+aP���7(���Ex4�4�S�dy����w������ S���`FT�o���>Q��T��������'���b[jr��Z��s>ycO������T�Ɏ�o�U.�£��"%F��il�!�����L9�`�z��HR�9�L����/v��bu]|�ų�D$x��/Mw�^�����C�E@M�ӱ/ݼ2������Ex5��ǔPĩ�M�4{a��5�����z�v���E�EB��a�B��J��p�	�Zx��,"���0���{�oB�R_Kʃ)�� �����r����gH`a#�&��5�ǖ�2G�l�.QCߴ%4êwqY�� j�%�P�Y"��B�PL���Z�ńD��)+׶�ϐFzi�������J�1IQ�U� ��ف��PV�R��E�}��j'�}��a\S�!P0�Y��["XL�+T�^���-�@	H��ə���o���kF/��eBm	�Y!��lB�G<X��VR�e�X�� d���w�h� �5��h[q�p&�˙-�?���V,Q�Ȯ��L�_8�"�@R������ӷ��Y��dN_DW����vs�w_g],a��Ɔ[�5�n� �\� d3n!ҫ�7�ڊS���qx5��~��h���B������#��z�x,J�7�,Kvy�}��ffY�_t�}�}R=��D=хJ��M!K�#���Ҿ�hv�֬ɳ��iA,�uF�)��~7��v���Q�ST�{�ges��c��:dK�h6�ϔ��h-�8����!џ��\�O��
#]9mCG\A�
��ؠ���I��G��<���$N! J?	y�Dr��꿽��|m
K�ʑ�|�"g �!�l�N|����"�Oڦ�������D�nz
!̂-h��B&�09?��TP9�ժ,|�j��n
��1T5�H�oc�rZU�-�ok�̽tϴ=�8a5�Hf�_Lꤜ$�U
l�<�B�}`u��:�cߋ|QM����sl7����Z�y���� >�t��,Q��\M75F�Ȉ�R��l���DOE0	�!�i�J9=q ���+�i���j�e�ftT���ހ�\9�*~�Q05�*!��MHeWyUi����R=�q�+4@5;� ?����?�@�p���=4�A~�m��]QK>[J��f�D��#���e%�À
����B=�������	��V�[�,��$��V#$������C7�Y�!��G������ʷ��A����hv:K�?��͇�*��s�ͻ���?��`y���w����f��+�E�Z-�|�5�w%|q%�grS8��n��A�N����χX���UkZ�}7?8����
�V��J����9�&��K��|S�%6}�l�ZeX�ax���aO��hBb.���L����Ȉ���4`�8�tQC�� �D���?>����S_C�B:Xb�N3����6@�*�gu�*�pE'^E�O�i�B����N��]L#��l��jS6j³�;-�C	J�Է�ﭭ��դ��B?��{6��ܺp��oٹV��Qd5�*�!�*\�[�UL��o�=�g������L�����jT;�+��"y�_�i��5�4N�2��Y̯���DQqI$��w���35�"zY	(ٷ�FT���B��0JfZ(Q+sF�ôN���J�����X�W��\#^H��e����C�{�D�=!>z��0-%b�1���*���e�|��t!�ι����n/V�U�u�F����l�X��Hp,�����;(���^��$�S���jj��V�K�t�%+��^��/���}�Қپ�Ȯ����)�i�G�'�:�=s��2$��͗��1ay�:��7IH.��r ix�}��PkF�-/�o�j������@�S�\NO��4r�-w��B:REK���|y7�u�t�e)gW��u�p�b�E��J���rՉD��Zt|Jw� ���5�\|)�rN8��.weWm2���9(�*q*Ƣ�K{��&�i�����a]�����1&�-\N��F����g}�ߊP�o�F�<�^�W<���n��S��5��5�.�$��D�<ؾ���8j�֣���0?Jh���Wo�$���9��/U'"��d����#�ÿ)�c5wz/���e���*	��D��M���gtb�s*��U�50��agR+S�3�R5�hu�P�rF�7�f���V��Q8]��b"����@}I֪��r����"�j�q:Ȭj�̡�ߴ��QN��4,��:0�HE| qG=Q�-G��ع��"U.SI��m�2]�ׄ1:��[o߀O�EG�wPc��F�v[6����Oc��v�/[�Cۇ�O)A����RsL��!�E���w�l�?�N�?�y���E5k�����ё����x��;@�*G���[�\����:_�0�&�����<�<����yC�m?���Q��vG����b��@҈A��tЄ	^(��ؿ����$W�80�٬�`��L���t�Ku@�2Ը�\8�џ�da�I�V�)����4i���w��W�.�0�~D^ti_�>w!<31@�c]@-��{�2������D�[�t�sU7#=S&�uJ�3�;�!8�x�{��s��� �BDW�d'�؀��"����+T�w�Oڃ�]��' IV�\(��M��i��*t@
[�	�N��)�0-���;#�Y�o�/�U�9�<���<���O�r԰����az�]2�S�D��|�]���b��Y�>�+~/��"�d�+{�-�󞐷\	�R�}��kLn��Ͷ�'�{8����[�$u��ܸ����h���èu݂���ț?�"����8���O�j�ò�d$�0�~����[�sC�"Eɩ���I���� �l�l����
"�ċ�MB�w�ƥ{�����F�w\�aα�r�U���$��*՛M��.�s�_8CA��oAL��:z���i����@
٢���C����9��庚��_�a�CDrjF�-yOӋ��p����&���&��B �,p���Rt��"e<%s�߸\cT�xPu�S��hoG.�T�N�xcõ�����G��}�"}�w��oܡ=�zK��D�GP�O/fϟ�{e;��#}^�~�<�Ewt�ߡ�'�B�p^�i��s���3�$���6���Vd�lf�'td���c�r�ط��#�'��C�pc�#N�*g������M�����TzД;��ڒ~<�׽ā��}�@E��B_!�q
k���/��SըDwa \��B{n�v<�'�:<�c�i�����{��@dєv�녦~��U ѝ��-�w� �5��,69b�(q�A����ދG�T�x8?7�Ē�.��o��E"�J�]��/���:	^��,�(�[K��6�J����,���B�Q�i�r�10 Μ�C⮗@zʧ�)�tê6�#�_�9�L�X�iJk�t���d��ԓ��B@�W\o�g�9�:���.�%˂�#m��c�!�Qu]y�/�E�䔕竏������K{O��T�ߔ�f����:��<��g�h�v&���P2��V��~��g�-[��c"���(����w���w(���AJ�}���75�>0�lŰc�2�*&>��o���P�O�AO
�k��@�
� RC6ԡ#oW#Z� H��p��,�����s\���2Ku���Kk��tN�l;��X��W+��e�H����vG�� ��/���1\��k����*ʅ�-۞�� �)��	i�E���dc��i$}9�5��lulC�4n`�ʁ�Aih�2 -5���'�8pN)�|ೖ:;���5\��[�ԥ����5�&�b�"�Zj=����9V��"�O�U��Z#�V�ŕDvO�f�<�\i�����"ho��J�!=�ET(q�bL|�N_��r���l��^�B�60���>g��q�@�a�6�-�$���rr�h�, ��`4p+77d�}hҸ)~��_U]��E<P�j��u�<
� Q�vR���p%U�.�����0�CN�*�fG��ԅ����$�Bբ���{��!trȣ*����ҙ�����T��(p,.�?���5X��R�er����p�E���;ˏ�}5v�.��eB|�s; �]�'w\�x[m.
�