��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0����_���3e���ӌ,n���6�2�U�|Ma����x����u�uW3��&/.FU��������F�����E4�k�^��~!ʟ�e��A.ִ����,��ܑ���m���)
b0Ns�I��/]���2�q��RPq����)��vHv��	���4J��e���j���nƸ�&��?�GP+$����<����?eG��#g�� ��k5����J��Dh��4�U[R�l�&5&�}zX5�[��d�P����}-�&�0�O����W鲚���d�2��~���]���Ch�\=�[i+~��+�\��@Z7�b�'� d����"w
Ě�E4&��UIc����wO
@]1�|QV�>���,�ud�
���}F,�d#�r �D�*ܓ?J�.>���e34����5�̻��*5X���4�0q��@��-�
"�	sW�z{~�Q�G��'��F�/.�1YJ�O$OY�|�E`8�q���SL�h�A�oX]���a���6|��֋��:�L��}z$�Q|��'�o+H^6攘{��W��[�P�X���Q��`��L� �1�ߺ'��q\#D>Ў�r[v�M�,�х-h�T�{���*�T���C���,-P����[}i��~�ɾ��
A��e:��j�#����w+�e�|���i��6O��״2�H�Sd�]�v��>�f��jK��f�#���5�hzOvf�#�>�SGPb�d�QM�c��Ȳ�A�y�GC����9m����Q�X�:�	_��e%��bd�͊��+�z��F��c%{���w��ya1���R���z�|�z&YocX�P�nq�:���q?� Eq ��a T����mx�ն�c:A<X�������Yt��,U����?���>���{M��|'�*�`v�@�,F��U1�w0>�lHR����W���1�>���,yl@]t��BH�m_�sQ�oEX��/}4�D�K\=m������oE��|y��kqo�m����$�Y[����^P��}��/~��e�3�OK/ߗ��<F.�sp&A�U�[y����H*���K��b0�ݷ������6,H�3��dC'�Ts`)�ek�[]ק�9�m���%�7�W:��,2��^ƞ�P�6]�@}�E��r�e�L�?�TVe_k��ԙ'On�kǙ�����g�x�5�mC�����vå�h�&V�E�dӦ��sqk�m����1�n+L�cg�+���Վa1��?�����l�FU��.x��M�5����������6śR��ק\4�Q�rTWx�D쎆�uH�)���!J��Nk��9��E(��P�Жs6��mM7G�i\n�/`ǳ!�u}���rLΧIGh�x(k1��o޽��Z�/:�Y�]�~v3w�ؾ�K�䁷�_;�;����VY8͔�Iu&&}Xe	��B0*��#��T�����lȺ揃�EB�1���
d�s<|�+���{�[	��m�7�.�eFޠ84
����R�S!@���G���zC�z���J�vR_��\�JNoJ?�	�#`�K���S��CA�S�4v,NfR\��H7���&��;NE	��묚E1�I�0-�(ۡ�Q�<�t"o�i�'�{F��T���}���,z�c�<�� ��Ǟ�FMwR>��Ϡ�<�L���.���C��X��5����ڱ��O�{C	��!D����~�XuQ������@��nT��@��w������-|@]n�ѝ$h��쮢�$�����~�5�+�+������4��S��[���8ÀE`]��
��>S�c��5Y�H�&�=�%E)rd���m��>`Rbws��L����T�c9 �yd�bɨG�LTj�?�A��S�	�d�f�L��Nϡ���_p-I��Ϲ��ؔ�d��C��ʌy�!¶�1��-�����B;Z���[i�}�z�g��Ͻ�����%��4�g�1ͦ�9ڑI@������^0y��(��D<t�B�^iF�9MUid�#�MT�Y�+Y&T~��0�d��rf�&�a)l���� �)�.exl�=�2~1>I|��\9.=���:)gDZՠ���d&��j<Cj����t]�F�*T�Ti�LE����Êl�tL5n�Yzؼ��C�	Eyy���Q��;`cZ�U���;
�GD���M�ny5��q�єn��>�!r/9��S����;�oی�}��]P���g�c�yU,	��AhZЎ������ ��-P��\P�������2�rJS�_�ϱ��yQ(� ���O ��o��2ðE�tRZ�_8�[ )`>�p9�7Z�^Ѧ��n] c�G9ߥ.�$v�$��M����\�W	Y�;�����4E���~ZF/q��*�;X�>�h���7�5��nX��45�vA?Ι�m�ll��Z���˗~X9�s]XS\�[s3�J�6�ndi/�V;���kz6�a��%�6r��st��{���E�tpߋNa?gny�I�п�8ݐ6�)�A���i�c���-V�e�V��,����2R��(C����8�$������k�ǲ�!>�1~#��M=��%�?>{�%B��M�#͂�V+�M ��?0�62�a똛1~�����2UV*ty^��-�	#1%�FUA�&��@ 2Zl#4�����d�u6S��ZX`���b�q`&��b�
mn&�����E��n�2� ��n~�#�[S�V����;qbֱ