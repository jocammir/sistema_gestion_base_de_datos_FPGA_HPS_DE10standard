��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0���rΉӲe[��'�齹̜��q�o�*@[Tb��۱,q�W�aϋ_E�'��T���H_���(S��ӝ�@^`���#�p�Գ�t���!)��#��'����	A1�Cr*\*n�#dV@ �����/��f��>gaG�4�+��ʳ+��J P���u��8"���!��JG c�́������N�Xz3�Q������He�(�e�z揆nQ�`G5�o��J�a��`[��SV[I��:4��\�P�fϮ������l����6�����漧��W��I*6�)sl<
��L}ͻ������ݟ�Ae_��")�>@�	�lRPi�S�L]�%��m�A2��U����TS�y���W�bx��;�6U�b|?��h!���_���,���b�A
� H�V�Ti!;B�ʘ�9�j�!�y��A�u���%S�e$zs:��T�n�Hm�C��m���:���b��o߾Ņ��K�?u��~�<�6�S�KT�~@1k�~��U$��;�݆�`��z���g{�)RI��6Nɴ��q57ΐ7�%���Ӛ�9~�ۛ�;oc��8��G��e�7� �#ƻv�P��u�Չ�Y)��zM9^���Ɨ}��'��Ta�i[�\[�N�JA����"a�c@���7��@\���ZS��%>��<��Ij��� �\gʱ-1��f�(^�Z�ԕ���
�E:�&;��1�7��H8m]��u�����̦D-m9�ͳZ�Q��|��ި6�!M_8�L��B��}����M^�fm�A��S����~I"!"�5�%��g~���y��eZ�?��*i�R����r�bh�xj^1@��.�i$Ο�0�[Q	�~�a�K�[�U��]��[e��]��D���Kv�W>ah?��8bH��������#���^3a�Zo<���96奊gձ?�+�ӢA�0<�s�H�p�1vVM���+����2�72�P��c=��h�0W[LC��a�h���(��S�D}	ׄFR�#���4jW5�	.X��S	�s2��p�9�߇�^� �������`�F�?��e�ym??�{�O�`m����Y��L �����7>�C�O>�Hq�M�݉#�|�=(�fW�L��AAzڔ��]�0Ol�+(��^,#��wG����ҋ,��=A'�a�`q��.���w�]�#��1�{�M�Z[r�3�4J	U��Z͟��2֫1F�W�?��s��4�٠o�_q�^5㕶OFj������',F��?���j�E�\���	Y���
B�O�q�1��~B��Ҷ��}L�e�y�u�D8r&2��NŨz��z�#�;���ꤻ7���%e_�0e����
Ĺ:���P�Θ�uə'���E�Ub�	�̮�s��Dt��{��� ���jp$9"z	���������U��������M�냷s��ҟ�T���1p�<���S��Fݺ21�$0����`Y����`ɷ]Ȉ3 ��H( j�i㒕]pP��GQ�κ�aP�!}�=���j7z*j�N=���|�!�&A%�-��7y�N/��rO|�{��Mz���+~A���]�`�iz�K�O,�ψ�`:(��u�g�sz!.������+,B����d]�)�؁�hܕ��ޢV����,�>5�����\��g [n�f�[�y�O� ">+�f�u�g����J��Pd���+9�tO5Q88�ll(���%�����}���}�TFG�����gaz��h�g@4�6�T[��O���#O�=�d��$a/9^��W���#��7�����ɓ�O�/(nс��]9>.�+�6���t�M��q�a�v��C,�SJ@5�L�u�lӍ����6	�5R�?�k�P����~����.��&C�!*�ㅔiOښ)M O�cQ�D��o�4k�Q ��  �+N/{�WC�^�~"fwrI�)�v0�QV���>A7�f���|T�y���U� ���8Z������R��M��a�%̡��+�0p�Ph�*; ~��@�>��o\�`���{ބ�Oq�z��$>+���ǹ�]D����>����I����W�Ů`�:�1U@��h��oa%ᵸ�<,ovV
颡�i��(�ÚQ�~�f�\ӝ֚��ڪ�h�pi�g�D.�6H�����P̋n�-w�\B�� ՚�Y�E�8<"⭛F��6au��-&.�q�:�J��'�M�Mב@Po��CW��1r������I����5=n����WË�v>9F�d�5�J,H�Ԉ!I1�48��de�eF4
&��b��ݭ���D%.W:����A�d��*�r6ȿ����V�*
�7�E�	��P~m7k����`�f�?�Qڜ�i��w���W*�rh��زVR���̊�g%5��e94k��u�ǟo	����)fVsﭬ��ШVC�z�P�ӻ��L=k�g���̖������1��n7���J%�B�͗|[�FCrO�����>����?�w��֝Øa�7�0D_���Q:���	2�BU���� � \Wt�,08e�Zcf\:�{ƒ}�*��-�U�G�L��~W�|��o�VL�֝��ƪO�w�	��7 �B���.:3p�	pc���D�q��@3`�����q^g���ĥ��+D��`�[9�[�)ӉY��t�Ӯ���p�e]g�T�r��´=� L3��]��Fx^�����T�(7�4��xy2^�$K��F�<s��#��)9%�Y�}�[��S��M���\~y�譁Z�0����/��ڈ�IA�8�S�I{8/S�� �m>0 u�>�RS~����f�L>�w�x$�:ĩ�x�O}ݩ֋��������j� 77�a���c��[+�nc��k ��Zܖ�R�Є!NNr%}ǅ�{�AN#`��v4�D���e���[^��h�2�=���>��Z�A 3�t.���,#-j�@`��f�I�v���wgn���,�n]�OE�}*��Ͷs�.�xA\�_N���/;aF���]�Ws�PZޯ���%�g�g������sv�	���M�t��Z�a��űT��Bs���V�a��2�`!֖W|�<�'y���8e����n�yn�����������&@F��%��\�P��I&����!c��ǩ�E�-T)ё����T��9��j9�3��Z-���NP&���+��A�%,�����վc���1���OsX64ch%�R�9
���4�:��O�m�b��A��tW+0�u��)L�c��ڕ��W��~tڋ��#��$�n��U`/ߦ��U�zz'�<uZ��6tP=ľYg:��d%h��/0�ዋ�K�q+N��,�x�wg0�&8�aD���a�Sb5\e0�#z���� \���-"vƝ;��g}� GWW��\p�J�Ґ/�'��u�/[��j��X[x��lJk	��OE�i�����9?	FK�d��� ͏$�O=N'����y,�jBlO/|�U�uY�?�ś�5��6�-����&����QQz��K�<��Z ��#L�����6�/ܐ�j�<cB�6�R�e(��&BS�c�8��i�,��*8�B��^H*�a4�5�`Gs�T+J���~�@H��4�fJ"	���lѹ$��X(��K��x�����k1�|y�~�uJF�4�+�-�y~�滀�<OQK�Q�	UC%x�yX=�E=�D��m�~���5�K~�RA���u%H<J3a��[/�B��*�����	#�;sXDt�%�Ϟr#c��8z.p4k���M����
��I�B�	<�ʓ4oW�����\fKs�3}Q�m]|�[0�H�o( +�"�Hln"Ҟ��2�{e72�U��1~$$&`\ק��V����	)���K�h}�2��ʲ�� ��&�Z����6�b���'��#�TTP�H���Ӝ/�R\H<�6�Zj!B�&��VBo`nhŵ[�����k�.`��T(��-���$q�I�̃f��I?��9�� ߻�Ո�����Be?�|w�J���z�|4�Z�L���O�2���8�b��١[*���{D-���c"9t�N)�,���x���Z:�������{�T�}���ٜ~v|�D��Py�$A����x\(*G�
\�?�`ɕ�yS�g(�i:�� o�D̃�%í�-��X���"y͢��J�E)&ܩꮆp���o�����5Sy���8D���i�`��t݆�� �hB�$����%���0[�9��K�.O��%t�J�Hdr�oӕ騎�8��!�,�9iN��a�\���Џs?t�o	"���Y�k��xĀ��̞�&����;��P�FýG}�9��������I܌������=����b�-0�vY�Lj?9PoXCXrUN�.�b��@c��2�	�w��b]��C;��X/ad�Zo��v�,ܢ���vQrrK����$�W�������?��18>}Wo0�'�}55��v��R����2]ߜ7p�ī�q��*�qF"}����I�.��,��Q eEY #���"��K���;��k���v�Ƃ�����sjq5\��Zi��\ۮ$��P��I��&<ǌ�Ig�Y)���L>����"�j��N�O�G���YU����*��!b�@+U78\� �Ih)ȧ�nf��A<K������>O�x�j1%��|^�u�:yY8��/n��ut�b{�3D&[�2R����-Ƥ�-)~�g��a{��qn��^�h�_~e�;G�G�!�i��t��R�=�OX-�￶v�xg
��4�>��g���{���,:�-�^?L.�
�(�ѩ��.�1���'/k���7��ykK������fo�t��n�s]v.�����r�����dZ���Qu��>�h����H+V�0�7��o��RZE<�z>�bUK��A!G���ek$'�y�U0���θHM����	 I㩩G!(L�=X�T�@ q5ޒ�E�s�lV���N���^���6x=[�GR'�d�x�L.�9�4Kfn�/���/���6�/���#T���(�W���G�Yy|X8{����5���ǝ�����Z@yvܵ�`S�8KBG��=�j���XkL��Z���"Ǉ��wIU�Lઍ���_eQ������ⵈ�PDM8]���ҽ�7��yВ��&6T�����t��!���TxQ���b�&GAf2=m4�H���?T+��]���ګ��#Z�/+����e�� ��b�I�[��Q*83�,���	z�~�/��5JY�"��� �iUQr��u�z|��т(N�u�m�2��� ���4�\�P��r_�\��}������aɫ�Ajr�����V�l>Qa�ߞ(��m�Y��Nek����ϢE1)��_�3F������q�=���q���l&�kG��y����#�?�N><_����3euʜ1Ɨ� D"��� ���P�ؖZ�Q7�ʃQ$�a 0ݲse��u�|�!�za���.���muk�_�RG�:.�I�V�#��˸�)�ۼ�J�w��:��6�v�℞���>�G���s�� �Y��j�m���Rp�z<v�w�#��):��x��⨣xN�LT�q��
�4`�ڼ����X�h��Rۡ�	��n-LH�7�.�-}l{�V|�u笉�,w������BjI�_ԶI87+Z����G;���@�?ٞ��7��$ߗ��M��{�Y��J��2u�a�c�1�Vø�Qbi�u5�@2��lo�.�T%��{��|�Xi@ 3�u1�QU���Zs��E��&Ds0�~�K��J��jP�/b� ����W%�X��2�~f��)��o��D�iu#��\4�����=��1�vKO�+o�~�*���W
�+�V�o�ܤ�&q�y	U����(s��Y���?k>���]N�4x�BItm&u�t�;�E�k��@�[��F����V�pw��	{�"axu��%;����o����L�/U
�4���L��D��[��Y���g�VЪ�.�A%c�Lq]K�?��c��+��G�.�̻"����������1����J�H�����Tx�=�s�$<&��x�<`c�u�u��<pk~2��g:�bs�4:q��U��>X�M�c�I`-�;��zM5`[kZ�KOa��e�@ǿr���0�e�>�ܽ���a�^�|f9x%"��</�#�?KӠ��wnH�#d�]��S�گ�P\@���e'��w���b�`Td7�b�{J�%��`��7������?�B/�Ea���4��2e�L=MG����5��N&¤�Ӽz;�;� NA=Ԫ@;�]֗�!Kr�^B4�q,�yӓ��k.<~4�o���P@$��Fݏ��G'qڦZ��턩�� �1�َ�n�	"�ԉ����*J
4�ab{�IUNP�M�����5(�qܗ�c��� �Lځ��@ɸ�����=rd��.E�J�&�'#����e�2���,v6qͺ7�Iyӥ�7��EC���`ڤY�`�,!Hie�G�g��9 ���5J�gI'=Q��=n,$V�ab}&2�YV�, aT�}�h}�J���A������1+�ԯ���g���3s綃��?A՗&��>y���0f�1* ���2�A�G?T?d-�K�7�$FM?��b��ޫ<Nd_1�6.#�zz���EXJy���Q�Y�N�4δ�D��n�'���C�Q�S��v%�
� L���1��/��pj��:�c�ċ��ZfV)��.�ҹؔ��Ũ���D[�.�񠒞�9�I��l-����XS�U"�EYC&՘pz���5�"�����N�{��0ܫl~H�l��~TG�t���|�:[�P3���;O���nr�F�8}�!\�/,��H�X��e�1��Iu���Y%�Lk���r��q��A.��)�I��p{���#���ͧ�q�Hb䤠X(���FՈD
*7����=i�G�
�Qo�ݱ(�>�X>���VD�aEU���1�lD�����ɖ��T<=v@!JJ����-��;B��K�m����d4�`��Vlw�: ۑ���(�3"�pv�`���	�R�I���=Ꮮ��4���Sji{�WLѹ~3�`^�3����g��F#/��TN���'������o�H�l���ٮ,��+���R��Ǜ�T_�����c����d�ٿ���61ү��SWYx�U�Cu������j3Q�eCʧ);֕;b<�R�L�E`j�6�z9�'y���k�^��Ǌ�x��'a��iT��-�J�⛜��y���(ᜲό;WK�Y%bӠ�Iޙ	�{�:��O�/� @����� �)��mF���Q�dIG��������
mhr6K"����
u.u��Ӛ^_�y'����<� ���^�8�C�������FQݨ�J��
�Z��3G���x�EN ˺�迏��O~XQ2�vu��;� �6X_�8���x��rE��V�����ಎ�uO�n݋Dr"���x(�����)ot\�"�̵�t�9����~�	�9�+�;v�|���&��Х�~����B��@�ƶ�R���V������43��b��ވtt��; g�Fl-�,����������}e����*fauA��?Ǫx����X�7��DL��M��K�R{qԔI����Ǜ�jn�E��"%�%���ꪬ�*@<��a:'!� �u.j=;`�(�⬜`���*�Ql�%�ʏ�Ohǿc�ht@R�3�/uW����x��������)�Yz�kg�3h��o$@��{N[���h۫����`הQy�a�qq�YĮ�D���d�oKPzap��+bh3��#�Ƨ=TI�T���"��S�< !RK��v�<���g�R@1K��m�3���D�we�ѓܵ;�K�s�<��;���9U8fnO?5B�� sj��1����q�ڎ���G3O��W<�.�IE�L��)�)�أ��"���G�|�5�䊢>Ȑ< ,c��{�_��V�}�3_(yJ���H0*�-=�c#��}Q����F��������T�8�E�Q�]q��ͭ� �R�Smϒ;8
n�R� ��w�m���Ւ;N�,�Wr�Ai0���J̨���/���.Hk��փ>n{�iQ�����p��)�LS6�4�g�&/چ�YΌ�D��J��������\����f�B���Ƥɶ�_��D��1UKMf�P���Od�U��L��&�dae>_YwM~�q��
�h���eU����(�s7�*�_VA�ȱ�8Օ�"����M��<d�e�S�P�g�6B�J~�3�Z��ʟN���AFq�G&�]�<�D��]O�_��dZ�y�r�NQݔ�V���M�gB����cY_P��K_�\�,��t�7�(�ǈe>
!�3��*��EȸW�D��t͐���8븃0��8n������0y�`-}�69��>p��)� f�p�ss�F���]Xwu6V1ƳG��95H��j�0`�_�S�%:p�	)�qLU�_
T�C<G�ۍM{�����I ���Ȟ�	��X����6|G&��r�&���䀘R�,흶��8z�=9�Η6�7� T��Q�m�#Zb9��D�5Aty�u�d8�s�� R2�1ħ���b��P��I�K�d��^�����Ƙv���W2��]9D�]��4�hS�pϐ�;d��A#�tG�x�B%�U�֒0/oN�-%����q���4�|��3[:���+ %�z@��tƼ�\D�Q���C0(��߅y� !5�2���t���_�Jq��_��X�C����?q
(����{+x��Ni�hf�\��N����� �7���}*5*zF
^��B ���9w�W"�N�BvG�t� պ�3�� �K�}�/��hҪhK��"
5n���żSs8��/2��������
��|sr{��)��(��u�:o�_)'v�Y�S3����[Y�+{JrǆF�UL���T,G�)E���p��o<;��pc=�I�cW��c)���?�'���),�,�@�Ӌ�3t?�J��K3$�'f�V�G�aN�L�����-�$�|�d�P��B%�ͥ@��U��YQ�e{�mz*	�Tr3$�Fﳍ��Fǹ�5��R��٧r�����;�y�ҏ��>woTW���)���*�{KE������:Ol��܍e��1�b�sfL5�n���z�֥��=���ב�-8)����̑]��s��@Wo}���/n0,N���]��E���E���Ɵ}O��nk-�4�ݥ���b&��p�(pz����+���˰�n"G���:�3 �]`���EyV��N��8ךC�&#���^$�>�8U�j�E��:�9��Kƣ�{�3����Y��)�|����>E��2�#%;�D?�-P�)63v6��#/;WH����H������d��Ey���ܮ�]��$��U����#[���4A���X��K��ּ~S
�:����ƣ�� ���a���0��2ǅ�)
y��I�>T�z���j.�,e������A$�v��5�&i�U�(e�ۚ����wo4ߓw}h�"��u����1�lf�1��z��bQ��?"�J���'lʏ���@a�+S��� "�)ȱi��3���)�FP�o���+�! T�C��}�$��	d�3&���9J��?�V�;�]>^����I�}D�0��`��Z�ޕ��ɵ��BXUh��I
�$�$�R����
�剶?液z���=Mx+��=��؋���ʕ;)��P7�b�L
�����/4�?@�{X;\(�Bؾ��9��u�H��&CNܚ'�.:}I��� :HadYCOw-���dl���fQ&<�7fPM���O5�M���<��|uNK��K�.��S��PDG.!c0�`�
���VA�q�*��vefXL�$\+/+���H�GL�甙����V���p�����bݵ+��j�Er�_/��N��Km$r)^��ْ'�� ��^D�Ry���4����0��8
�nk�2#�]su�#1�,���e0#�%y`���[�����2�V����oB����}nQ��xFBbH��\08��]��Ry�H/����4aie:���~n�H��<���*�,����.潄`�l���9�{�&����Q��� s�1��Y|�t�� ń��pŹ$���i�1���r�Q�7>+PM���[$�0����rY���e���Q�#�ӛ�Z��:Z���$b�YI��*���K��#C���S8?���^��uX�ή���:H�,B+�o�/�r��|����Ͽ/|
~��A�c$�_��ۍ�h��i��7
#s����p*���M\�(>�ofg2���'�R��d�}c���"A.��o�k��s�I`��}vf`���!��}&��f?�!e��\|�r��|ZR(�hPۀlvyU�^2S��T���;�y�r��0���C����`�wj*'T�B���G��t��V&<���2$Je�H�d���%GY��|y*]�k,�M,����;a5h��A�Q�]��"~�̚�Q�`����X�9L#��v+^'n�Ibs!5H8���F����Jr�n�*.v~�|D������F����L��3�*��Z��t�j�����ǘ�$JB�x@w��j��)��x��|�	����G�c��q)�i��-�+xV�Qe�N$�GYgH���q�w3 	�
�#�Jq?A�j#�}�iH��d���`.����\f���I����grY�������`R�IjrE��EF���U|x\����v*��ʖ�8���y��#Ţĭ
�������K����m��Q��{^-��뚬�m'C�p8Dr,T�jy��^�(����\(gŋ>��F�m�eHA�<v�v\�RD'��5r�����밉���䐵��[�� q�ޙ�zx���ޓy]�O�'B[1
��s@d�@�Z��'yCxq]*��������Vֆ��'�g�A�
��D�{5>��*0X�����nu}�6˒M��r���5�2ϭ̩)�� � w1m�����T�*�ߛV�#�rx�Y����*�#��EW��c&�����C����<�s�.XΌ "~��V��_���P�X���b`G�x*��"Ñ�K N�c�.!8�u㱎m��
�^ɟ��>��@�1�M�M�W{q�� _о��-�T8���X�������Sag~�m�n79�E(�����%��� ���h�Xt640ިN坣�l�����W���d�p�(Zd ����w��p��5�jD_W9�a?�l*?�?+�3�ަ,�8�P����$Jԭr���濋`�5[ꊐ�h�B���^q��>!�G4=F���c�� �Y��kѰ%d7��Y�;�Pה���0�	��~��E0�p��5&�9�ʍX>I�����|��F)��A�O�A�фw�@�V�3�w���-�k@F�'r8��J��;}ˉ#ڌ!��i�*��:�B�G����N2_�&��sv�[#�����j{�G6����W��h�LJH0�.<�Pɶ{},���!p2���R\�-����YN<�-O��V}Ad�t�G_Z=lޮЦʡ`x
���ã��T)[b�ًK0ܽ���a���~+N@��<��\�H~z��tQ�"fd�M�-��j1},���!�qY��j�m@ Tۂ��->��ԍh�i���E3~vz��o���y�RrWv�*�+�/���8�U�����7�d"%�_��W�*D�Y��"�eT�,l�2�:��i�C\����>r�v�{3���� 
���5��!J�2���0(�wAX]&�k��YP�.�o>U�W�����h��H����e����,�l*Ȇ�s݆�e(�Ӭ�_��}�*�������&;�}��g�6Q� �u@��T�1W�� +�,�\)8d��3fRD������F~�;v���J9���f���a��n#Fn�����d�F��c�D�|=&m�S��	o�AT�ɢ�sWԕ�������f��o�_�����i�͏K�@��mI?gq�t�[S(S�m��Р�DB�RHf��d>�{Gi9i��%;'	�5�}(�<�ҵKڱ(e� t�<��K�|I��Np�B]�P�c�4�=n/-F+7���U�O���ho<��� �v������v�G���Ll�����f���n�x7���B���Z��{!Bd�3q�I�0!�54�$ZF���� :���$�+��ru�N�X��+��z֛�61�g�C�87+j#5o�Ȧ&�0�@��en?��'wGeU���ȍt*���,�h���y�����/�Z׏b��8+���ܿ�*]���A�;Z�z��gM��r�'+���nf�-h��l-��K��VU�ԑ&Y��?�m�4U��~ߙ��9�>�ÀuY��p��D�z��x�~�|����*|������{e��~%"�Ɵ0��=�z1Ж��њ��A�ZF��,�6�)޻�ڽe�F~��^L�!tcڬ<�i��h��M�j� A�)�a�ى3���P�����G�g�k+	�|).���g NǛt���P�bW,�kN��v��a��t��f^'�g�u�XI�7t���5��Q�Uk+(:n�)g4��j��H֍U�E�פ��P����ڹ2>׆�FT�/Iպ>pp���y�|����Law7�z���n� ��$�� Y1z��u�Va�oF�TH���w@Z��b�+��vl�_�&i�.�p~	͈K��OU�G���o���׬�ɸ�r;��kgr�҄��H�����;Jb</�����w[��W�)&O���C$�!��8XPn�3�5Q/�� �r浗= ÀF5���Y4��I���Jf���*K��	�ly;5��;�ٯ���8 �9��N[o�y���;�Q�(Q �|J�z�I�CZ�ӆ���;�Ü�ͮOc͉��j����l��D6��)�M(g�l�2�k��h|�PwYK�kK씓�����f����1P������	�K�~9ʖ@`����hϙ}~y��ܖ�U���<*�6z�k��� D��%vA���꒙�s�-��;�]}o�:�w��������v<'I�Q��F��e'��&�+����W�{���UY+ �W���B*��Y�L��4D��r���S�Y�呖��Id��T��4'�]HwM���^P�^�;��}ê�q�e�;�{\-C�CO\w��y�B`�
c�b���.�)�a����'~*o#��6!���xl���D�S_j��H�k�-���_PdL�r�p�[�2�T��a:�%���e-!��^��ߘp�f���!�֛ݜ���$�
Q#l�ڐ�)���Y�-O�L��fg�y�i16�t뾷���v�5���݀_���'7�Wp��ff��S�I�f"b=s�q	ծ�ѽ�;)1�ke� ت�ׁ���,
ƞl�*z��c��-G�jV����d\�˕-۵{��Da(�����;m����(LJX�|���A)���Q���/F<���o��'�K��G�Jw�l�T��*�8Gk�׳>�;]Y�G�����c�U�\��B�$����I��:F�,�q���q���ѣ<D�,��ی�Ŷw�a9G\��y`j��'�b�7(�2L���>��fƛm�{��L�1 ]��l��:��b��.�����j�\T��k�$��H&��
�9��g�ib��JK�M=�Ϗ�݋ƅ�hy�<�M���嶂0}�}����Z1K4}m�b�GI���1�G&NB����?cG�Q��Gټk���]���ןl�R�'�0�k��[���@b��.��&��	4�{E= ��е�b(X8C4Qt!��`�Z�������ua:[*��S5̼�x�]���Q��(�[�Z�ş[l�s�&M5H�uq��U�.�L�$8���g���܅+X}&�g�ߢ����X'TVω"b��ε���@�Y���^}9O���0N�O;���C)5���1��h9�&���3��gҒ[މW1?x�^j=E���vwoR� s�#��� �b�H��/��]%p�oT���qϮ�'�LRp��۠�Ӿ������ S	�?S�ܴ�(I@z!�rE��[B�P+Xʺ㫒Ʉѧ���-��	�<g`�^�=0yV���M�`Z�EtԸ�������%����6���iUC=�I^��mR�]���8�K��/TP?�c�����d���.����Z(W@��@  � ���{��)����u3D�a��%;�aI���T�FH	Pf�3
/e��t���<�
#Q�ڙ�G��p�F}�
s�J��3R�Q��h�N�12z4��m��:��3}��"ͷ�G/N��L�=P\�hB�x ��2� R	J�r�r�0�VƋBU���hf�BĪK$Gzn݊���ߊ��lL@�]yԵV���/g����<z	h�b0�B�0�ûe�B�#���e�;�!"�z�+Q�)n�>q}�6��e���l��h��-�=[��~�mk�1�zه㳓��|v(�7y-x��j3�3��Ft
�g1��!������눹,lMo2(ȳ�M���q�@�
��Wꍤ�'|]��D*�<��~�I�4���m^�;4g��w,�x<ClU�㘾T�0���C`[��C�ї$` ��ȗV�ðJ2S��k�i�@�tp��/%�ث4/��Wz)��0���H��/(��Ʌ����|����x���P�d$����.⣒��`��}��(�n��u7���焽��4�P�-���M0L�aN�f;C������{N���<��k�+�(;&�wiG���:k�>���3n��ϭ�p��4}�c��d_�%��)�PbO��.	�1'3��qH;�M�����qxe���d9��բ���3��!,��(Le��~��V�������^w�jM=�xy��`b�C�t���