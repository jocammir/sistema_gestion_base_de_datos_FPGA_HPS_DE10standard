��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�s^W���0AP�<7b�HFC,�6��^���v��T�F�@3�e�_�Ѿ�bl�^��g0�1�e���`"_�ҳ���� �*0po-�6��%zڑL�9���B{"p���:�g8��ׁe#�ӽ�K����>0/c�	J��:����&SSN��/t%����y�@��%�v[,�C#��<��ăӖo��U�]�k �σ.o	�Y�p/<��!�gd��tqd�B�)�Ǹ4b�y��;Q��WkC����������wC�p=���?��2��P�֠����M&SO G��K��J�D �X���YZ�S�u~��J���ɣ�|�b�)��RI;]�$~���)۶VH.#��Ѭ�~�,^կ諏0�}�d�+����G	E#}����.Z�2T_���g�e�9�
p��.�O������S�g���g�ad����U򆯚	�ـ����$��tw!�_y`��r�9%����Û�w5\���	Դ�P��r�A���~/f{٭ڷ�
%�.���k�|W��P�9�xc'<�����I���h�cIw��Fƛ���闉�����zd������5��8�y�1�\���0�_M 9)N���DJ��PQ����$�k�.��	pPn�\�G&�ٷO��}M�╌�x/�p�*��g�4��NA;(����2)?���[%}�+�3�sv�|��J[�) k1�ȝ�_�u��$�b�ְ|��fð�ۤ�%lxm!�:ԯq�����A�w�g��!���dh@���%mo�:E�&f/=�rt�TMȭ�������"(ßSE�����#�*�ug7�3V��h@yGmLa��Q��(A�o���.�u�:=��7u��j�b��K���M	��DH W��(� _a'�B;�m��V�(ɹSQf�L������9�7����ʈ��+������w��OTS��¬p��Ĵ[n�U[���C�n���΍7��Z�� ��-\#�PF�Ws:k��	zq�!��6�hM�8H���������J]ךsԽ-"�=-y&O�����P�����v�-�� ��r���I� j����-}v���� ���HvQ�$�_�sX۬�a�Υ#Y��i,�\*XL���Ǽ5	���r��W����1b�)p닦WrC1i��j�ϛh�%�^���s�U������Xc��ܞ����q��+�:H=I�X��R7�����L<
T8�Z����dԘX�0���7�;����u4ͻv�9�%%�1+C��(j�k*��]���m���������1���S�f�N��%�:��SW��r�]uzi{J�E��ڗ�D�ȕ�ԬR�o��/�lX|��P��iHh��Hd7Z��O�`�ҲW��h[O��=���S��׻�?�%��a��f��q� R]�,Y��-�-J!�Q�ձ}���T�^�s�H�f���"��p�s�4!��P�J����(0 ��"�J+�8b�&O�\��o�1凍З[74�5��Y�����,�1P�%��qG^S���U�DLU�e�X����z��� g#�%����r�D�&ǈK��(L'Y���v$i�ӓށ`�V��8��u0Aw?�ccpmC�*}l��j@��x��\s���cXqm�D��9�/TЋ+_�B"S���!����e.]wM��u� hr������2x�y�ѡI^�i��/��}� ������	��̶���F�U�%�
AE��#�P �B�J!AW�;"+����<�[5,�Cv���V���F����J�c��*��r�lQ��q�j[ȓk�QU��y�{�Q<� $��u��L �P�)���H�?�YK�����'j�Y{O��A��r�8a�y�I���l/�y��;�Tt���B\��DS��5�� ����e�����]��<~])���̙�����z����,��=��l-I	G����֚�j�)ײ ������XYh��d��������9����~9E��I�5�Zv'���� ��ҫ�h�E�lȣ���$;=���c}��2/�tK_��XPg؍�f��� �(�ֹ�*��1���*���� O�Z�
��;�:�˶��^��M�3�s�3��Cp��H�ReT<,�=��]٫�Z�y����:.�9�#}DE^���-����s�T��n�6#Ēܭމ_�t�̽eK�e�߿�V��O\]fHֶ���̄H?"�4J.��LF5v��o <�pD��@L�ʲ����[~�:�\ǦMp��8'��A�AV�<���bT��`<%��B���t���7F��+�����5#�D�b�N�7��>sa˼=����Z���:Q F�s�
�y��#��aU�����&�yq�B���C���ڢ�F��C.��SxXH���cC��%^h�;~s���z����<��|�,L��?�a2�%"9�6���&?����`���iyǮ]n<�B!���1���B�Y'�_6'�^fV�XD0���a�>zW�@w���>����4'p���Y?���1f����[�o�&r��Co@�J�X���s}iȫ-���@��(��~l�!��(��7�����>{c���~�66��,��d��Xz9�-e{�B}|�[L�gG�����v��|z%�MA2ދGIU�.s�͍G�k��,�\�"��@nw�7�1���-<��/'`O�RԔ��kh�����#�U2������fx��N�$�c��ŋ\���hLԁ��S�V�,�l$F6)��%������M&q���'lI�pl&�$~�)�[jQ[�Y�ӱclJTB6��Ղ�䇪俣�Y8�I�h3�Xe>��Fbܛ��[#n���8�d�R_aЩ'h(p�
/=kA�mI5o�<��ǫ�{��"�!��>0۬S�*[�l�7jі��_� �� A	��轢�v�3)Ҭ�`�������]���9B�Õ�B1x= ��e�X��g�W�
_�k�N;뢱W��iʆ�T;- ���5�����ԙv�����Z����5I&J�e��WW�"nt��X���]f�ʹ5�h��R���Pw�ޢm�_�S����Q]�6Kb3��I����}�Gt�?}��>`I���@b����}|��ٹ��h��)yJԏRX��b0z.�~]A�6��qAU"�:��.���2B*#Zy��]A�Z{�� ���g�X~��z���m�b.O̾3��$�9� ��l�T�y}�������q�ķ;>IU���������������ӗ��5~W$P}����<w�Ou��eV�[����u�z͇�X���
4�M���ٮ1�9~�gm4��[������{$�%��,��d{]v��aT�bO�"��dm
��Ct�U­��h�-f��E�_,gѰW t`IBN��b�`�ˢл-{�rR��".�^0:���iu�e���p}�%���B��vӿ�z������	5��$#�l
����k�Z��o2��"�@u�R�Ӝy��}�y䯐��W��ʠ�P
N&�B�[�ń�̡��5W���r�`���[�|P��B�\���~��|#��o��d�"u�o~7�3P�0��AX�V�.�,�	F���Y�'?׀����%�e�"� ��*�4�a'xn'��}�[�7���?����lOrRnn����X%��p@)�]�^��&`쫱�$�Y�ٲ";�r>L��/��'�_����+28"(j;�rmNN2��.f��7N�M�C>��1 ���H����sj+FfS�%+���&xƑܡ<<�u;̴+Sc3]s��"����X9��B�F��p~0�X�p��O��ᐑ���u�4���2���Fq�L
Э@H�3N�|�ݼ8=:����Ϛ��J��@�шsAw�a�����&��4�
<� �XA��m>��!�ȑ/C�"�i����P9���-�?��Є�,�"��tSG�2�Z�B�N�8��/η����NYz-,���!�x\��������eiZH�P06q�R�"V���~\^f���}*j
��+�����,�yز�i�s�4x��>����F��=��\�Q�['ᖣ�I���Nm�PB�C8'�M�7tD��Ũ���@?�q�sћ�H���"m	���/!%�$<ù\F/`�P&V���2�X/|Z�œ�~s�����9�U ���j��q!&B쏕F���R._�����LO�;MX��B��{_2����̠^��b�s�t	թ�H��[�J ���(Q�`6�+Q0/G�AF���^.0TǸA���$w&2𙸕'\����BcC�z��I��at+d���6 DX��,yOHj��⡉�q�i���@&բ�΁R�Ah�]���xp�� a(J�)����:��?�W�W��%:q�l%Z��>����\�%	��@9H�_� �|֊�����_3�
s#H���2�ڼ��k7�F�+)��='�Fc�V>��d�D���"!]I���t���}������G=�q��+"�{T:_Mm>�6F�0�N;�nP���Q��1zP�j]F�.�B	M7>���gZ��!���Tp������.3�P�m/a����f��UyqY����f1���{d���e�ԿѺe�`O� �ݳ%������G�j�6��*�%�
[22J�Ko�BQ�ܭ(�D��-�csq�E�?^����ޢ>�X>Fe!�����י�+�K`���7���]^e�[~�O��Y����B���:@�nS5�4>#؝�Xǅ�v���q��$G��n����>~<T����#T깨H�?h 6�~��V��.��Fi�AS�9T���g��x<`�g���w�.O�XC��F`0�ؒ,t��Y�f��=ω"��N	�A�s�0I�9q���䮬1¥��o�;M�!���w�L����$\�r;��Z���?�ѿU�*v�.���S*�RU's	�UH��%�V�Q<Đ�ʮ
n����7yj��O�AW=?'��	�㵓�b��5�{ڛh?�^�Z�����b�#�������o�w�5�^�2��xz(���o;�(C�B(���C�k�m�Ζo���`����P����8�s@��gJ���K]���=g�j�7Ⅵ�Xg[�t��ɍ_&��ClpcQ�Q�"$�)R2��n����,lˍN�V��h���|��]��w���\n�XTQ|�3d�9̲1�d��\�?{�+�1�P�D�-5�xE�6`�2�I$u��"�L1�}�ĭ�yRB�@B��pmE�#<4����}��ȳ���B��������'+aOV({���7�UO�&g�1�o��dфȼ���~ J���S?o�>���E��>}��$n����O�N�c�`�{0���v�,Eg��(�19�-VB��3QB�.�}�`��zf"j�2�`#+?������?��u�V�aW��?�M���� R�m���Ӗ�R�'�.��*S����=J>V�����FY22;#�� Ğ8�^8jJ�;w�T�P�޵(��H#��U}?�������7U�E�įx_s9��c(x�k.�|��Ud����m���.��*�9yZ��5Nb���g@	H:x�My�	f<lOQ����nj}M�78�/�tk���~��Nhȳг��:��el���H%�=Yi��!���wF⯒�Ɵ�\��J�m[��0*��"E��E%��C������p�B[���< �4������h��^,����ڣ�Gn�$������Jq�)6V���E�W
��r��}z���u��6���%v2}�$F܆�;�XL���"R�>d�^\���$?�KL5Hv�~i�sQ#�z�=s�L��@g˟ŗn}5T�<���)��0��%��PH3�ِ8����P
�Eܵ��A�9�8���q����{2�u��)�6ݛ��LC�%�8V-ߵ���R����q��1�0��&�z0�	�j�DT������Rf���Q5��7m.�4+�?��{ڛY\���fy[*V���b9����d,�J�5�[���~�ĥ_���%z �9�M�(%�c�&�aѪ�'7I��d�־�S*q�ଫID��r:W������{�K�}��������S���{)s�����u',��X��v��ٟ�9$KR�'7�U�~~'��� jE���.��FHq�KT�PJKR6�/b����0t{h~ ����pJ��M���ԗ��� =K�|w��7��h��E���-Vyv����Hݐ�愚x:�g�����
��X%(*o	+�.z�������C�7��Z�e/���Ҳ�"��x}-��R0/�
uN˂�� ��*��"�+v)��a��s|�ũPܤn�Z�-n�Z&g3`�j�J����f<�ς5q�pJ��?��W�+����
ct�LnE�by�۝27+庣Dl�?�I�J^�������_|	�=c��.-_��ڜ�b��jϋ���ns�9	��M��C~�̱�`_1D��`��F�U��Bf�=ʞH�� eM����QM�X���a�����m�<:��KD�[�B��f�0���%Ýu��J��ҽ3��	CL�*�ͮ�M�a9j��W/�i�b!N��I�x�%�`�V<J��zk�t��F����P��{����C<��g���8�I@��mzIa	����$��j?4�00׏����Ҍ��o��)�Wy?%V�	��J�HO���-ݮj�F�?M����2S��E��KS8�'�G`2��q��9��:�,
�Z��,��h��;}c����y��g�;L�z��m�����g��`�}���b(�8����hQ
�V�D_A��>ď2�n8 w��������vFp�2�.��������R�兊e&?�kcl ˸��d�lJ��,9'_m�Bg����y>�8:��;�nn���19p�L��
.Ԝ0���c/�^w�d�(��;=Y}�uH����Gz݌1wt�-�3a���!&-3���C�V��o��u�#�ע'%Hoȝ׮j�n�ZN��U�>��w��'���n�d����
]��ʄ�3:`�h�l��~��`c�MH��N9C��&H��q��$�`�ezz�_���K�LqY>=�Or�`�����G�N疰#�'p�_�.{9���v��+V%A,N�8�j��{�ƌ����mI5)r_�)l�ğ�c�tʡq�?ն��8 �ltU�`��C��棌��fțf���҄J�hH��s o=����)Bx�>]�=i���R��x,��V�Q5jM���u��8c�y;��,`=e���+t|�yD��H4��*��k�+��lQ�V�{\D��2'KD��[TUK(O9|�t��Ӄe�~[Q�w?�:oP��?S�jd�>����.ow��������W ��MbUx��Mê؇B7o��H��u�����G��Y�\TR-�`9����(�kQ^�{�"���j�l���$���)
-ǟ�3a�!/X]�-A�~rl�Z^�'5��f���!d�.��mJA� QȊ��`���G��o&A��H�kl����4TUx��G�>��w+�%@v�˭t���\֤ȕ�_�$��Au��<��NԨ)��k�@��#�V��oy�c��6��Z�'`;:hs�I*�5�-qG��T���\OWN��7�r���cV<Y\��u���OՍ��T1Wz5.�g����)ř����9hvi��󻛣�V߿d�4�{(�6�+�;ш�<������?�@�M{�%�e���Y���K'�:��Z`��NUg�J�\����Y��f��(��8i�SG�0�b$r�����r&�դ��̮����,�r#��K%��SmsAP�ӏ\�Z��Iz�*�H[C�?'7��,�Qf[;�$c�s1��T��x�g�_���Y����*��/���C��(�̌��}��W�[E�x��U��ԕ��G�2���/m�ZJ]�A;���3�t	�t��%Ƴ��;ʶ��r.�bTDJ<9�U8L�`mw�-H5~�c��(ή�;�r�:�|�QL�P��
�L�:@��Ȁ��{w��o�Ad�/�}C��:����q�xz��Jg�ܳ�<���D����^�}���:���,
7�+w�7x��a5��h�xQ�B��a��7��*)h�1#�7#2�<B�o䝜��3X��L�����O������dq������^�p JR.T����&qgl������-VL��o��l`�,�%Ѯ�ɓI6Kꚧ�&P��i��p�����w-����.��7iP�o3�&��{���}ۊ�`j��J�14��ۧ��<L������ԙ"��
+R0U!�M�qE�x����L�_�M?��d�U�WXp�9Yod�cy1<�s�'v��8CH��G��h9ɳ����:밦�*S-;�g���jb&Hy���)��U��x�r�vw�!ҕ\]��Z˾3~�xsIF�׬̧����$�w���y	6U�M_w���%&A������Ϳ�C+�޳3=��P5���[�9�b��eGl`g��nW���D�|bK(ӕxb&��M�g}���p�39���ο'�FCj�L+�텆�V-��9qll0Xm��/؎Ep����sY�A�@��g��ŗ�ӗ	�6暿`��DO��v_7h5 ];̇�;���s�AB�'~X(�j��z�$�L��z�'��lFZ;۪x�'��cp�k�.V9�J���j��4�A��<���x�,tǒ��;��t^/��?`�0+4j������J0ج��vW�Ƽ8cZW�+�ԝ��y���x�l���%`P��5�6�/*ɓZp4��>��d;��#b�<�~ -��w������;�+܈�I�S+$����~�����!ƢE�OB��OD�o5����b��4Z�X3,C4��xD(�b%V��_�MrS�Wg�a��yڙ/B dH������5���9��}Ex!�Z~���n$��VC�MOb	%�����L՚k�,�N�q��:�?Ӣ%|X�%K��q}/�79��*���ܭ+��C���@�"(�� g�W���6}�8�МNk��ˋ�3��T�h�Ԉ�h�6��J7fU=]��i�X�Y���6q��J:��уp�iV�Z���M!�����tE#��1�be��G4n��G�<�p�л�~�%t��>��ĕ���[�)R?M��b�=��!�V�PVئ �^�
�՚�_�x��iq'�1�i�������D_}}�����Dc	Xޛ����G�Z��{&�r��{�ܶ��Eo �Jd�.�8���N�O�n	�,³�|��lpË�KN���M&0���[�`�u�4������ͱG�� �y]��։rF~)��V��*�o�I
��2X~�3Mc���#�������hԑxk��������?`��
��"�*mҘb�3�@I�Z2ot�m>�+w{������.q��@� |Y����v���S8!q|cZʿ����,RF�df��/���K��
z�5r|��xmZ�g����-}W}3��1���bۯ7�cf�����,pY=�ޑ�+��I�#��!6�������0�;�$�sA�ǨT�4���7��k��k#�����X�U-��/@`�.H$�?)�8�8�i߻X���kp��[:�����;�N�A�(T�@S>�;���ld�w�ðOARp��}�&��=����&��2cӕ�Uq���6����D�E#�޿Y��X���!�ΓB��YbU���n�r:QTIi>��-��{(є�}`��18���[���BMi�U�f�b6w*p��r��xz	�Y�b-TF}�� ���e)h<��j���Y�A�7�5�^f�g��:=��xu���V�,��|��%�&����!3�� ���H9��G<�zT?��R���x)�����_y{��#��m@DGg��A����o�ٴI'z]���.R}cpn�{�65�kF�p�a����LklhX��q��w�d[�&2��'�e����\�вj����l��k�9-Å(���&U����S���.�g��R��G��:�`Y�t���x��ul�����4�?���P�
�9�}�0�|2kF�j��lkp�b0#}"��#[�}>B
�����(<��T�;�f0m	O����i�ş�u�eb=�0���u��#�B6�o�(�I�a����.�XհC����[1>_G�P&�'[�R���1W[f�4�� ��˺{7�5����/��
�ƾF�T4w���<3�{���,�gk�7�Rv�t�c��o��FwA��iFW�#tf��<	X��=�WFF�b�s�:D���񴊑Lv=A�e��flM���y�>6w,���(Y/�G�m&x~4�?�()ƺ$%��=��t�W�9JX*m����H�K��C)��5Rj��(�B;�V��\j*����ebh:Dȼ��~7�;l[�7Oe����dC��Ӹ��E���Uq-�E���w��.�Q�vQ[L��W
`��yI�.�=My���)��C�������9�ۚנ6�g�\����ǜu0$}F���/�o��@��J�r��$��Ո�DV�K�PG�r[�Q%a�l}\�8n��(!}�m��$�Jo1���	7E�IX��j`տ�L�ǣ������dE�V���1��Y4=֤k���6�zZ�/�^��P��Ғ{FDK"�<P�y��4�� o
6*�˯)�|�����ƫ�ye�����=M���RlC���zܭw!�d��T�R�֐,8����q&��a)׺BbL��X�[32��
!���'w�hK�j2f�H�2v�Z[�8��HYO���u�&�\��H���$�w�ݣ2#�Ңz��y�hI�ug�{"�%z4�-P*z��jip�L�k_��nɭF3�)1�S�@U�e��KGD\RR�W�|3}�m�=���%��{�hF�a��2�Q��&�֥{��;�\�Uvz�	 �n�8��޼z��⏖�o�u	�k[np��<ҿBw���`�Jyփ	�""E�zrS]k�I��jK[UԄ�� j��m �e���ǳ�J+���h��(q��9pu�߈n4����+��H�G�����s��~O>�P��j��V�^��d�}����"�s�/�,t4mH�2MTy⡜��K7vkh�gy�rD�H#t�jȯY/�Jr'Ɓxp�ԭx�;zI��th�/�M��V�����	@(+��P`��v�1�i��v��8'�g-��hɗǸ��#�������_]��E	�po���6��Y�o�
�V�~Z��˾�U�Y�x���T�Y{���]1�(��8���l ?�RQg�0`��(Uɏq=a��Rw��� �o�K���
)&6��b{��ށ�A��!�4Ą����&�.]�t*���=��;�gu~}��j��E�2�UBc�.�@�❴.���8P�Wj������>f4W����7Q9��kD�k�����1��2��y�A7B^L�G��ô����<����+m�i-���0�gq�@�j��I�Y �=;=�-��T �,z�Yԓ<d~�t���1umO迅/��E�LA���/f͊dY�B�?�dƨs��M���
&�}�/��n�\��XKǢf��9�Z�l�6���.�)�\U�0�K�D�D��Z �8!r�|�R��>~SpD�5�Dߨ��[p��=<��+&`� �̯ z>��ڟԬ9ytδ��57�7��T�Q����m�D-�[z�Mu���6f�1f�s�/��lA�>"�6h���F�h;����=��J�qowoD���tBk:���g�L�-8��䖜�����|�
�m�M,��I^kc��h���Wg��=�6����}���SJ���e��Iɯ�Ҧh�Oɷ4� G�'����c���'vS�V��y;SӴ�@���+|b&b�M�m2�ƶ�ȋ�=��AM9��C����_pg��Ȫih��I��Ф�� ub62�Kة3���B�V��MR��1���Ο&�e����6�"�+J�*&��3��̖��#�zr@p�R�H�Lf;��Ǻ���{nPi^߽�ǌ�2�cY]���B���/��������BBH���H��}��Ri���Ԥ.�#��S�#y ��Vz��ԶpԨǱ?�Ly�D�QIpMW�/�X�J�w�����ί������!V�u<z�g�M��뗩Ʉx�FSs�l��\Ճ��r�J�}��@����4@����7�p�c�ܢ ��Vх�Rپ~ȑ��C����Z�z�a�1t0d�Iv76�0�1B/^��Ի�◤���cB�b��j��Q|{K�ƒo2&�C[h���p���:��ߡ�>~�w{h7_r����u��[ղ�O�P�zNnE��LLU��_����9ٛ��C.E��cs][�79�I6v@��)|O��_�jU�F�␉Jǲ�P(~<�&��^J"Y���'t�����R�d�+��I�ݣ�~OV����=�d��u�jʖ��@���ew��p)���-��Q��G&�`�a��<؝����mR�K;����<��/W{N���g��}>`'U$BO-PQ�q�҆�kq+ʾ䊈���$��2���r['�X?�x�	C�M��E�)�Z�[�L��{@�ٱ�Z���t��אqS�'2�3>�)�9=���1���� �4�Jӳ=p�b�g۔ٕ]��Ԁ�F��.?�BRb�^,+�<�&�2�"�8H�٥�	�cd� ���VvrB����$̟tݫ9l�T�P�l����xH���T�T{������b�{�=�a��Q�S-`RS����VϨ'�]���ɟ���@��i:U��{�V|�Ws��o/��o��$@��[�_,��Nќڽ#(\qS^�&�.�aA�0��W�y�m �yF�GcU���� _xU1z5�XR�3~�@e��U.Zr6��~�O0���g�M���5!Ϯ��x8J�{��ٯ�΁�F��4�[���s�@j�h�`ť��A���v[�,*;�Q_\Z�^0���/�.\gytٯ����Y�2!���P,�u'dz�
m����[]�KxO���5�w���e� 4(.'��Niu�RI2�����ấRӳ��(Ϗ7�^߅�y�7��}�7E�{W�dfB�b�����l�f�2$]$�9�J�75�>	���\���[�}HQ�&^]g��4˖k^zLt�8��D�]���I����E)��.[��mE�ő5/�7���]��͑l�Xrv����f ��R|m�?l�9T��9��$}��=q8�L�H�<IX�hż�o�,��Ð`2B��`��P��n����m�6��h����{�Ds�2�6Q��w�~� N*U� @����&�4��%�E���Ž���S_���]<�0�+,`�����G��*��Ю�u�txaUij�4���?ڰ��r��F\P[1
W�b��%�t��K8�~��IlO��e�~%w�D����X6��]�O�q�L�h�T�*D ~��"������Jw� �p{�ꪶ���Hb�(1N!0�NO�`g�v�����f^�5�K�Ƚ���ʺ���� �ǿ�U�mp��������
e*F��AAC,�(D���N�ħ�	��E�@B����_	�ϲ���~�����L�%`C��oF��B��s�����Y��k��	�7����r+;Re=��%��龦Z\)V04Ĉ�NΈ�ߤ1��r+<�P�ĠG#|j-nV�\)�$wb�����8~B3�����5��ʫp�i��ڦa<�;�Ե�wN�����2Z�P���@Ҡ�g�?W�[�a9��ou
�'�� e������4I��M�Gq�ŭtܽ���Ig~����	��P���ҽw������elt�P~1D�9����I��="p�Zx�}l�v9�æ-�L�i%r�o>��O���s���L|��_��VI�����ip.���� ��{�e�K\�1�5Z����`¤�^�7�W��4u��.K_�M>X�?���p��#+ ��,C��"�f^��Ϟ�|�O�GiOҶR������2�*a6�U�Nc3�QO�w���~\�탧��ĂYh��hȶ���p�4�-�|Qzx��L?j��jp��+�]�$����㘬־C9Y��MT</�
�]�Y��fX/Z����JϫQ���+�^�"Dob�<�I���>�����	E6Na���C7C���X)��&�z�emG*d�q���K�&G�^q�5���`݄����ӜĘ܎���$.v�u��ޙf"z@��*��7���b)�%x+�B���;}���C����m�p*�9.V��r�p�ֺ��l�DP.�AY5�E(VՂ0s��1m8�
�eYK���8k�̛-{��s��0��:�� �~OQ���:ڣעJ��^F�"�꽺tJNj�Q0D
�6���,��
7��u��<�]�̟b��a�1vPA٪>L"�/����|>
!.�fv�/���B�@G>�*�;Sb������h��)�/��
���yZVdB��=��*�;Ps�H����v�
&�I(%�\��&��@����KCi���~�0'��R��m����΢6v��_���ȦB�F9s#_�y���p�!W��G+ #rP�=��7�H�fH� ��G�1��& b�O��M�#/�D�A�{	�/#U!�ܒ�՟xc��b�;�����UJB���ω��@G�B����]�8"ش�{4�gE�N`��9qR���33�S����_�P�c���;��(�)Y�7�c+��9�F���c�Ne1뼞>�.���`�!�ߜGC�:I����l�nP�tDTU��ӹXq&����`���~Q<�G�XaĤh��m:ƳF$'�ְ�
�Xc��*rn�hFG"��SO���@��y�����P�֟�^7io���1[!"�HS���h��)���Z�{h^�u��m���8�1K���2F�aL��I&�`2���HC����T�E���/W+ۅ�(��6�ֺD&�!F���YP�M׫AX|�߇��1.��js:KL��j�CR��ő�Q�;&�$K�z'��GG���#2�s1��7�O�W����,_����U��J	;{؁N��?�y�%���;���ҋlK�����j9#$^D���A��@;/ M�-M�R���?q	0s��Nh*Eyڦ��WB=���4>��R>[����҂Q���G��R��W�>B�)��F�����Y��{�T��ȝ�N�eZ,6_����16|�lpُ�.C���C�]�"�T:竾eIVȴ&دy�e����.�ջ�n խ�z^�ĊަA��pRm��^V$�س��po�>f�
w��č?��ʠ�ݶ��x"�k�E1����M\������n�@,{��.EН��C%�Nu��o.���`�,���PWX���4�x(xa�)����844��J5�Yۜ@�u��#�j:8�yw��A�v�+_�̘L�A�e��?;�䇳	�ő}(���z�vo��(�H�1u�F�g��_�(`w�a��eJg�L��'�ˤ��ǿC��${K�<�������_���f�LX?�I6ַB����D��[I������k&���9_�cԨ����b��[�`q>���.���P�Ul��-4�e����z��x���EO!��o��fa�-BSZ�H9
P&t�@)`;+D�Ͳ,������c�R�\�\�o>�H�Z�KS5�5�=5���`��������4�gt��kR`o�x�NF�F#���t��.#Fq�+w��PJ�:�2���d���_�L��E���6FB�؍�(�٫ٺ��͠k�r����ҝ6���w�ݕA�C��1��|F�fqǹ�`R~-�p��j~��Qp���� �����GsV��@f ����?� ���7,+вneg�,?��o����Wvr�U���^�G%8Jܳ�L�f�����<{�Pؖ� ���>,����p��i{��^*e����:�Zh8�Iq��#N4..�i%�%�<�K`C�ѻ�ܝ�7e��)�+i��U�j�����ւ�ƌ>v�Fw�t�E�&E�~�:�����?�O[���4�|�7�f�z���U�Y��W�~V�9�&��m�L5̝*ͲŚ|�Ӌ���S8���u��`�wn�Z@��ipM���v�-��Fh42�A�܋�Y����v#�#!BFlȬzzʇ�
��A�$���0}i=��L3�)���Yi\�arx�&>��� ���<��6�QXb�$Y:	�0�oz)���X��a�������J��K�����g ��)�^�D�u�Q.�*�_+u.32�6�)��W�kYzd�"da�Ch;� � ���v\Xc�ᲄX/mg!6�FP� �-v
��Lff��@)B��:��b&r�/P?�,B�?�g���:%��"=PR�h�H|.R�7�@��Y'�����/�Y*l�*�	���;����/�x�_�&���ࡌ�&s-ќ0x"�ؐ@Ȋ,�c$l���%с�d����k6|�h\�V..\�x�����A_���h�q9���S�N�+�eą��6��f�����e���� �~�L��b_������'}�ב��e:���A��Nr<�ҏ52M��4��1���e�W�)R�:/�)��*���kH��e�kV0����.���mZ�)Ѫ�8����t6)3!���F�F�=h�Km��,��{��`�8��Ę����£-hd��
�4hI�ɣ<��a�F��R�l��}7Ir�\�D�,A9{;�+\��׋?L�
٫���"qL=������\Y�g -g��xT�2	�_a�7I�;��/�|;��x	��6"����ݪ2�N87a��v�;�h@�� UC��hMf2��)�|E�����C1���&�ma%: �� ז�05{g��5�ӎHD6蛹ز��d^�'�������?���@���>�R[�����#�C%����Na�;묑���E�c?-k�$�*�W�+[��~���&��:��/c���5�3]\u	^mLY%�	����X]��R=����-�ۑ6�8������7�a�*L.��E"x;�a�AT^V�����;T�6M:\[��~��6�Y��~�#~�����CG�{��)�\�/��⭬�S̺��~��q_A`�U{���'Ln��BA~f���p����U��B1�)Q{7o������~�2x�[xR���d������! 얤 ���&��D�&g�R���I���ad �cH8�5��6�mS��C�J
Qv�!9�07h�6��L1N&`���pl� �|�n�xP�	6�|L�w��5�W��$}|�0����f&���$<гj�2�0�y�=���4���h�~V��d? ��)�lV]Q��=�D���ʊc��M�����?M�V�\���-j��a�̚���%\���t̶mYl�OZ�o�����n^�ӇX�|���
w��r���N� ��_�@��Yl���s 	fz�,�F5Ƙ���]���O�n'��m��*˗%���������,���θ��~��l���9n��E0_���l��i� ��
�D�}Lco�W�l��j/b�n�7j΃�|�W��yK@T8~i�� 
��jc�/3��/���V*	�������"�a��K���L������Aj+�ß�lPZ��zc�3���� �����@�Y���Z�Lދ�nY��s�h;y�{ɏ=wK&1w8ϻ�a�$�lm��)��Kk����FB���/���U���9��Or�R�Nrpm���ː̏�����_@1����\Q50��r�������hԜT��TD�y�གWJ�/��w�ٿG$43jţ���'��Dd$*<����~�!�=��le#�]�Pc$Bp��u����K�Cc�s�\T���������SS �k[b%��^u����~���F`��3{��V4��Z�u�2��B�{�n-'ǈi��"{�D��Y�W��}4A��	��+G�jߠXW|���*A�Y݉�j�j