��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��ᕫ��H��gq�f}���+����c��0�7�*�y�HXH�+��Y�Ar�#�<�k���bu�-��.���O�;����b���7pE+�������v@��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T幭xX��8�hG��kr��'�n�IK�v3�[B���fP�e�q���7V�&����J��v�(� ��n^�ӄ�`� S��JK��W�|�	�bL�Ԡu�%��x��@:���Vì�������V���M-�`8j½���[�n8��Vk���FW��ϔa�lA��v�ZMy.���M�$��K^��yZ(��E��6��y�鰦?��7� �d[B�J�������G�l���!G~1���Y"�틕���ޠ
j�
+���`k��`�=,f�kD���dojX@�Sؓ�6g�Ҕ���j�FMm�����k���JQ�����n��H(��nYe������('d!�i#-ҕ!fm	a��	�?����r�B8=�|!���L�<���hçI�HYG�E1/��Ǵ��r���j�HZ�+�}�ACi���~�|��G�v.���+�Y��Ӆ�^����Ht+��g3!;\��2-֚@�d�u�e�"`3z�͑}1�(Ģ$�b��Ԃ�Gf�s۹����W��[ij-Z�̾D-�  ������K�b{�
�Z�̜�i(Oo�
a���q�mC�|��ej��[�۝X�jƸ�`3��#P6�&g����
[^���Z��#���o/r� 'Eݳ���ٵn�˻��G��О4[��/N�2�<���kQ���49�;����`� ��|Н��5�M�����(����x{��C�"Kp-�`�x���I����� �+0��@�̗zP��ܡ7�hv�q�I2��$�g!O�����T��[�#U�������{�}<ƅ��,�d���9Y�̜m�)PrE�n���l�}� \�ܭ��R��e|�����b�C�̺�>0�{�d�7}-�f��\���)�K�0ys
@��zG�ϴ�=C�L3����:��Oj;�hS��^Z�E�N�}N*�&�(�ap�Ż�~�̊�C���E(>Wʣ��ҕ�6�8%+^v�.�kb��.,�Oǌg�;?��ܟ���+������ž�R�P�
]�@���|^�"Q�����<�U�m�Z ��I��Ak7��=�o�A�m��y��I�C[_'�^������G���e�G.,[^ز" gN���gj�l���'�]=H������ �Sr\׸l�ʯ�cUі;s+�p`b`��O�l5�A#�J|��� �j��Kb=AL�",�ۈ��W�l
]�h�Ԋ�m��l�gJh�_oeX�~��pj�V�C�?'}�S���@�ao2V�X�5u�eJ�kȡ�|��Wh��i���x�E������+K�X�b�5Ъ���C�<஗b�n��?m���q=C@���*P�Q��Ũ��Ë����~wܮ���y�Km;fś�%=}ݫpP�Rs�d��4�����l"�K�B�S/����u;��t@���'t��(�j$@��>�9e�u�T�	8�!� ���giE+ÊٛC�!IU��E�szC}�ޫ��C������,7H�G��=@p��@�o��nB��n�#%6�s�DRxV&��N�RB��˒9��g�^*ͥ��v[��:!,��������p3`�<2ٕv�g����s���rIbq����wW�X��08 ��[�us�_��=(��(��	+B^:�D�1ԩ"��aH#%m��j�9L���E��mS �F�����F<��Q�h ���:z�B:��U�<a[�_ƄM Ŋqy�����qE�f�n�"r^ݳe�<$����l3*K�N�kҥ�+�>*5Ф�4k�CZm�s��Af+���%i�c`Y+
�����~  1]Uܖ�Hgo9�6	�Ñ�Z�:_B�A�6����Ah�� �ظ]׈@�4�d���Q�����I%`�n���Y<&��簬����V��pL��z�Ч�_�)�t�z�Q �a^&��i�#9 l8��&k�P�K�K�m��S�|��=h��@'L5dp�>�֟���s:1�l36�g�&ή�!�s@i�X����Ȅ�i'�U�"9�]�s�N�V��,������=V���3����?a=�t��<ts )�}�v Ic®�iv��'O�-�t��Ȕw!@KG-�9m�ӕ�G@�^L���1Wb`2�RCsg�B����?�������c\�:�qY+֨��}����+FX�a(�l/�s뼣H t���Ìi��D)D+S�����洣b���� j�s�IO����xt�BY���Լ륩�UDC�Y[��\r8�{,�	��r�"}۔@���#�����w-�^uMYAnNk��#?DWRt�8�	t���Ȇ�	�]�^1.��@[XG>b��i�ŹR	����,��������F5(ЇsR��ֹi�݂f9rMBJ�T�*����.c�Q(�6p���
k�m�k%�)A�L�HBS5
7`�]�֧Ƈ#��S�����}�~!�a��ϓ�8n��m6 *��Q�谗��\QlI�G�o���m'ͥ�0��ޢ���28������u_����i�����<���A_Mф�5�o�:ex�c6MՉ�g&�����F#CU=�uT ؐD�K�Gl�$�H[gy%MyȚ��#?�6���nVMG���i�<P��W^���t�/㯡�ql�����M,�#U�伈W>��������e�j������䬢z�`^��u��"��-��<\y�B�t(B�qb��S���2�+�� 0he�#���_���H�>P�7�y:4��P�-���#�,ʌ� `}��ox4I�6�O��W����|���̆brAE�Y��)R�'���KH�g�]����R���|�.������.�K�O��2#8�s蘞\��1>Y���\h�֎����>2>	"K4�Z�@��gCr�b���
4�LwD�|S���L�k�� "5�"�	 ���ꏇ�Fra����'���Y��ϛ�u����=I�<�^�v��z�ba����c]�b'T�4v~�����z�!G#��e2--�`��L�ŭ��K�"��rg&=�����Gn׾��������ܶ��C��;��Rl�T�Y�O� �q�I�μ�t!o8�G������S�Z �KL:��(银"�rcs����s��Q;t[���$K��,�2�%���eQ�u�Y�{� 7
���+��������O׽�z�תz*'�`_�Bv6�k�S�b&����b����)���\����GD �,cϕ����[M�{a���5)�1���1�����W
�_��)���&D��~����1g,�YY�`O��g��oB_��;��w�����|��a㘷�n�������u���z�L]�o���$.C-B�a��|�CMI^	|M�<�9��D�o�õ�1���t�&�5z�7�>��,�(�M�Sȋ�M�%�b��Ђi�{�tJ����s��������j��3�S"���0�Ѳ;���1�YW΁6�7T6j��9:R�ZJ:�K��uX�;��5�t~������!��������O���B�$F�b�$�$�j� ��	�=�@��F�oG��]ǕP60%��5"V�L�h�6���{����I�I�e>�3u=���ѡ]=:���'�rj�^p�ʬb���O T��Cx;����X%��F ���IL#QV
>�QU�ƧU�4��ۚ��l�z�p�;��=,�8�l'&]��g�2�w�ݧN�Q�!�r���l)~p�WJbs�>Cu?#�m�-�ŧ0C�1���5�*����\޽7p�&�/��$YT�KCK�����6!"`�l�`M	�f�yW.Զ�vy�*H�S�Ŵ�����2��ϰ���Ei�����.p�3����_Y@0��g1X����|r���!���ٚ�m��F�ߡt�C��&��~��\���B&���߆��������ي��̈.1�ټu z-�T��tT㚬�T����q�8��� ��y���!�/�mSq�9ND��}�=��c%�����ر��j�tH���~�z�
$W`�)C�-?Qp�m253��@��-d2S���w`����x��U���Vt?�!�I?n�@�	8b����I�b �U�񁭃�>�;��>/hI}�v�=/�@�v��R�9��ة1 +��80�;h	�3�1�.��i��SU;�Uᯉ"��f��U�C+YZ�	�<�G�����I�-����U#�����I�E&e8ծ���b-v� &5�Cu&�zQ3��ۊ4��P�������ygߦh������j�� *��ҨG�C�>؅���J��=�~
,���'��Z'j�s�v5fz�<�c��:�6��[�6�L_�^��ѭ��*��:��':���rP�)��<Q��!��l�v�����Ip�"
4I�ˣ�!�pp���C�ո�ȯC��������?mC��f���c�n�����{O�q�m��~�5X��#��d�����Z~���
G������IO\"�2."�����
�L�gÑ��
�w���DP�x���@�K�vw���#j��}�3@蔽�u�d"����KS��d��i�s��)k+#����f���N4��>��)z�.�ߵ�r;�4%�"���J@B��偩C��}{��EV��������}~�C��-����[����nh��v2<C��	��pc�νk�9:��#�$_�4���z6�1�s�R�;9oYɱ{�t��E��v��!1�f%KYO���|s��Gx�'�.��Aqw�'Z�Vn=/+z��U�[�g�O#����%�4C���)n��m̪�K��N�Ze�����$���J^(�Y珟{�e�ԴÇC�c�/m�D'^��;��4ZcG�p$�<P�ԸR�'�y�kkب&��o���dƍC�c{���k��|��<^j9ﰔ'v�2Ї�ʰ�9A�9��`�#����H��ߚEmV	Dք�4ͥ":�	U$�HG�9�P�(9|��5�P�.=K�{�Gz���)���)��������9��Mē�l� Z�gas�vª��F������������89A�ԥ,�6���-JyQʜ0��)#z>��o���O7�>��ZR���I��#h�?
`�T�v��@����?�<h`����s��a�<h��)Z��d蠶�b!�I ԭ�~Ӓ����~����o�0���zn��l�M'�K������h��@���mōxK�j�c�~�_�@8�I����Ė��>�G#��y��-������z�V���dȀXT��H��1�ab@�}�D�'��� ���ŢM��f󣎖nn[��܃O�,�����;7�W�a}��KbM��s�*'���&5�9.0"�� �7=�Q�K�HI�[���gmR��p��!�s_�ʫW��Σ�Q���Ҕ���6[>� >���?�����[*|d>-�X�tl*p>� �������Z��-��ܝ�z��5o�M���~�Y�V(��!%�E9Q�����2v���V���Y�1�Kw���d:Q�;l<��Q�S� I��z�%��	6���aû�F���Y�$��yx��!K�.x����M:VAW[�C�����S�)�ku�`���I�%>��C��l2�	���}X���O�R�&荖{�n'���L��#�.	OSD����O���ć��g�b*�l�B��\�����������,U���w)���x*SC�߳ukӸ��:!��Nev�6��}�0��ZK�0RFcZ�Ü��l�Lu^{�^�.h3Ήl<�(�[���I�ظ-)���E=R����#�PtD�kt��L�Qڃa�W~;���nS�˚�/^�I���B�u��BX���0����K�/~`�	�d�Ќ��Xn�\y���P͗KI��(�E�I��G��m\�o��6��U�ANQ)պxI��YK�
��ap��~�(�}ѳ��q1��&���[��=�P�ů8��x�����м@�>0f�L��[&W�����	DAF�t6��_vv�1E��<���<�^��@L|�,�~H�����G���֐��7'w�b	9L<y�Y���p �C M0��G��0/d�q:{��7�uv��J���g�u��*�u�k_Ŝ��]�»�!Q��������H�T�e�y�^�t{�UjϼJ�K��N�#%s�G,&ʨo^���qb���3�aҋ�kw�����ΤVq"�U`/q��^�7�7~(|\
����f+�©_��
���.��d�Q$�ND�n�\؈�>I�.)�K�HZ�P�{�w���5R�@���	��β�LF�l�ⷾnlõ��hklԥ������?�h� Eo�/��H����H�?�TLO0Ȗ]�Sy0��G����HӉ����
�*z�zGsQ�l�1c�$G�������|�3*�Z͹�	i �����FO�	I�i.����H�B��N�B%O%.��~b�G�S����b?�$��F3�#R�E1� ���}(#�� ��+���89`��t�+`�#KŰ��W���4�.2;3Xx�fWې���������bह���� %4Q��ˡn�N�u�O�l4�Z�B�K��,e�5SHE�7���P�o�
K�ң�L+__��	r�d����#�R�nw.'��\��!�F!�꡹�HJ����p�@�$uuj�Ś��	�vC��z�Hр�UQ��e�H�"�*�����!!cb�j2Z�������М{���CX�����M[zE�q8c-�b�r��߲�Ǚ����W Xۓv�_��>�~���m�rW��3�-p��70d��2�ߥy<�����F�6��#��1ÝP�W!�?�;~�M�e��O
����?�8���ˬ�u����l������Or��SB��%N�z�z�"�`�7�������L�?�S�,V�����
	|���⌽������Gp���r���֝F�"�eƄO���ߏ*����Aڍ�z���uԳ��`�!.��,��RI?�Y�H�x�lu�6������֘v7B8������-M�/L# �'� )+x�,�֦����
@s�)d�c�{"�U���,,:=6��*`�X����A�̔�P�tW\n�f4K��/I+��ܤ�w���|�cN(>Tzk��w�z��*��z= j]3a��� ivt�R�q���u�K��!鬨��#2�&��R���*E�+�Y�T��F��>cT��E��aS/]�E���W$?,��v2�l��o��ƀ�4o�y9�����E��M+إv'�&���M���Q9�dF\.�v���ۣ��d��!$G��L0K��h�J�'�}>c���c��h�WG��z4s�7��K�}����S\�Y!2���]�D�,�"#������O��η+��U����p<�B�,�_U�p[�mB�j�#~�Y1�(�	�C�ե]j�B�`�#���Ex�k����u�il���uVÂ,L��+�\ ���PV=�&�����-(]�L�ne
�݈w����7ȴ���<"L��NwA�l2�,�����^fާ�3hi~�K;U!��:%����p�ϓ�B��I(����v��<����~7={h�ae����Կ���=�ꇷ��-#��<���kÑ�}�����DA����H����EU��Nҵ�4cϱ�q�)ep�`+�=: ����i���g�ƐXae~�S
�6��M0���:.у������]��h����Q��6����	tэ+=�x�o���f�[L�۰6�!��di�V��ҥA��[V��o��.wݑ�ʺ:��U���R �?׫��P�ZI4Zu�?87��z�3���-�i}���xp���J��rW4ǭ�2;�����Tl��~P�v�]qi�]�(���8�d�Mbeq.ۿ��«1ӊj	m�����<V�D�Փ[�%4%��J���E:q��
9�]!T�zr� ˥�A V���e%� �d�1�5K���T��-;�'N��ύ��x���5����OBP2�f�=_
%��t���X@Ɏ��K7{�9�@�w&#c."y\BI�̏C{/� f͋;��T�Mr����@��@X�#�>y�B<�y`�N�n�V���K���(�SR��-�L>�|�Yh#�W�3�a�� z�j��7@�AI8a��s��d���l	�$K�a3&�`$�>���x�윎���Ĩn�����M����3���ֿF���@�����9����#�At�/��0̓m�ĳ��-lz���= �wM-!�鴁����GFX*���Ix�oA5U�z�k�ړ|�KQqY�)E���~�~m�"c�\�#�<t���[H��G��|��O}�Ib�V!6+>RJH0�"�ʙIj�9HK�}�<�_.𫸡�8[���>;R#puT�SG)�_W���	�a�d��ql��0�+��Ag�R��j>mx&U[���ҹ��R�Ob��Qչ'��ܲ�JX�^m}N�����gz ��*�*�mMo0����(:��8-��Ϸ���b�M��$�J���FwVe)�¼G�@Sӛ�rp:Z��8���'	�Ww�\N���'�I�7fŅ��Vs�X�D�0�,��+��rO����7`r�w�	��?|��j��F�b��q��~��+�S<�N���]�I!�k<�,�N���j�oK!O�@fΉ����U(hU#�C�����=5��;gv���������T��$�!v��U�#
q��O�"���9P�%�ʈl�U@.�_�=Y/�s�3���F2�["�7�wNj�-ۜ�P���v����i�/���'&(�~���^�NPM��x�è(�}��E�x�ުSNB�?m��S�Y������LG�f��OqП�J��fފ�QO���H��m�X�u��<�#���"|���>��"�`��l�s8e_������� �O�i^X���=Q��k'r���K]�-+)`����h �nD2�W�r���KUx���M��O�Y��8u�C���&�$V^3-����	L�x����7$t�kp�S��ج��FG��{k3 ���
�%>ϸ�q�vK�Rr@�t��#�e��0t4��h]�z�G+��_o��
	�o_�V]DU���gDS��ʔT-qbL��Y�6����j�q�����~aޞ>K�X�ū��J�]1{,�FQjGԘR5��RG�P��S�Hb�c|N���bo�Z��L�D|w�`9 #{'���C�ZU����8�TwM�>	�ܼ��>��s�e/*����������α�Ŋ0�4oH;����3�C��L����A��18��C��<7vLmb�j��`:�E}Β���������n�@:B,Ø��[���$T�6���Q���k&I�RUE����}�va7)�W�E���?��AC#I�V�����1bP'����/`�2��	�9���=��gy����~�,h��kQ�z
������ܺ�s�C�()���#�F��Ц⍺N��W��g9�����,L��_>_�8�āZ9���Զ����*�!8�Ūu��g�	7��!��1\�I�����,�'!P�|WH����=���l}��r=}�p2��1@g���J��r�s���%[��v;.����9�dv��)��,C�,�Sڜ��ZQ��+����[х�^�֞���=��6�q 	f�]+hl(P�z�Y�_���6�)��W;"�t�} =��E�A�3��ZHJ}��v���G|�Eºf���c0�-*��9Ц9�F�Kt kO��h�[�>|��.gR,��̓���a=�ț�(Y��y6��� ��+��]!�~@G��j}�4���{p`>͓ ��r`0
����[�Q���ν�@E*x�3�O\O"Sx,j��o�S��
�@ ���?���|"�$�����6�N٪�뽣3^�_*~�����~x�ٖv�C�.��W��b�"�E��'�� ����Fr����SҦ�׈������#�N齠!Ku0�I�t!Q٠�n먐Gp����gO����n{۠�>1�e*�ۀI��Nʶ��ȫF�����Y�(GT�*	� ����Vn[>���B�HQN��C�ٱf�^̡��:�pB��Z�z���^=:�=&4�l ����zv���ǠV\�֢�_��;�Wh��S:��������%�]w0o��{�[�)2��'��x�mU�����T5~�l7υ�@SQ��&���̦Ʌ7j��]�oS��7�%���KX�4� ����`�މg偬�pm���7P�G����[�*&au�(P�����!�Ji
pU�
9���W�Eb�d�Γ���z�xc=�Gr�<��T��
cVv+�z����`��(�������	�3[�o�EO�UN��݈l�AO1�IzKe���Mݞ?�<���̰,BR4�EB�kp��E��D�:\Ԑҡ�8�+�T�e�j���n��cxRK� �t`,�s(�Q�E�Z3C����0u�X���
�'¢�j�SE����ʝfݖ��{�y�%��5�~'S$�U����T��Y�h�a������X~t #��X�H�<x��[x��g�]�[y$z\�N��l�lF�����CSk�Jz�V%D茯
���CI�,%���D�{I]�%ѐ�8󬲴��e��R8sQD�D߀7�>�y@ގq��xM,^CN��$���>ܭ^�;i�ze�ĕ=��8N�"nq����/�)���5�|G
1�G���90�\��r[u:=��}��-��(t9qG-C*��bu��r�������Y���d���;�T)6Uh��b�%����*I���0��#�_ꤹ�EC�9K��n�D�UwAet�.���Qr����&�?�B#�N�c^>��%0��s��s�e�HM�U`��NI�<�����0W�����ŉ��7`l`$1%�i��l�hy���ޕ�tE|�m�8��+D�@�{h*w*�g1�����u2��� KӞ��pzmC�ϥ��K�r�\���� F.I5���D��Q���`����`��VW�B0]����\���N<MCQ�Y�_�� �7J�b���Gֈ�2,���ȨuɥV@oL�OGG��Ш�	˝=�����jv�0 �!sݴ(��?��c
�)��y�_}_e
�f:}o�qwo��o���r���,��T6Mr�����j���۰8ֹ�a�Q��~AhV��[%__��\=�����)��z�QP�CR���w�#�p���"�0^j6��τ�y)�0D��ڠWd�b�v�Bp�uƠ�=�d}U��H4ijc8!wK�U����\MmQP	�MN�P	SRW ޺��R;�`����p��O:'����-x���y�U���kC�G�&�Q�y
��@����p
����d�B�@:Atp��
����]��;�zW���A�ӟ��:^�]x"y��Ñ��>��6?��u�j�'Y�*��uGM@�$=_F�3���P�˸��(L��G����Y3�%���y9{��i��O�k�f���q,�
As��W���=ȓ]m��G�OE��t����JcӇ�;���>��5+�\�}n_��]Ht��?��彀ݤ�r�ݪm�J�l�.G���Tϻ�F���������6W$%�Dc��1,�d�}��/��[��^�_x4�G&7WQ1�7�`K`Zf��[D�I�@}����eO5I6(���z�*�+��������������l"�4@��,%t].�� �[��'Qt�g�SZ��ب)�d��Y�ٹ6(���	�w�!�o�t���C��٣l��������GE�T3v�v�!�.�C+M��D������M
�n&�k4����eOh�1��U��vNXg� �x��)���U|rŕ�aT(�:�.�nO$�@Rc1M!�H���ɻS�}α�B�9L�p��]�ʆc�?#���Q��ٴZ���R�5y�7��H9G���t���t��x$C�}A�yy?B��P?u}i��/Z�MK��ގ]�P%���o+���$	~���dVE���ڛ����������m�]�^q#��ZSUG5���<�h{J�Kw$�L?�hՀ#i���H<�s(��P�]��y+���NW��̸��q�id�?��Y������U�N(TW)��1Xc
J���E�A
�~ڗ�1�0C���r�@���X�/�"�uty������2*��-�:M��gO5^t;�+MA�p���:�F6�_A��AE��uA�f2Uc��*u=9Ya�>dH��&������i�R?6����+�)��z�197h��3��[}[g������8 ��c��b\���r��J+'��,z:���dM
��;�� A�O�΢۲����᫞[v&4��wϾ_3=
a,ϓ$�~��7����mAş*�T�;ƕp�L�$�p�`�<s6{_Pz������6�eؒ'�Je��W�9��.c��l$�=���*kec��7lB�ThaƷ����#�����1ٕ�D�8e����(�r��T5�:�PAJ��:g���!?/�̵�uė/BbTQ*Q��D6��Z��'�¯/+�j*��58M�f��X�I��g�<�{������C��2���k����N��0X�.k�4�:srs��`5�7<~�O�(�:q-O��-�e�w <#�ęz.[�K�KyE�FH|�
�pb���t�Ԩ����p}?��-CV��gŬ`Lq�z��xpY�y����I�gU�H��,h:rP��J��Ȃ|��S�
�y�^C��jyIR�$�:�ky���V����hK룸����P�Ь�.���EGv��705Kɍ8ҴlL��p��W��������{���-H�
u�w���o#$B(jc���Ce���r�6p爧b�Ѱ�}�$�{�/���A���W�O[i��%��v��#��9/�C��<X��T�rֳ4��d�iC�sQ|>�hŚ5�&�&����:Z���ٍ&�:ֱo2y5ŵ��}C�C���ee�d�hcl��9��38L��E�)�G�+gG�X��{�ղ�f�n�A��"���P7�7�[1�D��=��}҃b^��Q�`�#cRgFleQQ�N�/��. r����+����HǾ3�;|��#�bDs�d���6�(��N >��g��B\T�鸊���`���~�"���~��W�:*��j��v��t���]	���HZv��p�:�Hk㲕Qu�T\�%����ȝ�ݳ��puגb�7�!w�
��&�5�f_�=sbA}$��Z�.#�r>>����w�#7xB��*����0/�Ŀ��䶀k/̭WyD��T,|��aSĝ���R.����L�'��z $�[�ܑ����5�4b�ͫcd�~Z$,j���0�h%aq.�$S�/Ժ�|���*}��Yw�Ro����vT�/�JÂ�I��t�����b[A��O�R��h���� �P[&{ݥ��{���=@{��,��CO�(���ܡ�}��ˈ.��i$�q�dE�'�SQez��֙�Z{��P�)x�D�g9-V]��8ԋ��(����}��1�U��� т&t���~�c��@�j*F�A�A�c{�i�`F�o����C����}'�j��������7��T�u���ap�awE�av��&�$�\���K��*@�1�(\�Zu[�,)���x���}�gF���&ⰽ�Y�s�r^�����z}��X�/N���!CN��CB���r��V_Q١x���q�͍�>�|��_H07�5���+�y�&O���NF��h�8d�P�m�}5u��Ӏ�
"w�RF֙Z�ɲO,�|O�6�;��'&�O�K�I�>?�#�h��R=?%���N��'��f�� W2�Q���%}
 ����x����L��J�����#Y*��صI,���$�g����Ԟ����ʠ�a��yW��㛡`KJ�L��_&
�4���h��%+�e�<Z��uw�j��ol��n�sҵ�����C�x����Jq}j���P�@04˩6�[�3Qj0��%2��Q<Ɋk>���)����E�e�N~����dYy�����e9_�9�W�)2q���^27�>_���f}��d~�W0��\���W����/}��uMC�z�? bKb��(�%�æTP+JY��(ތ�gL�Y��n��7�	C�(Z����x�
\W	z'b�K7�Ch !�������9�ֺ��\��qa*�70��5�а����� �*i��|��xR��΂��w����!�$��󵳐�c�8ܐA.�]������u&��RP@Ԭ�( ^�.�Y=ˈ�VF"��XKs"l<�����.�8�P#�z﫿���[)$'��ͨ����y+ �E�">Q22����$/����.\X��,D��� ���\^����i����������B��XK��I��� �h~���}lpJs�KY��^:I�������m{I���l}y��Ćµ<e)?"��
��/8P��^ٴ��p:Wjqu���h%�����U���BUloOn����5�r���%���M���خ�4��<U%�D.��>�" �љ3����n���%,Iw��`][�܃Z4��F����@�t��8���m*��<cA	L<�ص|2�L�������(]�+y��t��}7��3i��[�+h������n�ᶑ����bg�v���[�=�-�W*��^-�۞�?�Q�����UL��)j)�cI�0Hi���b�������٘�n[�Uk
#�t�(��=.���+�5���%VE�*,��M�z;�i~X0#k��{F8ݼՃ�~+����mx���PO��>R¬��e�95��V�f"R����M�����-"�f�$�-]�R0�P[�,��r�8��+k������ݙ�m�@�H1|H�k�%S���q8׼��x��ʤ��.�5�A�/��(;-pӏ����<�Ȃ�2�w_���?٤J}��V+��t\%N�6*<]w2&���U��4Ɛ��"Z��{�UHW!�=��Z܄�h�����IEL���1Z5C�a,��6��y1ƶ���}Y�S���>��`|FJ�{���n��+/l�0��F!�fhSY�!
*;�g+�.�p�����+�wVA��.���x;S�.�����(K �Y��k�y�,>
�1�Y�J����ڇ��>RZ<�M�J��)<D�#��
�X�Yn����㰮�)�:�!G'�C��
�)�s��3�\���,>�W4�������)��k�2�}�zdg�g����������:-*
h�.M����`����ɐ�aA���!�������r���{�$�?ݹ6�!!��o5n��,K����˷jފ�2Nd].���F�P`�D{�d��-���2��-�:L���p�A��i�M���K�M�X�'/�<hf|���h�<�W�қ���5�|������ uk�?�'��e�k��x�;��3qimr�&��![_����5^LՇ;W�k��jZ;i�C��1�,��3=�$;>ZD ($���7"9TH���C�$�#���!����
���jI��W�n���^��1B���ؖ1h���/G~��q��Bk,�E�u�)e�O�.�\P��{�{T�oj,�}b#�J�(qRM���RmB�3�m\@�ѷO���Ur\�HڄD�76Tw �J��z�n���q��fi���������DW��������Km.V��2ܡǹ:�=;C+{f�=��ģ^���j>Br���(p� HAD;�uІ���Ќ���6��H��BcXKH���l)<+�`j�k�%�����M7� Z|q��I�A���e恭*�������G�����%I��E�e���Fk�#=��������F�T��&���E���+�z�&?����=��6�i����.�}$���lUs�e�:{�,�����xQ����jIގ��hq7�
iL��>�x����҃{����9'\B�K3s3����1�I�q��vWJn�^����z��\@qZ��J�W�"��Օv�r�9g����8,*bL���&�[������KR�
��^5u@�����&d�JP��f>�3{l�����Q��L�KEZdV��y�V23m��]�z?�_�֯���+�ؿ���.|�a�M\K��
�dl�aM�T���o��F�-S�F����ߜ1~=?T��e7�?�l�w��a �7�g�p��%�M0�]�b-O��K6�Q�*^j�I��;�̍�iF+��kW�n�d.�	������E��F�A�$O�}�X�-5����6R��]ƳH@y�0o�)��g}�����?@�r�:��Jc�r�>��-���y=3�p�~I�/#�3�σ޷"��!!s�㭙�!ܠ��2,UNg0�0Ϛ�F�[�`����>��y��B�&�	����������5��{�`�l�,��	�;`}��~���X66�4��+�6�ꓮ$u��a����=[]:�D�iy囯�CY=��[��*sk7��?Sj�g�˲��:	³���x�v"Y��0m.�@�my7s�%�I�v��(���}I���&�K���!0e�{H��<�dV2]K0 ���s���ī�]9�Xb�d0���Yb65�>��5�e��IW�@�`QQ�?��7;�����կ�!�Q�[\��9��\���u�O��"�||��	�A��T��D�^3f��o��S �����V��T���f�$p==�L�(������w�D�0B�;���<'ǔ�d*,�6�2]��d�L�������H⣮��*�z��T1 �qo��D�-\���鬗:@˷`	T}1<�+4�Mai?�� 3��9��%r��v���i��������et~��9��&�����ǐ�K�bT��=>�a�|�w�I������!cƹ�r�j��5�^�*-� <�rJ��0�BU�߳{��~3����{�b����R�N�%ֹ���0��<����mT��(4�~��c`c3�-�x;A!�f#8�5O.%�*n}B�����~.���M�}��T7%�Y��8��U�sG��LO�+�h:�[�����*�f.8��7�i���G�H�U�0���ܛ��^��^6~��m�e⢒�X9���y¡L�X�ېS�����喵�)Ģ��E-���{AU���{X�`+mx���Je�ح�X�\��L��M�|�ӛ������b�˻���:�n+��QGAY�(���(d�K7�#�6���W�'��.��!M��祗��S<����]Q���
���%3��H�Hfy�a�N�2]r�1�E&�1/V*�7P!*^v����T2_�/*��z��Sb&
8I�_�M�%ƿ�~��� V����NڀZ�4!���P[��4^�]zmḐh����t��\��Fz�l_j�|Ru���q^����2� t��I`��g}mAp_9�)Bf0\~`�W4��Ԉ����O)�M�\�٘�,�u9�Ob��hD�y	���{���+�u%إ�^���}e{���|o�)�H%6��1��"ຎt;,v:M�GG1M��D�ߖ�Ӓpmro`��oS��Q���.1R�3�#5A�z����~��i[�:x�����?N�F\���X�<V5��@�90� ��C�nLl^�ԑ�г/+xG�sP�t�G% �VFP+�,Ӻ�o�=ؘ���*�Bu��1Z�v&�C�[���=��m���*��L@[ś�o�ӔN����Y���b�lqӑu�p�'a�͐��l�<�Ά�*<�Wl�<��Y��	ϝ��\�8*P�� D{�>b]#��yu�N�ܵ�;~8��E�|07����&⻶%����qo'�%����	T|'�ğ�A4��٠�����&�-�Oh���I_H5,�g�;��7�A�(�D$sW�T�6�_���0?š�i�o ���՛�i���	��*�l[Jao:V����e���g�����L�!bTó���_����u4��m�&x��Sƒt�����~]VN�
�'"�[ W�������{�Ǐ��Q�����x@�OÄ K���Z�p�ar�C�-�Y�^F��S���ڄ��8�b�͹�׭O�9���31�dO��z�ۜf�i;C��p~8p��zb�8�^�f���PN��
"��`�/2�E���p����O/��,PM�
����*`d��7@�^�a�LD]�R_6!~u5P�+M�-�#Fb2���Ǜ50u��t3�
�ԃZw#1ޏ$���A�*'}��Y��U\�8�!t\9�r��(M�Xf N��P$7���S��ݴ��m�=z)����{�Ja�N��Yu5�mՉ�u���>if�P����f����lM�%�K�:ل6Ճ�[�zRw�Ȗ�s�D�oß2lԶ6OL��S�j�Z�̷���:��W�ڌ9n�v��$�;~	�BY��9m<�=�N�S$�"�.��9�wRDP1iP+�	\��� �N,��@���o���bf27:��8�#F@���1��G��q����o�Ë�Xp�;�p�<��ugA���{�8�m8�,�<���RחS���tg=ɶ�
#����z_-)�y��ǹ+*�//.��Rv�`K��6�~ˬ���I�d�*քޭ)ց���\��S�S;�S��0��vX��9��ӕL���T�{�c��@W����D�Of��e�<�&K����Ͽ��h�[���'�֕=ɂ�N� a�/_��A���0�[�QE��Φ�%m=�Z����
��w{tDK��|���p;�� �Ia������V��ǀ��0C�`���d:��9����P� ���n���[���v�Y퍎|Bڗ)���8�A��Mqv]wI!X�r�z�قa�h�u嚟�t��|�Q�.wl��l���ç�W:ܰ'�<�M��~�T�ۏ@�c{v��.V��������]F�J�Ќ�Ӎܬ��W��mb�Qx�F_>�ŖW,wyJu���+ �q�>W��(l����ō�B[�3crO�4?��V��T�bꊏt%��'7�vT�F�M���LJ��}���N������T�S-�6/���;_y8��6a�jAq��bl_C�n�KK�y<�O����,�U����E�<
9��o������݃���Oᛥ]��lD+I[=�5����6n��[*G��}�e6����v��U�9��O����,�}�2�1[o0���w�ͬ�X^E=��9裲"D� ��D�(��s�����K�z7���W8�ҫy�:�$�W&�^�lw��R���.�?KRɾO�6�@KU��u���YLN,
�HoI,�����E�G���~_l4�	j�=���u��������X�<Q�:�k��k\nސ@�r�z��8��\W��8�c Q�<QW}D���T;�g���,/���~x澧���2P��b7E�f�<�r��+Q{��B�X ���&��sQ���3�d��F�
��ZI�r��:T�o��'��s�&���<�E��u;㳡>{�ݱ�q��0o��d�Da*U-��d%Qb��U\��9��`#�}���j��:W�v�ZtA^� H?����e#c�H��t+�#�ê6�'SU%�*:<z'�ϭ˂#�6�'�oukv~Ӵ"Z��ՠ������ mv)~� 2wH����~ݫ�g��Uv��vXs^�M)�~)RB	�<{�J����&��wkѿ8 9�t�p�7B�A���	�a�$��	�Q����*"O����\��Z��,^7ܑ]
g�ޔO�E ��o<Υ�P�+����("$�>��R2P�nA4��/���={��N�Kw�gЭK��H�!C���g7�!"��]�G'ԥ6�G�Ƞ3�턔O*�\��+ v�r������{=7t��H	ħ�v$JJ��t��ǜ$s%'f�(!��6�Tr��cw�LSb��O�.J��G��e���C�z־/��K�4L4��Tuq ��8�S}X_JpOm��Ӆ�}�3y�:Fl�������z�K����[.�c�=�:�k���>��@%��̨u�'C.�R9f�]UW��{χ6y��P����-���u�kk@��jB��l�N;I�,%��4~?�4}�L<�	�f��y>q�\ɋ����Z��7e���rzݼZ�SӻTx�qt����$�H�v6Z���v�>�)�{�x�z��������9N�Y�6:�&�Y��~�f�N	b��i���*�+UL�ɡ��A"��d��+iZ�i�Q&��Wo�=`�]�C��5�`�@��N8��P4��_���e#��OO���V�;RӋ�$�II����<�IG$�����ݐS�QOI0��4Pp��Du&
z(�����(^��?��l���>,}L\d����b�L�W�'�z,�F�>%�vN��K�:��"�����d�Q�Gov&��E������
�&NV��?ͷ� �sȲ���n7���_�.���ۂ���Bmj�2�����C�!)�Rau2
��`�{�x'���7��ʧ�넵�AS�t*So�8�i���Z�`�W���@�N�X��Q��+��|���!�ی/���D�-����ɞ7w��ei]PT
5�/�]�M�n�}pYh��/��ܺ�b	��Ϭ�)9j2f����е�]*���4,%�� ��=4�a�bHa_9��Q;Wy� ����,�v]��t_��#����ɔ�ڎ��K]�c�gka�DN�?��6�VJM��!X��[��@_��^�=�D]=9�:�}J����K��R�.d������wrM��thI��t�3g����������p�B��L7'�_���L��ьb&��&,�nT����X9���E5��~G2��{��ɷW3���T4�2=	B�4:��Qczϫ�d��k��ɘ��'��h��94�̢�������ߋ��WlKɼ���oeA�!A���  �j��wZ�I�Xy�+�4���3}�-�;�%��Kc��cW�D���罷��[��o�	Q�4�p�S��ԅ�L��w$�{#����E�-&ia*�M�x�Έ�����)_'
ސF��:��5�"�`7TfNv�(���Ug����|q@T�����*��h���]c�j��קڍ��n+���qf�iP����דaUA,=�fČ��G|EǉZ��8f��V���E�	���&3T������G��&9g�u9c��({�Y�Ϭ�[eD&sJ�Y��gZ~\P8�d�b�b�oV0��!�^���@Q���.\��C|�ʴ0�F�^d[~���`蘍 w�dWL�~��r����v�,]�A!#�g���4�©n��s�P���ZӶ���r���[�(�e��u�8���W*��7J9�t��Vz媰L��p(�Vf}��e�B9�$+�kE �
�;�
���Fa�w�����&�P�ڰ�Rfޏ�6�]��������Nn�6���P��|棢S��m9������̕��Y�l ]��<X�+�9������,��v�B,��,��Dbٝ3�����Ġ7�e�'NX��bO��S���Y��LG˙�'������LUt��#]�v��{�e�Jg`m>�)b��;���g����	�%J��S"��t�`�ـ����->�r�v{��Oϒ�<H��(���y�ಯL�}���[X+�ns?�P��d[p�����~/I�܏C��qA�y]!BO@r���Ff��X��T)#J~$�h2�[���(����iq�fNM����\�<#C�D`v��`�Q�i��R��lj���Z��Ǖj�y복�c-�γE�IE�Ju�3�^���=��"DQ�ݣ+��SHѮ��F)�S���D��<d�#H���p^�on�$#֖���c%T��G�PS� �ڥ�A���k���2-�(|r-�;b��M���ѝ�7�~�)�5 ���ڇ���=4E�%��r�;wa8�S�A5z&��jg��3��=��rR�����@!*� ���ν��<��q�������y�
�y�r�3.%���c#�3��=�w�;�#u1I��2MP����*��	���q��N��I%���E$��h�S-�vSЬ���W����ND�^�?���:�7��Z>�n뗂����w"��Q<7�@�SQ�`�@c�'����܂_AbQ���m֯=��BIq��i|6���Ňò�j`"�v��Y����o�V��(֌n�i�Y]*�.|/��ζ����-��V�[��o�o>2�vBn�0��*@[� h�ϊ���[���cՔH�B���m;���L���ߛ��a5LNH c��u
a+���4�N�1��4�H�jv<��,Uи!@
�/N{��4DR�# H�]E2bW���G�������ޒkZ��SeЃ"���K�g (zH�%R���~X`�N��&D6󭍤�d�\��D�IH��Z���hp􋪨z��F@wS����]��xߒ%�w��}DJ��M j�i��-l��Rw�=�l�ͫ�[O�/��[8f����&�0��pgz��2�.��I���E�����[� ���pn�~,��qy&������H�T'_�d�G��z=i?ȭ"���^q� ��}�9gY�*V6C���dzI9S�'Ď�m���w��5�A9Jv��-�hn+z���PBD�H|D�3�`��|��`�����}�m킔����Q��V����:�

T�٣Z
�%r�I�@���#�O�k��驭s?�,��n'�s�@%il��������]���	��6)ч&�wPP�v7<+�y���xޖd����#�*v�<㺳�-��j��n=��c�s(tuP�틃����A�7=��Mo����ڻTR�G��,���v�D�u����0�T�̐XN�.�@O��Iub�L]�����RO�0��G��6@z�n[��^�|���!be[��s}2WQ	��B��f�@���
��������vȑ�\�?��>р�,}��]cER��'i�O�b�n=>�>��͎ͱ�tga��V��x�l;�}��)'�s��|��P����O�a]�tŒ��>�ߤ��7o�#���V{@��-�G�C����E�~��G5�BE��Sl`���k��:T��\��?�/�y�Q�����#�@Q'լI�!2�D(aۈ�^)�r�����2?
��(��;�9@����Ywf�TH�����d�ُ��{m;�w����8�%axRO{/�K�eS���"�Ʋ�cb�Pr��d���J����PHW���������c��(7�;!SףT��%�׃�c	�Ƚ �F�z��M
b�8�y੪��?���=�FV'�'�y��Ǵ�U�ex�ݚҿC��X������_uܳ�:C����1�,�]U��'�Z�kFbE���ߟe���8#-{q�0�֭!�S��xZ<6��>X�|&C�/Fz�������~G5>�FN�b��� A��nʛ��N'0w������;��'���dj�Db� ���(s��"搽���2Ynʬ��K��p��5�I5Ȣ��C��G�}Q������v���j8����̖_��0N,�H�`O���m��)}X���a�\�G��Io>`x�Z�|�����fDGhz��P/�{g��3�E˖��φv����PLo�0���ځ���y}�؎x�~��z���4J��酈 �%]�7�tK�αr�H��旮�3���o�*������N�
a�A�>oh��InK!Ov�>�'�P����1��'Io�|@�lw	�
yqhK���N�K�&����\i��`-a�p���\P��n��i�9Kz^���=�}^�<�~�uE%��z�����ڐ����}�7��\�w����1�$��+ըk��9�@g�Wiˁ;z��mѳ�;�=tE���r�pѯ֦�;)L�MF��9���^�k�9�:P��� �?�����a𯺪8]?9���ۊ�)�l\�]��wftݲ���-��>J��[��� ?S�G�
���zq��YN��K@#��(�N
���K@f;�7��i�rzQ۷[���/a�:Ҡ���hF~^2�\�V�-�Z=�$��7�~��Pg$�Ya�~�����4ƸUnJ�%���c�r�)ʰɣ��k��i6��rĳ�#aĐr�G���[c�� �϶����S� ���ZJHh��C����q*Z��	�5It�P&�9�X/F>�8 	귖i�o$G��K���ˌ�{����2�Ľ �@>�i�	F}�-��?Ƭ�%��V?9���a,$v��-{�M�]�98�#�~tjP%����i���(֪�� ,���,�s��Eہ+����;
�}��9Q9v>�K�ػ�
�k��KjxG�jη���8whS��øѴ@��})��\�6n"DZ3��ũח���<�}���[�P�unM��Bq(g��i���O���h2�:��I��O8�95^@��ə��2�.>ò���2&;�]gQ�и�D� d��2����~n�l���K�e4�]�Π����sǅ�U��R,(|pX�E	��A+0�A���FJ�D���u��?�q�V����s�&�"�4A����.][i�����.g<s�#�p)��7/E����^���w�̗S� 
��A�#�]�M煽y�wZ�f�Uџ��F���RJf|�Ǆ�U�7��l�Y���V�`�w�4(c�xJ�-��n�M�/��!2[1���/��b���4���LF���q��y-pP����ުa�/���.�~�l^�֠6�3c� DN�?+aO��c�*��=������k��F@�8$���$dD��`����c�+ε�%3���x]�܉�u)�(���j��E	���uHw��Vy�ֹiؘ�swt�1�Y��*]����G�`��>*;���a)dY/>w.4�c�q
�}r��>)u�����ұv�×"E_��*�������n�|��j�u.�M�D�{�1�O������D%��LK��^ġƲ��:�@�A��q��8%۪�$2�$�gvm~���S"D#3=�Ʃ�Y^�&����V��6�u�y_���I�槂ftD9����O=)�[�j G@��=�|��)���G'�Ս5��+�鄬��P�!>�ٝ�������!W�q �z��X�L#��=�7�˜$	����p�O|e����c�h�!B^���MT�5��9�p'�H����K=�]�adbW������$�-1	�G�{��j���l�B��M��[�v#��o\y��>�ճP��ڐ`�;�켇�A*��W��)�f�9��8Zˉ��6���D�Dk�~S�N��c�)J��(2��B�n�����f'TtV�lѣ�ˀ�
u�ݡZ����N�I,K���%<��A�H�5=���Pw��X��4id��@W�3~�Yyus�E�kg��;84��S��^����!W璤h�Ir��rK �IbX��|	H�f��v�-r��!��;�e��7��q~'H�!��/!'�ڙ�Q+!o_�V��B�];ad�tzQ�D]����&��ŝn?�lO�c��V	,|p,��yt��@O���<~�L`��담Lr$it���M����A)�q��_������(��_��ٰ��Xs+���Qj'/���f?R�{���!��p��Z䥟�Y�=3#u��:��G�ڽ��R���(?�ws�N��(n=�R.��}�O�J�W�Z|_˵�w��]��8z�*M���+��O���e�0���3؃Ɔ@�D� R��fsr�Z`c�Cvb'E�痶}�t�t�����p
(��㇨�0TQ�U�bU�ǧ�]s��Lx&�WN�a�W��2C����A�V1�2U�B����]�}8��pi~<���Ʒ/����Q"������K �j��F��3��^�ħ���]�>�rP+}%�H`�(���QíP�B	O&|���o�S�.�J�NJ_<��?4�7_��M
7el2sԧ��E�9Qȡ���I Ӥ5�iM�}R�=����?��B�b��;�M@!�����
0��w ����
l � Ǔ�����E*�O�XR^<�0?��PsyV����W�nG(�Bp'��<���F��4vǿ��w'�w�`5㉐���=goP��y���N����W�nR+��7�t��V�r�O�(��Z��b��$��� ���.�u+���F�3��8ظ !��������%�/�Y��Qz�֒Fҫķ���[i����P��
��/�4���
�@��ڵ&�j*��j|�)�WōV��r$�����Ũ��Y7��x����K�z{���n�}t>I�#�v�ÈĤ����	��A_�p㱰`��x���[Qv�@����]��>>4�~[`1P�X��hKd����'�<v<���<Vm�@����s�nf)8��wm�\wo��=��U|j�e:!
k�,>`,�������`'��!XtV���NR�
Y�Ƚ�-j��g)�8]��/`�B3�F���Wg�����%0��m��l��ּW�#���(�����M�"n�E���!�2U�����o.�=-_�M����Ng�q����yh�m��˾Xc�����-�fB�Q!ЭMWbgٙL/��v��ay<J�!��T+�o���1i�`�^U���#?X��͊V'�=����X�5y�N\c�`�zp5�'��n�A�	4 ^���$H	ƮS�R�wtF)��dgj��A��B������':�A��� R��9P��7�`����������< }���j\̃tpB��#W]��CN28%r�&|��V����R*�p����j/ ���m�̳x����f�����F���;kQj��t���Zk�D,��=��|�z���q�U9�i��=�R�pW�e�����rKbؒ�t��%a���J����d�J����Y &b05�q{�{���(X�$(��i3��E�r����.����������d�����
�]��G�v�S���t�k��+t��rg��K7Q'\�կ�Í?�}Z�8Jʮ����W9c@���W�2ia��<��cLܤ�l���D ���%�,
����pB�Q�.�!��(�P�=�8ܟx�u�`ЌVQ��pb�ٍ?��P�w���8.v��g�QQos)�[�v	O�ܔ��D.%OѵR�m��,*�� ۽��y�l��
\�=:~��=93��E �=o�V�7���
XI\�mﻍ�uط�& �˴� �,�uދ���]�� \������f)������.�8z�/h�?U�HI_q[� w�E �ZBc�� �:ES�f��y�P�T|���P��.�)��y�Tkw#�^�%����?�y�!?�>`:[��2J�ia�jY�8��[;W�9����2��[����l����8!~���ڥ�
��hl��T��8�d�2r�QP����Q�2�>U��:��U	P���&<⎧�ifph⍑쇧�o�U3P�yV���BD�粄5�˝�D��kۮ �:���=v�ۇ��̰5��-(<�|:D�L��h�"� ��(��_s���+P�Ղ�j���<r�hף}�N����L�,��f ��}�������.%���!��#��;��1ѷ��.�87��$�I���KJKZ����3����>�4�u{dv�x�oe"�v"~�� ��zbk��v�߃���T��s������s��?����]Z7��]LH� �;RP'����Ym���k�E�T�&�B���ގ8_��e�L3��w��~޷z7�8_!j�#���z56�V�/f��F�A`��f��L:��s+�#nG�pE|��Pந�9�j2��%������vӿJ1P�����Id*��
�V4!���a�M��� ���2�:�+Qi�DEI��3�6ƹ{#���c��?�D��@�PM��m��H�0�a)�1�+5Y.�R��\3�����D}���tE�S|�e��5U82�u��n�Ϳ��M�π6�#����7�ش\~HZ:�=_���{���7�g�h�.��qt���7�9��N�Hڷ�r��T狙Q:m�dv7�����t���L����

�qt��iy�l�C�+���z�CW�A2>a�6c��47��2K�
F��Lڃ9���j�jWm�Y��t����3;By��wF--tYФS��K|ȟٟ���q�~<�d����눎0�u�L:���Ft�)�@4��=9�
�$���uN��tQ�}p��
s�������zկ�A+>Zf����{���)/��l�,�P�����J=�|�A�I
��e�v'��y �4���*�%*��W1T -�.�$��tE�,�k��kBi�i���R�Ūt3��bŗ1�8����,\))���v�(%�����U��e�BH�nt��g������~B,2���MH�	���Q��I�J�/u��5n.뵶�?m��USK�y�6W��_�����3�3�p��:tr���v�U|_)��\�߈�0Z���w���6	F�C�����O*W9X�D!ћҬIr?c0W�.�%:R��EސL��[VQ�� ���;-7M����A�~X}�a��0��X�F�>VN�#���	�ccu#"6b|��M�Z/SX��]"�T�a�3�:W�}��n���E��f��Y5�h�x���VB�3��
ͤ�Ν�"���Ȕ&9�F�-"�����+�EG�)}��{�i!�Y�l;��le�zr�<7�t���f�y���Ơ��]������Ǌ
�Bu������n걾s�;k��3�X�
������W��6U�,]E�b'�k�I�$�4#�Z�y�b3�+ؾ5U�+�F�!h�/I�u���?ѳ�vH�'�{�9L����c4�@����=_���>L���!��h�r��,� <e�Jo�3G�T� �!�?��^o���Qb����?�v�_�H��ۺiI���_{��8��G���5([X� 8S�G�fή?���|x�b�7�!�>7j{�oE�y��F����-I�Ӂ�Kb˜'�tAh=�wi�n��SL����=�]XC>���2�I��Ӭ5�}ʃ�v)z�Vz�gbۻ,��$K��\�2��!���A��\O��-�b�X�o(n0$喱G�$�N�/�[�j�⩫�7����D�}� ��	ڪF�`PlV��c��3�n&��h�K?��\]3ֆV�z�����lQspk� �͡�}lW��o�&)�١O��3pmd>��E���J.ex���1�cy�q�������F
px��Zz5��p�Cci���Ӛ��_0�e�����]�d�9+��n���ڂcY�����5�E�����V�"�	_Sehq"��Y�{�\*6���r�(UǺ�m�׫ ������	U8 ϒH+,旔FD,����z���a	�
\��aY�E�M=�J5U�'�Ѐ�9��ߔ;���E4��)�c�aR�L�����jB`'pf������z}@�(�@bSv莢�()o��.�r����@g�p��AQ������EuQ5��Nɼ������m����--��[��X�}�x���㏬�J�}�v|ϨTa��v�lEPX�/�+DJ�#����P��8�@��v"+:0T�<3���C���D�VA����+2����K�3�׀"�ۈ ��!�aE���f/l�N����`���H��9�1E�7DQD'gt�8�d�6� ID|�>"�b$��G(��{�����C�18���+{O�E�*nP��-5iI1��0i@�$M"Eyd'����?�׍�=�qd*ѫY��q�X��|�c�X��%������O��u�Z1��]OV7�5OO�zف�,7���a/*��:��M��K4�6��DË6�O��kA��"�wU͍,\�{b�~c��۹��W�3.�n.c&�^�t��id���)��:�Ϊ�{(�9A�.}�Ur+����3��h�>��$���8-�8� :�,�|� "8J�D��?�"C*hN3��n���dWd�ݶ}�nS��\	�����W�j<U�g	�����E�~D�ʽ��Y�����鮏��|+�����63!J]��nށ^{?��H�>�	u��eQ�9E$+�/9�,�O�!`iOQ���L��l_	�*3�k���j�&����[��^�]f����c΄���\;Qɑ�t�խ$���ĭ%��^Z�21l��YQ�#�,���	t��_Tⶌc�*��p� �|��ۿ�a%���q M�����+P��H<�:6}����<�־!��e@#9F:��}�9r��h8�\.�'d<:p�eB���>mn/�UD\�]��R����1�z���l��f��H���A���	���[�o��݂����Eyߓ d����1���i8��4�0��z+*,���fV+ujVy���*��ʔ=�Sb}���a1!���j.��]ĕ=�|#|w�`c	�=�8��J\4Mr���.�
�l��-}��ۗԨ��%��4���/�D�(~��7v�鴕����jU�Aa"��k�Y^J�䢐���xM-+�({y�!Fa7�q�� 'O���.)���^G�|��F%1ʥ�٭2@��[m����l�Ck�^�ۦ�I��"elm�Nd�2�2�Iav.
��#��R��j(��R�lP@��Z�t��t��vS'z)$�
��R��7��J@7�~�+k��
f0mF����,<)_�C+;4����g��y�Qu��T�����|�+�Ȥ� �_�FǌcH�X[J9��B�B�I�|������n�r
�9O,Ps�������`���p��kĐ��̱�������f5,�w݂�)�����S�\J��B���|0���R�d��3n�n"���ց��09�\��]]�u�J����ʈd�R���d�J�{"a�Yy��B��X���5�����#��}���G�A��Shk��tO;�c$���x�Mc�#|�J��g ݄�t����Ǻ��۷J�3٪�$ ~���o!ŏ�0e]pCO@��
:?s_�]���T<�.z��o֓t���j�N��/�u�����Y�u�c_��'7 ���R�vR�wP+� ��5<��;�<��)�V�$U�,U�i��P��a�N�M�w�f�r��i$���n�TjL�R���r1�/"��{k�٪�tC���HwlE����K'(�wV�Zj�=4Qx��F֥?����Sz���4�AX�މ]W���)�1�m�#�F�bN6��n{a�	]�׉��M�@�qL�o�'kS�B5O�N��Kw�Zs긊[�w��c�&�	_���$�56´˛l��Z�'�b��ң�1&M�	ϚC�����0���93����!�l�Z�s���N�xm�_fN5W+���'[W�PX�y�4�����vmԣ{�vOr��y��6���Ys�-�Ї�K�1L��ǳ��/���i[S�r�?��Vtg� 	 -��2�KW캯�n@�hsOjI$�u�|x�RAڱǬ��@9����D_Ð� �&n����q�W
��9�U�	.� ��d5٦(~1�T{λc
�%�)yy���WT�t���~W�f��b��AQ���v������[���@.��6��s4��SZ0�#~�2/*~RZߗ�e&���I*�w ��X�uFR�{���*�[aˡ�nq.E�%8jH�X�"@W���(���N=��4BS��/�=aS,w�����=\�0��i�bҮ<)����/"�������Do����8���L���N!h	�~:~��")�]��Y��/M�������HH��xc������^����K��Is��:K��.\�D����P˞ �_�;~��4��酪N�g��2��+�c��YK=��2�a����Z�f�l������-�� ;ٌ`-f5%�$������ϸ����?i����� ���O%g*!��Jh���ҕ�`V�z���ū� �&�_c7��@��y�e���j�+��M�C��'W�u�Nɾq�]-��ڋ0H��t�hHx!F��i��"%�[�8J1��1D�6�E6��kd�V�`+G3�5ޖpV'����'�4�a��$�;���鷓孿pF��qcs͉*cA(�V�b����"��)� ��5(O�r �ޜ�;��>��^Y=RrF9���\4�N����� r�`�uJC?ώ���������Z���}?5?����x��-�����2_��k�}���+8Lu�* ����o�G���M5+���C�	��MPŧ�h'c(�M.5M�����U#���i���T����������1�ݷ!0wHS�Bmq�mQ�@o]��G�.���& [cϗz� �Y�s�gB��	�d��Em�d�UR� �$V�U��_=$��"AL��쮇JjھT7ΐ`仸ߵ��W�[u т�<��4$5�b�R&�]z�U�A~q�x������<i��p�' D������}��V^'Z�\V�[�;� \���;J�[Z�^VN��2��$�x�Im�N2���]��E��6�|�KJt(��0����֩����&�*kV��_��P���,ױ��ZjM~�xt��V���Q9�Ki�u_Y�|�"�e,�L������&A�?V4�
G�B��x�SZLc��R4���ҧl�Dn+H�����E�zXKߺ�c���0K�BEG��d�8�F	�.�/V�L� ]��x�<�
H��u4}Ճ`�42T�L���˕�d�}D{&�>1c�OKTO�Fl�d�]m����M+��(�>K+��aPf�E���(�]���=UO�,� �-g���t�+O�u?hhR,�̅��xGy�=���
�0�պ@�����Y=�V&��x�|�E�J�R���a��zwGl�����'p����Ivb�L#��� 6�{�2('F�{p���w�qk���3��|�o�򠀡	8�1�O��>�����W�5���	������7��ϝ[:��6�[����3�fO<.2τn��]�z|�L��$��$�T���A�lƞwaL��1�TX�C�lf8���S�nW����P0�nF&�H�Lo�>t� W|X�k[��{D�Tw�ˬ&A4B�܇\dIѲ��,��o��_�
��wR�i\X���Ȃ�	�� ������ZK.V�^�9JX��}��k�U�a5KA�jrsi� ɂ�V��?��C[T�8 B�Fu!%HdlsO��[��`
E<����c�"o?�����	���K":QV���:���,�J|�I$��w�Š���}6!�n�[�P�i*��l��Y�'�e��s�����O�LF�H/<r��L�K,Ԫӓ����6�k��1w��9�
J�4��N�L�9'?[���H#��x��n�1�c	�p6sA�9��,��os����9�B���)�V�e��9�������H�ag�N�W���>�3M	��*>�bY-e��9̮,*ha�*���7r7��7oT��J�w���3��B���"�RO#If�:[�d�{b��6`.��$��8��˴��Ŋ�u]J���X�|ͳ"�]�:,��1|���$���y��j��Wih)�y�b���v	��%a��x^"�g҉	�� �+��0Tx�� Z�_�u�w/�%̀������x$F�T�s�h+�	�w��}�ح�$�: ���]����85xy��c.��L"��O����L]x�G'�X������'�����7~�}|�^�?��S9�z#�8_�p�ת3�=D霥��D ���Q�'C�'?���Ve	Ř	�h/UPa� MY����(x��?�^�&��뼖�����yA�84�V'jd}�0�}5�B��7e�~�O�i�1�@!�懶���@麽B≮{@�&_��wfC���F*�	R��{]{��uAR�ׄ��=N�SC9/v�����:�����T6�x��0L�Y�&�QeHs�p+���HS���v��!�Ȁ��=;��$U$mA��e@M��=�<�:(���Fi��|�I����fܴ�vy�Qc��V-�Mbv�M.�`Cv�֍9n�����B9�&�P]x}`h�k^��O�JP���U���]L@�#t����]u���0ʠq�/?�B�~5^�0UӜ⚵ki:���}�mU�����X��P� p)�t ������*���Z]��[u�ZgN��j�F��4��Vs3x<��E�2���0Da	6v⽷�>:��Y췵�T�xC�a������!w(m���L��ytd6��Н�݋���������v',��@ʈ��9>a���b0�?e
_FP�/HT�ݺ���b'ى����+�b��f��'�1��
�{ k���6/���b�Q �U��ˋ��bt�D��	fa��N��+h�u�T(��ӌ�bY*ټ~����唤��v��1c��rrs�|.XcGû�2�3�7Cp��%L�0:G������B�F9s�CW��+k�b�s��E��; 1杘�*��N��׹�:M�h��ocO�&�$ b� ���I��́����5�ۺa��H�H�qf�.Я�ҫhG*�O6?��xF��$�h�j����˙"����S�������|G�O�h~5n��M���>�Y�NgN����{Qҟ�u�xܣT��;�������S�r9֦�Pp�����חZS��U2(?͍�ڤxwj���0��G[�	ҙ�);͙P8��y_\��S�FJ����� r�F��[� ��@�#T7���3X�j�cް@�����Q�)�ת�0r��hl)��HK�f��l��y.vw�&;������JNk�-���=/e7K=U_�t��l���ܫk!?�%���Sz&��}C���0�4΂ z�L�e�28��
%&#�����Κ\'��_�P���Ex��<��Q0tn�%C�������gĵ��9w굃$#���y� -u�m�GA��'�F�0���M��\�^Dc�'�T*�/��v-��#��K3>ۜ|�F4e�S��9푬����}?�BHf����	M�|
n�i^>᎑����>�Jw9�6�Y)G�ю�Xi�&�?����"}�]�F�����#��e��٢0�T٦�c��?~���j�U�3z)���c\����褫�k�K�j�6o5r(��H��'�YIe۫��D-]5Ү��"�3ޱ��|�$����9�~O����p����q�;���<9՛i�r��e���)^@7E�O$�&���c����߉�@a���)jܝV�u�B��[-+��i�\��Fԡ�x��,�4}L�?�_\aY��k@,���G}����.L��\iC��8��wj���&�_�
�I�C�A�ĺ�l����%�K~*�R�=���cR�<-{�!!�_�ܾ?���d����j�Y�.��v��<;A@�2c ���rޝyPO\�s[�Lr�`g>�Mʹ<�(�o�-'&����Fd�;}����`�A�7�R,������C��1M�y"k7��d�����{�o�R`@m|��mh�T�'��ռ^��	U��i�c�=( ��fpSfp�
�V��Xbt�0*M����9�c��׭�/�
"'\gl}���g��<$�q;�HL�1�� Ѧ�1�!r(�����E��R���P����Vp�������$i�R.Q��d��\u��6�0T��3v�oXc�J
��s�
2MiE��<j����7]Q�"NM���P���`��SEU�1��B,�S���}������p����אe�d7�ꝉ������m#餩R��|����0$0rj��
�C;��z�3nXc��0�Q�l��Ĝ�έ'i^:[P7o:x/��C}����Ӻ��+��F-�Ek�k^[�\���E�1��� ��]���Cw*�<�@G)���A��Ko13w��k����w��u�J�����֭���UDh6����eϏ�k��:%�pH�s�����W��'��
t�i��lY6St��S:~���B��C�+f��{K̉��K���#�h��� sBg>�́�:}TG�YD�a�T��b�p5O�l0�W6A���l�w�>�b�HV:�F� Ph��|'���\%��u�v�7�`�v�����J\�E��^;����O� v�W>r<��`�νe�4w)/��OS���Q�o�x�}�']�#��y��uG�t a�82>ゾ��� N�����N���GC����Vg��/�z>�.V.�5���D��R{�S,�uw�h嗤�N*�����0mKP/��W%oO0���ji�6(��w$]&�My�u�D��{`x��yiTř��[F� �6�\������ɼ�Fg�^>�>���#WC�y�� �e��o�}Gc �=�c�!�~��Ӫ�9��&q��#�t2��ND�+=��A�UF'�� �8�,��r_�E[#��ش4�{�h�En��Qe��3{~f��c�� S��|������6��(m��^2�t^�Ƽ+�l�,~H��w��H�h�o����>��pW|�G=+1��@m_¥U���qkC4 ��? �I��m��E[�zW��>�9ZQ��G bU�������'��'	@��Y���Q��Km��!N�w����?�u����*�+��_��|yڕS�0;��#QI��9ғ�a:����Wv��[`�2�tI9i|Xl�$
����:x|/����,����S��/�o~��H�[�1�Ev6ˮ٦��#�%)�d���tG�d��˛�8���[D����IX�O�U;�'���Ņ�2'�p�
���/�'h/x�KL=z^3�
f�Ir��N��*xY�u6?���쉕9{��/�������7=�(ڵ#9��O Nɀ��m�6Z���~q���_8��nt���m�����������9K��)�'�zf೼���2C��Hْ��(����]���Nf>�P[�I�W�������N��چV/kX���6{ʔH�����܊�=vٔqRA�X�в����2Y�ZJ��ZF�ե(�<aФ� �L!��w�^�1��tJD�0N,|��V��p���S�'҂އ�QH�)��ka���4b�E�x��l�&DH���\�M����q�����z,���@`;�Dl�ջ�6�^�2��!�a&A6T�iӒ����Y
8���9	�`��ֻ�5-�������L�н{�l�*z3����i�~��qޭT�G>�A����[��촫W�0,0%��UҦ�A>�����r���*Cx�� �O(%T��o��Bg1X�NӪ��Qr�|���h$��L��N���5WՐ �(>'�CIK�Ƕ�Y����S�%�:�q�q�5��#OO����7&�ޗ$b��U �K$����ΪNO!�ܒ'Ň�I1n���e s?�P������P�R�Y�"��������_S�]6XdV�e6��*ڻ}���v���A�Jkr����7�)���YG-��Y�q }?n/aY��EcVy�[il�`!�H�u�3++�ϙ�*,�~V�)�R�Sr�Թ'Y������E��2ܢMՠ�Ϡ�x|�d���\KN����Z,$ӎd�:�H�<	J �Q�	�1$'�\�<M��J�ʭ9%��u���G��������PL��(ea��w�O�n�i�ӯU[�]�FE������ʕ�$kr�@�@�Jr�#�I~%���œt�'��UWw�eܤ�)#���_׀����^'��_�=�ʉR$k�x��7�0�9�]fB�hyH�&^�;Wv�-�i�yC�@+k7p㿖��_S2�Or߆df7kZ|;[��?���m�ޏ馧ۓj6��t����a"�U�Wq����:@g�%�G�Q1�&S��e���\yNj갺�^]4����h}��QDv2�-o.���V]�d&��ZBV��L�8���N7���;�X�;�[�+�g�� �G��Q�� ȇ�Ek?Pϔ�Ls��`��n�W�Af���A�L�e��7� �����A���F]F�]vKq�H �����)��^̻��dy��Z��C��)�|�B��TV0�a��;�ه�{�'�07�$�<��gr@2kE4�*8fU��q2�^�8�B?m*7�����It:�ZG��h>�t�(Y�������Xc^M�TaV��$%��wux��z�$s7�A�bs�I��4&���}�uH.|0�NY�'F��8���(cz�%MN��Tg��ţ���Q���f�%�_\�U�~����^��ܽ3����[�טs�<�Q ���o�|�M��%�"��e�B5�5�/Sظ�sb�[־0�EP�'8��I[�cO/Ϛ�_u�ݙ�0ǜ�M�6���x�Pm�m�hZH�9��Dh�(-HX���� �K��|&�ޝ�Q`2�K:	�dI����o����>C�'��3mϳ�mW�U�-�P���ެQ�T�fo��	8Z๼'Ѩ��ʠ�S�^��%��`upo�9�b�qs8s��N�vڤ�b�dv�Ƃ�"����C[cU��=��e�+��lQ�ϴ��žxg��	f��{�Q!�Wu�>�G�ؐ"���2�$��c{�NW�:�J\lt��:�Rƌ�W_��5!����t}��vʁ�Fү�<�uٹC	�aSS��4��6�5�'W򘭬f����wA��vr�Si�2=j�]I]賟�')I�M��?���8����^�JyDG�.�Q4����
؛	e�(��2������tj[��W(^<kR�>�8���Kd�]r1Q��������\�~�P;>uo{�{*��\��P�T����@�y( �qr�QUǊ'�}��3�-R��yx%-�Q���"
Ӧj����ˇ�A�	j�mW������UZ�1޵��v�4����<���Ɣ$��M*d�����q-�)q�Bs�A��I�D\Pi��$p�yZѦ�8�PZX��{��PW��=]���p�f�X:>��C�fA�d�B�/"��,v�Z�.NU���#D�v��x�X8������Pmh��o�\X�� ��d@�B,b�x�+�2*�;�j_�m�Cw9F3���T����ï|3�ck��H��0��������H�*��"��9�ղVຽ��5B���rUڇ����r�,V]�TaHY[�s�9�-�o8j��y�d��.�����+�S��tN#Ae���h��C�I02P�v��{k�^X���ƾ6�6���v�y���5���ڰݯ�z��~�����|řMݻ�s��-�Pw6WD2]d�vomY���}l��
Ml�d�,���E�W�`M0k�qm���3��>al�dk|���gx�+��Z�>/0�b�����d����yi�����[(X�=��V$��3kJ�h�==ϧ�����$Z�<��*�j[���2���l@aλ\ܓ Ql��#�A*N�+�|ZUk�'�O��Hn��n��ti]/ �b�HY��!9k[F�����Z,�^��z���R�
�h�J�+�� 8�t���MQ^�ʯ�^ܹI�cP�����c6���草y�MM8���������I���Z���˘Q�˪�U-}P��\��d��f)׵��]o�- ;Y�_ㄧ��a-������FA
Y|�o�����jd��V	��HN����lM�/��z�+Zk��S�F���掉�
��ld4Y��>s�����qA�+�m�i1�`��N�
�Y�f���oE���̅pg����;{x���A˲)b���3Qp��ν�K�!�k�u�����~�u�H��r�JN��H>͢ǊV<l3����t�HRU�e96x�T�Vށ���R�jk� ���n�(`�UJ��dɟ.kO��$��s֐�V�=/��L��'����9�Bt�K�Oq� Ie}ֵ��E�DK��&o�7"�R���5M�8�d����@�!cC&�b ��6Y�I o\���o �7�v�-|wZ�BvQd���S��|�i%=���@eq�i��#�5c�c�h�;��G�T�YR�2������\�"�}�}@,��_�*?�>�᝚6h����Ok����I#����,�[������ ���:�am�^�����xl���߄�\���Fŧ��Su
yW��"��՞���S	99���@ֲ����,����@�?8�>��L`8������_���<o��_H�[阨�~i�`N��x�2���i��q���H���\J��'���!)�-��5i�.<���P����P��:���6_�}�AfxU��7R�ޑ��W0�vD�=' ���5Kbv��󥃸�@ 
�!��dG�Q˧���ґ|r5� L�C �����3��a�Vuq��	=�4I�F��#���@a�,�ݣ�n}������AD/Z ���>��qSbM/�k�L35�{��F��0�H�=@�Ѡ����L�ب�PW���8�p��2����-����aC唈�ܭ4�V����)z�����X��4'MN�xRU�_�]���}��PNNt��_%��5b�;��h��>�1��6�I�<��X ���I��*�1�K��G�绬�zK6�������<�u32��_�);�R���<��%hf�����FE�G��U�'G�%b����k&�G"v�d�A��@XP	�6��Y�>&�ٳr�T/���+�x0,�S����웆	.>�eyCֱB�;�Cn��Gy�p5�������W������������B~��;��_P��g�J�xާ�c룴)��H�x�zת�8a�`Ȃ1��*:���:(���N.��@����d+֒G+��R�M͑�Og�[@��	$# ��?��D����BX�忠K��b8�X�.�x�~��V��V�v����d���R�0W;L�9h�q�e')�KT"����-�'=�@�5����[��4��M���Wg_Q`�b`2��S50=��VT���@Uds� Y���:_���J��Lx|���XQr���#!
�dE�O��&�c�jr5����T}$W~�9�j�c�M�s�i�@2���� 2�ЁʁGB'��ŷ�h�n�s����;L��� �)R.kƕg�X�g�������{H�Q�C��M�+Wԥ����2���kH:���8$�y*��s�#04�m�@����o�?I�ҵ��R���:��q�{E�� �#��YkQ�ôC��34�Ѿ�g��k��Zz�}�Y>cq����`��v�t�T,,n��%���2�y7��@�r� ��N�4w�I��Zķ�U�̱�&��"��v���4��^H�5{���2�sAs�i�x��U:�tIvY�rME�ݝ2C�%��b����n˧Y�_��M��e�r	z��t0^g��q��P��$��d#��$Gmp�X�.�,㒒>s ���7�ȓ(��ʓS?K' I�-Ñ�Y8�%���`ܗ�w3G����;��C!V��q��* �u�?	�v���::�����������,a��S��C�ZD㎖�o9I������b0��{��h�����w2'���O
�o�;�*����S��qI��E�#3W��jĺ��ٯ$�����J�`b����#�4E@f)q��$ݛ$l�p� "x{��}G�6��e�	mKi�<�=^[&(�ӥ	��pqZX��boԙ6ݔ���Y0��z}�a|�!��Z�^������oq���56U�^�KAc,xe͘���j	�PC�2����5�z������R:�FF`܍r��Q��e0�l7S`�����n��%��j��/<���Y����F���#k,�D)D��o��d.=ּ�]��#��?U)"տ��!y���vhAfg�!�?y�Y���ڿ�!h߼ޮPA0I#�JsXՅ���)��Kqjj����n�Ĺ�w��b�0�$fz�'�&��%~�M���o(R� ��J��
�^T������{eu	�
��b��pl�e�@����X�^��I{�I�>u�Q9k�������fͮ�Oﺼ�M`a$��o�3�jNp>���b?�h'�Z�َ�q���@�3��X�7?x�)0`;�R�K4\�w�v>�C���N׆ߚ6��?TyIpa��z2��v�T[e;���漾���1�@��e�ʰNܵ���9z��W_^��ڙ�s�Z}��6�4��H!eA>�P�)���9�p��N�qe^�k�ԒDp�p�˕����c��U�O�ی?k�����k�i
Bz/`���N�3��8�s���hN���= $'[����+������"�����/n��)����1��jݶ;}D�rVu5;�Z]n�m~����cRP�����|��P��V
m�Wu*)�*��}�o"��v?^2w��=�Z|;�]��A���	��oֹah���jArtKl;�9����b��~����Vn�	�~-p��1S&��?��5��n�'2`hp�a"��k'�&)�4�SJ2R��e��e�L��s|�4�{1��k��O��F��w�>9�W=���aP���T�ʖ#��m��[�{�v�Ξ*CA7R���yG���u�E}�Va��9i���\�����:��[_�2.���5ɜk��h��J k��mϑ*������kI���jͦ���{]��{�i�&����2�?X�q��7��+&�Щ꺩�i�"u�
�g�pt}-{KE}�WЇɳH+�c�����J�x���Ek�9#��X��Y�렾4���*������
w�I�9At*�6���$���拱���Wt�W�s�U0���E�g��dZz�K����!�(E�Wj�&<����ZB�bxHB^����.H���aQ�ʿ�����m�� ��!~��Ï���#��h�s K�g�?���*��GvScyV��ߦ��i1����%���'���Y�����s~��3��\�;&�Y�ʦ���uͦ{xr�vO�;��U ��]o����Gǆ��=�d&��LuP* 7��"$��k{=H�!�m��d}fY�"Y�7H��}��xhT,��@y9�L��� ����P���=�js�R���Ƶ�yA����u�>�S���Eb�������.G�� T~�yK��S$�U]�N} ������Ӓ/((�$�iS���O1ag��"Z�R)<��6,[�᭯.��:
l3��2w�����)a&� �8G��<9���[$�i\��a)2��Ab}%�x"tX{���zW���|�O�'�;����t�I4&v��Z?k)�$F���lj���G�<j���rFw�C��'B�m��}0�J���/_P�Q#Z;���ӳ��1m$�ëBeL���L�������G]8�91x�y� �n�	f`"�`���rɞ�c8(��O4"���W�ި 1�QrR�h�����?:uoV=!���Gc�����Xޒe����/�ݢ�T>��ekp��a%���t���|0V-d1F	U��V�f�b}�4ν�,���<ζ�cn�|o}j�Jk� �Gg�	'��=ٸL�@I�.��ċB�cm3�})\R3C���s<-�
?RG��mb��E��+ZI�Y7a7k��}q:'�.!�^�"⾦ �%g�Μz�j˕���d�D�X�~NBq�'`�9��8��[�G��g�)����!��:���{)�5G�O�@5����VUlmdYN)0p��:%���M^һC��5Qu�E:!��ȿ����&f�0���&O#%��!�h��P�l�W����vh]��sP�ޅ~��f�Lu��R�/Be%ʃ`3�６����0�q���h�,�7/$<��B�~��h�.���kfہ�a���`�߇�c��.Oɫ��������5��*���DI�1�1�;����&�;"�пh�3	4�9nI6�jE����Ak�j�1n{���ÐYec&����7;o2�a������1��W��<J��qn���k�F�J+$:kb�{)۞�����tA���*#Z�5�&~-�;$�)��r�fj�z}���aM�i���Y�\�����&���#�Է�W�R���Q&H�F�6��˔���3	���m��8VC��&9�f����2�e�6O��L��G��~����yi�n�x�^hr!���&���>CB��BL�]�9ۅ�1�c�!�"\n�ǈ#�l�	 6(޽?I������B�z�R)��J��JSHS<�W~r~�ZUB��2q�y�fR!�V�kK���+�x��wM ���}�p��O��@�`6�ȷ\�Js#3���0Z�� ��j����uJ:{���o2#���o>�}AY�s콮���qv�m�S���)H�;����[�{j,�u���n�}�-l�d���|��~b���[��dKM�7��=�<�$^�Rh�0�C�DN�S�!^W)j=� 1E��]3��� {KEވ���74�;]���<~H!������5t:�+�D
��`����n��:ԭ<��&	9τ�r�N�:ݨV�n,�Ɔ��g>�M�ۡ�B+gRױA�4q9瓈q�7�{�x#��&&u-Dr|4��|.GL���Te�;N"��7InR�/��=�x,�1�qhY�̠�	;��
���!��e�k���g���������ca\@�۔�FI�W���2�)�*x=~h]�8u��f=�)�������n�mp�%�3��GA(\j���-nN0Y��G��4}x>��}��G�;ư%I��Y[F�r��쟴Z)�83��^˺��iRzŲ�܀�#�� v��)L���9�N�E�;�A���7@�����0]�%u����D��M�ȟ(f��^����(b�����ai0�c�pZ��FnN3��8F���p�'�Q:�W����
�>���ٖk��=��"_�3��x[����訟l��R�t��gt��cZ0�,�`��P�0���ElOd�3(ᢵaO�H3�5j<��L�e�be�D��H�ߍN$��"����R����o�˲K��N����^P��V�Hdn*4�b��#^�o�y�+�PXEO�*�=�9���~����I�f8�jֺ�{P��/���Z���ڞ��'��M����Er����(��tɅ�?�]��(p���R���a���U���;d	�-,6!^V�!��U�@��[����Q�)U�r�����w�Z��'����r1�}z��>���5�����G�e��P��F>�T+�h�`��/�@���
��dR�?$�U��a_�M3�%`�D�k���I/�0O�
���#�u��[0i�jV�h��#^�9jiNC�|��ɜ�	���;