��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����{hi��7	G�����|��4/���YEs��Q��H�9e���ϒ��(��t�.�?�ѩ<�Փ�<�Evj���T�����B�ݰ7� ػ�3��p�����D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�D�c�;��ЄUO���?�G�����d����w��ܳ�5�@��=T�σCFV���C	��r���o��[��C)r�|Ϸ�A�4���b�� 8v$(������c6���:�[�IL�&�זaj�~����[|��|�/�xڑ �#��t��\�88���jG$��N8�t����#W0�����U̓ZJ�d�E��gr {��
�+9�V��Fa�\��a�7t�=gF�>����Z�峺|��-.:�KEV'Ѕ%�d��ᣠ���ڊ_V%��HO��c� :躪���8>_���F��u�U�9waM�NFk�"ϑ�iĻ�C؞�s6mrGh?�&��ߝ;���3����G���o,)�?w�#���t
r�s�R�v���|��r��ޜ�pc��0��������J����@g�������g��ܧ6��#��{�:������%�8-����f�+t��x�ט�1IZ��H�Np��X�G����Z�l�Hƚ�Lʇ]��>��]:�W�{{�xuYɶ�(�D�w;ӈ(6�Cp�Y6L7:�s b�u�C%C+��t�M�����eܨV�&�bi�M�t���&��sFaX�`@�VɅ���(ik�wp���pJtJ,�ל�oɧ���OB�g�/�hȌ�Ut	w8�d�sn�<h_�+j�{��S��tq���)M�r����s�p��go-���H��0��R ��"0H?����֛fb���N�>	����@������+�~��}EC&dt ����B�$s?,`A0vI`��w�J���(6|6�tث%��tkl�}4�;���a#=�UJ�+��M�.q���8)y�F���f<���q��.�>�m���}��+��.��XB���8�����]�?r��ð���S��i��{ʒs�V�3}�&����%��<�{W�ǟ|�2��J=��-� 	�_y���*����<�qF��v=��"��1�n������`��Ȥ�HM�������0&Y{�-�����(��e�<˚������' ��eTav6�7�IÛ� -8W1͈�
|�&�z����/������i
}T.�� �N(�?� ������z�� ��K�$�!�p8�w�e�$��E��A�Ȓa�c&���!��U�>m�-(�1�Q�&xj!��B�xR'��ks�o��
��R}�q
�2^��yB��-&pP����
��*qO��D�v�>9�?��~��i������f����?`^*i����]�P��wF�ڪ5�c�l#�� 2��+mp�8��|]�:�I�GZ�k�DZ���U�B�)3���K�������Fl�v^ /�{� VM���vb����k�݉ñ�#_�Г��L�vi��V�o�3/�Gw~�Z&�f�a�����m���4.�u�cd#�m��vZ�g2��L�qm���� �0\B RIä�M�VT��C 8v�m�,����(�P1�$}��!#�j��V[�0"��Ճ��B"��J�E��ٛi�1�s���������զ�� �U|����"�-]��iH��1_�8�)�9�|EW4�g���1��bl�{�/g3��ϢR��ֹu�x��9 L��x{ד�sq�&nL�y��;���#�����w�]GwC���I͹V]ӏ;Z}�!��b���CE� �Cynq�B��C��<�,��M��c��;q��M�ä�U�:�jy���(����*\�Y���;�PEh��(8�h���0�P�v��M�R�"A��e-*�6�c�#aE��<�!>L�F��B�+F�X�����z���s�aZ�y��dj�s�{S�Q4��Buo���4�n8��H�Y;��3�o�8��u����  ��thEe���vH*Ƿ`�2�F�Aͳz�RYp�њw��o�� �N:�)���{P3�ÓIv����+�oȕ���`�%�nG�a
�f{����|�1D��V�W�Um��R���u��7m2z�~�EA7�Vk�~�͚�i�zg;�M'�����6p�qF�=*7&���&L33�؈[yXd���:�W�QY}}�g$ F|�L"�J͇�j5U�� ����/���N�K��7P����K�I�'EUPk�Ut��Q�������&�[��x���
-]��,I��Ar����j=2AW3CneQ��������2��+ �Cٜ۔J��_[��xu��G6���,UvqB��%����_?�Y���Y�hE�Z,Z��E�����1�C����]���?ߡ�B��H섴  ���JL��ho�G�nr]4q���Aԧ^Shσt}��Z���E�+���h�ġ�����I(1�l֖��!r��JWƒ�-���m���u�O_��2�I��=v_��=[��M�iS�[d@w}*��`�vu䅉�XX7�	Z��97�݅r�;S�ݻ�ƀ�Bc���-�� ���|���f���u�ne�D�
B̭��)�hӎM9��]��H1��q�l��������#�{t��S��3�߄c�&YA�G��\i�p$�2x���t��F8�T��Qm�HV��y5v���?�mU���ߪH�E�m�}?@aMm�yx����x�CoQ�&ISP�����z.�t�n4&���6b~��@���"�#��
�40�����80��:�1e��p�x�ЮzK���b�1uq�{
�-��T)NC���c������_s���cՆf���ih%g\����J���P3±=��*��i^H?����.���tB�QB����W%a���|�qx[s�h�rċh��C{P�g���2������@n�8�}�N4~ے�����ۿQwJ2Z�|bX��1��3Zr6.4���^}ՑUr�-���C(�Ҵ��,~�&�ɷ6�|�=V`Bx
�?[�鹇R�$:#(9No��:HN�gLcc���m�!���֧�m�԰�~`�Yuw��I {�핌J�éz~�(���IP����y��ɽu�BO����/��������א|���ͧ�8�<��鄝t :��4���T(���N��ay�.�[U�B�x\�)���*9��і霰�Kj�:2b�e��]	����pn�䛽=�v#�5�D��4��i�����GDV�-C߳���@Г ��ԓGa��1pK/4��1���)><6H��W��U�f��1�u�`�ǎ�����Y f[�ն�(%���?ß��+^�z,�_6�k�&��4��0T��C�� �w�cix8h�r�e��a�3�$z�GDj���U*�$�����y�
��7����ax�=Q������	A#y���+��Av8/}�B���y%����3�u�?���X��}Y��!��S�	��D�`D�~2��ߝ�,�J
�W�K�C�.t��y��p�����K$�iߙ�k�&���|IƗ�
A#�i8�� ��8�ல#�5{D�B���H���C���'�>���n�ZI�Z�%��h+X#�,�����K~E9�S�Uj<�3<O����O�e�h�u@!m1􅨙+��9����f�T��5؞�W�������o|"Y�ݔ�_��3�b��%
/Y/��k�p�=���캄<����m �X9q"�B�ǤL'ޭ\M]��)��3��|�<]�r���ǆm�M�6�>�[9*��U�;����`�s�!L���ws�l,7�њ�m1K��n{U���Q�(�\9���VI��,zEU�S����u�y���Iy2��'�>^0���	�}�A�Z�wߓ��{n�9����W$��6w�g��K��'��X��W��:��I��짙sݳ���!�jH�]�QYwT�]e_��8�4J��;d�oӭ_��hR?�p{Z#����(ВZb�|��S�̤aM6�9 ��dn*`E���V@l�;R5W0/�& �0��IhJ�{����="%0R���*M:���WI�����9-���;�L~�'C����:2ZP?�/�܄�%���iGd����#J
�����������U�Ӑ�R�^6�����
�Q+QoJ�R�4�am�LpM����fŔ�L�!��}�:��A�N�!>Z,�=�\�t�T��@,�"�άS�����*ax I	j^G�r�(�����Tr��l�Vho^�I����V��d)+Ӆ�ߠJ �~q!<�v;)�+�5^]�t}��h3S�\�2�����BE�吨��- �O��s?te�U�C��x�7,�hŸ���t}ؗ��8���}xs����z�U񙞱h�!�>?o��~� �����J�U{���d���3�q����ӆ�B�M�m�a{�rpg�=�	U�E��/��4*��;���/!�@�
�]ϥCz����%���Uz*�����r�&��(�=�V�q�)�XH-ZL��Sro<������JZjo�@�S,�$���dbߥ�(���3���L��;9#[ֽ#�~�ϣl�R�>�=l�:����͘,�xIܙ�&K�I�K�d�?Fo`�M�4`[�G]6��<�B
@L�nY�`�1oFء��y���B*5��-Ԇ~Nr���t���\�J��3��� 엡�z�Z$g� /۠�,�D���i��f}�Q�e�Eθ�?��;���,���`B��Q�f���(��r�ꐇ��Q��eW��'�a���rˢ����_��j��v�S��s:���lG� .<��rZMqP94�1��2�ߡqP�N�������"�%����B�3)%��6d�s����EĈF�N��i�d�*<;�Y0�^�������e޹�0���u,�+�:=��t���<��"M���cH:M���v;ʨ1�4�̾����)��u�����<*\��s\�<t7;�_�Q]M���< Ʒinwc<w�԰OΠ�ʁ���,��H�9*������߳56���ԁ��3���^��WGZкt)�!�O���u�ڟ�*���UW]��}c�W���M�\�����X����ʔΏc�KG�hRK�qR�Er&��֠el������������!X��`��y+ԨT?{g.˶;�$��"y��ԋ@��H��s����_d%-�'��4�/ꉕQ��!��U�e���W�^'ضɶݜ	�����N����{���B< �����L*YGVQ��tf�ip(!�h�e\�d�!HI��[/�t�榸狒 3Xc]#�P�i캲V�V	����k"�p	"�u��8)��I�iʦDI�aC8���(�<��dth�d#~��R��o8�����kM�zb/!���������&�/D��*�(2D7�(
X�����_�PJ��ik��c�&*�!��1�E�����	�P�6��P1�����z�uw���n3��{��nS���r4��!R�,������F�u@��l��p0�X�v�YՕ����f���J�w����Sɗ`&=��m2��vbN  ��K/Ag�/z5Tv�w��' ӡ�)�����s��0��Q�K�=�!?7_���(J_��J�}�M�EjS|�?�=��,.���z(򟩷	���ğ���[{;�2�FckV`��mI'�	G�O)n�r�0\�������u�8�<��b�*�CMǎ�0��8�~�`ѡ�]�7Mb�r�}�Ċ�*�`�9�������Ĺ�����I�$��ҽ���\�ݼG����cG�������-[qW �wN�ȉ;���-ޕ�Cy�����~�]���N����ec�X��%���HG�	�$�=4mI�L�g���ϩ��DbF�(�	w�X�-\t��)�����8?�&�Sۖ>�q�S,<�j��'o��)Q�*��շX��� s��������1(��cbeޚo}�C
�K᯦��]��ŃܟW��A��h^�M��CN2�]��m{�&��)�^Y	s�g&�V�·�6�G�e���y�C�g�!BLLX&̀zB�ٌaCZ�E�����'}oi.Jr���qM�,  ���j�
�mRW�l�$�5���6�y�p~��BN.�z����`=%�3�>�����/w厙~VkJmD�@�;����6��,�w=���\�=��?�/J��LDI4��&��t��cj��2�=ݓ�'/��DT��M��iKx�B��A���2��XI��R��s9��;%���F�j��`�ؤ����"�il�]fO��f�]�"��4Aɷ����Y�mrt[�1.���ɹ���`;.?7T�LA�Ta t�k� 5��B��`�='��N/�75���L|2��O|ߡ��1,�`��>�H�>�v���!�?e`C�̯9�s�[/�T�)�`�^�K��T�*9g*�����l(Òy�c��w�%֌��p"i���ӷ2G@���:��o�X����g\�k��4�ˏ�Z�-_i�?ґ��h�0��}�L|a����`��|F���@�i`�� ���]�B�8���#��2o��zb��N��:�h�-�~e�$ |��b^��ZAw���xWD%x_��mb� �si�-0�'�t�%�qY&���";SRd|���x������]1�0��GёT�.�%1��i?_��&t�SzH`�������Z�3j�[�:?w䄯���]��v��s���X�7��X��/��3dCQr������9S�Q3ұ�,���-�qq�c�*�'�A�l�'�vD��}���2��1�"U����$�1``]�="-�� �EZW��N2�#f��c�`���
�u�]�%-YN�W��pd�v�����D�m��n�lwy�!�Tf0�7���t�c�l����@)W�I�D'a�φ��k��G��s������E/|5�F�>�z�p��X��~�0���񱞌y}�4x�"q��ixČoQ�_�&��4k�AZ�m����-v�%vÈ�0H��K�|°����o���!{��1�蓿ڋ�b���ou��S�e���i#љG'�|iJwb�F"-	f�F�W�H]Ԏt�-���=��]j�1k�B.�V�h" �v�,�Ucq^r�:�����~�A��~����~��W����W[�g��B�r"�{g����gQ?�����(,��ܡ�b�E�̉������`�n�m'�����Z'i�n8���w=<ٍ,�мw6�N��v(������l��X)=���V��%g��L�`K�e��eF��j��#Q��TB�};�9����Yo~�P�s��|	��Mg�T���L*�XԗF�Z�^�Ez���%m�Pږ�8
�'�U`��=�{ݲ�X��@N��J��dU#��P��/�^W�f�(C�`o�Gdz�9N�w%��$D=�t�ϔ��9-餜�W7Q��̨q����$Ǩ%�����1g��[�0\�G~yC�zhDD�k��8� Jڷ���]�Y���m�R��!j���'*��Q��TMT2�ћ��hC��m�QQ����J�����&`��7#P{WÐ����ʶ�y��|A&z2�
$$&>D!�̞���cZ�[@C��t,�8K��ÅW���P�6�]`���VJ��L=�2�WZ�Xq��ᵝ�M��C�7�2�g)�]��	n����c�+�[�IJ����uՁ�I��~K��_͒�H�)�!�$�����F��.M��ZdX���G�[;�G^qԍ�p �v��c��}¥��<u�M��P1N�͡nщ���dpf�oUV�J�,w���^n����/Ԣ��R�,�7|�/x,&ʚ႓odz�G����^��݆�p��	>����H��*S�4�����@�&b��X	�D���^�?A� t]�,���M�s�$���r/�TR�s�����}�����*#v��E6#���޷)��kO���b�p��:�7<o�Z2����|^�!�h�)HxE�)��@�v���9�Ǔ��vu��t(9L�ƄR�ͨ�0�aR�����Gy��������/����eEJ��)ן��������	�HA�!��!��S������|&0��j��S�
"F�'����j9(�4)f)�w��YQ����ܟ��2�\$~j���,�Io��K��j,�]��є�B@�4?�� ��[� C"E�@�4���4�%���M��R�������� x�b�SkL��S���W����C�8�@͢�������xt���k��B(��_\���MY9YY�xgZ�iQ�ꔌ�����$x̚ B���7)��$#	��	�6�%h�5�4�0�]dh�?	eባ���LlF��01���$b�EY �t4\�SЖkPx�Z�o��(��v<��CZmG��g����Q���:~ w��̔,���e-�L�@�6П����~��Ҙ#A�:��X΢�������Xq�i[;֮��8��x�m����ɛ��Z��8��Tl"&es�=jCz�����#R�!�/��\
�k��>��C��"
��K��\+��b�7�I�G��Z�6�\l���Ѧ��&J���ܦ����̻5���	����i��=��h�){�nhE�I��u�V����7Yɧ���R�-rC��X�(�b8ە�a�6�����@\3���5��E� �<�)�/���cV���'����?X|;hn���$�]=#ۂ�<.Vf�S-�P�;U��ʿ��׈K,�~�������	n��XVRs����/=�Z�f��!��`:$��n�h��y����B�l��i��N.�{ע��W![\�|.|ƫ���Er�d�.H�~��?P
5��IK��P�7�UO�>��;��4PJ�L���V�k�j2as!��_c*��Z9�Q���x����:�V���M"a�n2�}~A�^�6�*P5����3�-�`��t%:����ḕ=Q�e�f>�Z8?pH����ay��ZM*�L谢��_��v�E�7��#~8c�r�_p���/�'�'������*q���Ϝ VH��e�:�%������D~l2zf4�[$�����si8�U�O67��v�B0�(�f�B�˴�79r�� 8��}k��G���;t�����wN,�J���Gw������~��N���'?1x���m����px~RnHO �F K�ek1�<�tb5U����S��0r`�{�M�f>Z�
V^7H�@̯&-c��P9�Z��͉����<��9'�+/�J�B�xS����$	�6�l�4,��v�ذ�=(TΛJ�.�G�0( ������������BB/5<�j�X/��.�G�2��Gl\�bipEQݤa1�̎���W�M�gna::��e���l�Pd�S��ߨ^:y��R�}N������� )��������T�)y�nb�� � �`��ƅ��\l|��[�Đ$���N����u=�aQ S��fa{�H�	O�c�.���pfGO=[���m�s�J!�*Hש*X��-�Df���x��IO�m�b��}pPyl?|�qr��W�/�k�'��1Fth�V꾦��{Y�h	��	'؎�����2;�2����%��.����oI���x����Y�},��!�ͤ��=����3 ���"����| MNy�W���z�7�>j	�&UE&��G��AS�;�xi">͢t�LI�1���aY��zJ�{)�f�� g��NQ�[��]�� )�.�2��R��zF��������x\���r�;˛���p|�9:ej9�~}��y��سDx�8C�	��e���S��6$9O��^�O��	���ض���j��,��x=b �����y(�	0
G,:�*2n০�F ?�K�4�����z0�CY�5�1���q&X`�m_���Y�����U��X9���"s�↑� P�2��V�M����(3�R�.�,���Շ�2��R{�U�
f>�aE��K�%�
��,sx��F���C��U��6>��g$�5��G��_��]��HI�lU=�Z�p~����p�\�W,'$
60���e
pqT���Ka	M�0��\��d���_K~Q��s�T��gN��ϒ���\ڿNS�N��4��7���U���[n痓��Ҷ�3���A�>�ma	Yx���)�C	�I��de(�Mgݑ��(�ކj�ѯr^֞��MЎCꐊW��ե���		1R�ˏa�h�1���d���EM���N*x蘊[���T>���A���m���څ�L���K���{������w���t%O�lF��{'�o�W��a��OE]����`}_��b�� 5B����i��ކ���j3Bm�\o��/��0��;��5B@�܊�vN��1��tB�G�ː�W8��x���X���J��y,NH#W�Ȭ�������9�fbo��O�( I�#���k�o|Vv���sK��'#M����3��!��+H�'ï�4[�f.M�%Ti���X�t�V�P��ro~�wb��2O�ȄW�H}H�	=�赗O�jN���3aH�S~���fS$|u)i��+%���q�!��=9��:Va��m�}V�7n�2MfȾ"�:����$��˖f�(�_a��̪D�ǽ��#C]�\����UP'1���0LJ#k�^FI�mR�����0%Z�N'B�mҧ"d���39�����8����T,�)Υ�E��}�
q\��p�QA?u�l'��a���L}��HIPxDPǀ<���]��/�m,����S�[�:
f�t1����ۥ�T{������\S�s���^;�i�N�l�P��KJks��l����!-�]G�t!����`�<�F��-����|�%1���J��̓8���eHT�mN0���.�1\~(�E����2&��AO�׭ɑ݌n���{U��z"�|��d[�=�xŐ�h�[�鎔߶[/H�']ZX�>Ŀ��#5t���ڊ<����),'rtdX���q_�~�b:M���Ѿqd��xA����I�56��C(�M\�Ń}>�HO+�<*�z3�E3��V�����hq�Օ�à+%���nu�p��u$��T��J�e3��!8L���%+�j��}ئSAzl�X~8�ϒ,9B�-��km2xq�CM�����c�*7�C�����T+P�&�<�@���]�/[Y�'d��c���1$޺�Ϝ��v��I�C�a�s�z�IA�|����^p�!��LNr���t�/��FJ�E07���H��x�#T}��z�]q.�/$āV�Rzkw�n!�$�
��zG:�#C��)�ww5���pN�zO����tKo�X�"w�m�l`��y� ���<B��F'l_� <�+���'l '6��@���v˻�Q�*��伈�\��v��T�!��u�u���r�Ec�c�o���d���v�2X��=]|g{�Ƹ��B)������k y˸��4�D/� K� ������gZCF2�,� n3AѴ�X& �QvN��<��b߽���bG�a��ZqgW��h<�X���8�2`�œ����J��2_�H�^��;t[��4���7���\1�4�S�~|����IȾoIE��đ�a(��~��ߡ��`�v�<E%�-(��w�vDA����,�����vO��M6}���l��b]��}�{j]�f�r�ݸ`�2l��V[3ߗ�a��L��XJ�/4�V}"8<$
�	����|��h��i�Kv�k����j@nh�_��_�ezu3@,��+L�m�v��XA���^�u�eS���<�b�-���"8�Yk��-��]��?�:�{���S6�N^\bw�n���o�[O�S9!�[\�uH��'��BR�W���p>���~bh�B�0i��YB �!��'�q	�
�%g&2�����dA�YA�{���I^��N֤�a]���C���s�]t��3���ȞX-.���=O� ?W�� ����N,ߦ�@��4�=e�6�&������иF�#��Kr����6�w�\�7����Y��l�~0i��T�-��?l�����V,g���om3�>�:^={�,ڿ�a�ƟU�y��"8�>J�q�y���٩�v�r�U?Ҍ^�~U�B��0@� +Ii�FՁʸ �M?c6pz��i������+�v=��NDU���	jN=z��?pC�]�mK(=�=�0��c�@#��2�0��N::wc[��&BT����S��}^ e6�G8z��ۦ͛��3��)�JX����Ӎ���?�~ӤVJ�wR��2B���D��h��/j� �3ƅ���Vv���8��D�3?���/~O��x����$��|iI3q��=���Y�Ǻ��>�ݽ;J"�S�ٞ��[(�e<����1���>X�y��bN��T��6�z�=C����Jvkn��w��}E�	̛�{���^x3DVH�̅�!�n*�ťݻc�\޻k}�0ɘ��}��h�%�y�)gS�m�.GF3h���h� -.�C�<E���K4��h""_!)wCz. �I�b��!��A�v|�҄��=˘���8A��bC�K&Fż����Y$��Խ� g]��"�DD5� ����A��/'c���u��Z^�J��O��
�n�+3v_9��3)]���>�FL��A`2�6:��X�AZ�.ِ�=�7�������@�*��(x>��6񪞢n�K1*�0	�Bʓ0,�Tp�����9rg��w���I"�	�Lsޘ�0���e��C����G��';Q)���X�|�$SJ��]�AX3�}v�����dH�.��d���K�bw�@3�{��q-������om&���t��D-x�A�?je�	Q�O{ !/C�B����߷O����W��Y���/U1�Ș�b�~��X���O�H�,"�RtΑ��� e�o��u&4��oK�	iLV����zI�#ػB�i4�|9��O�m��Xپ��1�|���r�.~��I[ng���j&��7N�ɞ�ٞNę�]sef۞�u.9��<�wT4�ץW�y�([(��mQ��L8�b�迢:$}�e�^��Ht�:�����T��lk���\��_P�6r��1��p!�*Ǟ[�ZBs��̂;��)�F�6������qd�<�ڣ��KԘt�)n�k�<y�Q��D*�]���P���OF���D�%��r��b�Dg�ފ\2jy甧լC���߀�s��\��Q�ٸb�* ʴ#�^��r��mx
6^I����z-�L q�{O�#���Y��~C���D3G�o�l^��^%�;y���a"�_�p+~�U�%w���r�۸��EEM�C2���O�{4"���=�݄�Y=�e��Ň��@�Yz�0|+�x�_�,�mM�dw�
��W�T)��D<�Jt�@A�+N�wa�r�vH����3��}H�'���ȩg����Ȥd�vS#�L��9�Hq[֌z�*�(J�qS����̙��͙ڻ��g#�F�o
��:��`2����Ұ\��7yl?$<d�p#1n0q�֪�!�,
v�|�8Pi"b@�)�_sK��N�u��w��Q&N���}�lm&�P�׀�O.8T�A8X�_0L8Krn`	'J\��}�2�#�G�ˋĆ��O�Dt�owd!�a���QG�s���I���O�Ϝ@�4}��Q��K�4#�H.d���S�t��gEϋ0�V�I��q�m�3[q�,�s�<�ȖE�ʙ`w)��Ƭ���'t���~n2�-�mZc'�u��6��D ��p&N��4{*���&Q[G9&
8�����6V>�%�q�̧��%�F�gF �,��.��������m$/�
�Gp�#���g������'v#�y�x�)����_���>�M�J������aw��W��QR<�JRV��5q�/�df'E��qL�k%JR�>P�j��W�Ju��ԟ�<TQ�^��0����:�Z�{��p���Z�lB�ռ�<��b��]�J�89�8Թ�"1�^zb��C�}}.��[ ��9��f��(׆��}e�e���'E�������-�j9-P�c׽�s�=�	`�i�"B�0/�/8í���"̷8�s�c�<����42�o��x �P9}�i�T�L|ȍk���<4 �0����_�p3�����7oÛ]A��/�MV�yO��T�I;�z/�¾I�j8G� _zB���cP�æ������[��`���@f�������ex?�Y
��>�Sz����a�E�WD� #J��z�SWo�l��*�nko'9���&ɚ�h���C��P��)��F"d�O2�|j`Y$X+pAs��2l�(��yl�_
�`W�m���%F:Wq���GBPp^��eao쮅'����6N���f[qu���S[�����>JC���M!���v1+��ux�(�r�m��e�˜�HBMe]��?�����^��$$v�.���Rx
�e!�]Ћ� �n,�3�HgP-��.�c�}�'f���4+�5(�+K)���Ӷe�7���!�#�`1}�*ه=�q]R�O)�G��9ް ����6��x��=p��DaV����mj�g�C뼹���E�����j�D� '����2/��ʩi#��?\�t)*�!��&�)f��ؖ������#�v�U_,>�@��=G	)2U/5ާ������l4a�Zhؖ�·�"�JI}ePq��ȜAW���ǭ��@��8p���UIa_3k����8J�v��o}�P�ٖ��{B�3��Ҽ�ȟ_#R���9DRn�N���4n��fC�����W��k�YŵO��v��F�ͥ)E�:I�Y�0�Yy\!#�ޛ>�^{��M��|����ԙ�S��A+�EG��a�!tǇ�������/��S�	�3��(v�fH�x��	G=�ߙ,��Q�3K��v��m��JC��t��(�o�J @���n%'�)�ϴ��r�1�_3�n���љ~��	�{1o�yO���P;��U���BA����vc����xB�_������]�V�/?�˷�ο�q��:����_��N㠍y44�X�oV?Fr�X�
1:-@q�-�DK@N	�v�ŊfT�<%a]T���G���,��pʅ���w�2~�E0F��K�a�Ah�,w4���@g����-���3�Ԏ펛�ʬ3�_���`��f��l�~�&��?�J��\���8mL0.��yѣ+դ.k겻m�f߾�V�a��>E���� �AA�+�C�kU���S��Ӓ�C�&��&4y�8%[û-s>4S��KS�rN�����i~��"�ǀo�/����a$�¬�3`�����'�<Pt��G����+�MR �Z9�"_x�aF�ƀ;���R�[��k&j���v�\��[��mC�SM��s�,�g�ҳ��XX�� &�v�>��ѱ]���5�E��i��'�C��8ts�(���H���9^���cU���B�X�&J������.�F�V�u-��QL�q^h��18-�z��	������P�l
�IG8T��LI��өq�WM �됆�R��f71�3SZ$��=�����@�mʽ�� D���T�ͦ�GGM�:��+��ٜō��.�G9M�!z��B����?~�W�,��OV&n�b�/Fΰ��~��&�����L���%Xx�\y6ێ�6�)(���ْ��_1N��!	���eP��i�����>���{�����
C��-́�����@vD��T�}<;*jB/���;=xo�>ԭXc:dY.�P���EF���V��7���se���i�w8�;�1/ׯϧ<1�u����Z�HH��}� ޲�)�I�����D�|5h)�d��KW�b탡���Fwn6}�"Z�c&��bC:Bg"�l�Z]l�(?�p|v�qiVVVrǵ芇�d��O��.��j�6�蹊�Omjq��b�~H[@�5{bG͂�	[��{���yD>�x��bN�W�&���鿥pZ�u5��˸��1��V����E؆�V��w?�r����aq���X1��'��?K׼j�W����H�����E�-:&����� ����Ud�t�K�!��0�Q�w�B/T�/-՜�O���E`M��u�`�K��:&)c������>x�v�S�T�|���� ��<��3�Z=
3\>�{���s��Ri%��qm���Y�[���N��Р0�h�*�t�5�hh2����uX�G)�Ʌ�+�k�l�X)|_;�nD��=1� m.��K<kq(��lX%���{�ij)V�DDs#�&b�C M��`֑�p�Yw�Lp�Ґ5�d�g%>��*�u���ޗ�>�fk�ޫ���|D�}wP~��_n�K���b�	��Â2Y����2V�,/�$Ԕ�б�<sCU�A�U&zkx/
�b��z
gT
�m#���Q���*;X(Z�E�b�����
�����]�J�GE�i�w[�~��ma(��(9���cn#�"qJ�d��:��A�75paV9�BѺ7��qN���9j�/��{��կ|��4�f��٤��Mq��׈e�~T�HK�����k}WHY6�h]�j��X�5w9L!���hB-��x��E�B��z�$�Z�4�"~D$>L뱏�}����][�тp|q�K	�u������>��'-�zъt�	��-U!�Mf��-�Y��qP��`�*�W݌�̂I�����q�e��K�~��!D���\a�:>�CZ�û����ľ��3}���������3Xk2F��U��)�ӷ����ȵ���X	mf=�Q�f�,eU�������HN�E[R"�sq��7�l���[��8D�%�Pr+�5	����o2�$�F�f3�r�o���5"Q9:�`ո$�q� �0���M<��A�������y�^+�o�>�[�+!��(ǣ�1���Ue�����6��:����)���Y5�.�Ң
 ���,�ks@�UŃ�� :	�'>QX}ęg}z���DEob�u��"�� ��Ie	�G�1,����QG0� �[����w#��n�z�SAˀWD^r�lDz��p�ڀ���Z��6jv?˼�+�s��I�P��m�q"��"��F���h��w�BFJ1%��-6�M�73&��f��W%�*�������E�G~��+�/Fn����c���z4��sug+�,���D	`�҅wy���s5=+Y(��۾�}2Qp�bvP��ע��b��E�AЪb�eGl�i���wcJ�&�?��\ۼ��=�����_s ���*uhF���]���L���Z�嫢���ۂ���H��Dq����b|�lU>�*+���k%K��˞�H�U�ϋ׌��īc�~c�a��/ܸu�f*��zL�N9V!������C�l�}�xcfl�H�'�^P`<�w�ZE��d%~'�N�b�+03ع�Jt�N5�+�_T����Sh��V��0r�+�US���n0al{�D��%D�E���|�?d$���T\�і�q����<�;����Ƃ��봢n���}Z{T8�#W��*�����*�9j �U�����I�\�턡��D��E/��)�2:��0h�e�t>w������՗-Q��& 70aPI<�͎Ht��}[Լ8�o_���ũ=�B���%W�2 ��8N�h`�[!����vO���8g���a�(
�D*bfaĈW��h�������ձZ�H�M�H��X~�N8T=��	JY��j�eS�R�P�iK�|��?�;�ё�K.^������Ē�^�::��u@ԛ/J6����;x����.i�o�e?)�
S,��:�O�?�������ؠ�-�܃ļ� H山+��ɽS�!����ﻫ�!h�%��N'�)�s�S��:g���R��i&�"�Ak�#��snҀ`8�.��E�r�e��m���'��9o��b�����e�B�g�.�յ�)6�v������a� ��9*�`����c�J������s�d�x7�1����T�W$�|������Bq9�4/?���k�<1A3����*�#Rw�=H3͒.��_��NJ������Fc���"�o�$�āh��e���#_��,b��f/�p�� kg�`L���)؝"Y�eXNoL^�΅�#м�$�Kif��"���*�����!���e����U�kG�B���-���	�l�)�!�x&�k&،�M)s&9����^)�a�}�Ƌ^�ObI0?��"8�^@,ǻ`;{��@{{ێ�6�����R ��{���Q'��OF���H{Z��on����ĭ�X�:��u�	xD,C-����=�ƑZ�Tz�'��@WN]*CH�GIV
�d�%jY��%���Tu��!��\\��^ͨj/�E��x�A�Yi�Ҡ=�m����'���R���B���x"G�n�
�1?&_��0�!����j��ߢ�x�bdAdP ���Hh�j��tb�/���e.�5���)	r+�O���8��������Z�KP���9I'�p@ �r�X�ڶ�0�c�8���z����Pt�7��]��[�CK::�ef�����Z�eR�h���
K��?���?�|y��V"�F^��I�|�	:��nx��⃛n�Q�'����(�4<q�$��GJ��E�6���si�: w\;AY�[S���@�.JS�t���4����m1ι�b��r�x�~e�ݵ�6�rS�n���0M���\�r���oz:�.�'���%<ǋ�&��ܭ�HIѠ�V3���D_*8��Y��	SY�OVrd7$|�`fv���wsb��V���YA�ӰC��s����7j��	[�1j�6���6�+FF�a�������DPk�r4��VN�&�>Aׯ�%FJ�gķ�)<�OI5{�]�0�s]�L���3[�b��3�(5'l������S�M>6���%BV��~���c��k05CK�W5��)n��rC��cL�`�Я�A�\�Ցl�H�V�ڂ)P3�A����_��fb�Y�
6���ozt�_��{�sم̋�>��������"*bޟ�7�..^�r9Bi��_^|k�quv�����[؋���f��������e9<B��φ�Ȃ��Џ�	� ��Y�""�h_�Y�'��`�g�_�<�ƌ��~Sƀ��SG��(�7�W�"ƀe�b�Z3_ۘf0G�=�ZG�J�Lh_N��ߜjVm�c�`V���T:ÍZ��!"Bs}�(G�.:�V�@i�P�S.�8�M�>�?p΃�{��9�P�sy�ӳ�ogv׽Q}��z�M��T^mr��~_� ���� m��ܕp�D�6?Nr
ƗrPe5"�J�8+�6���SIkaj0�-�ja)^m�4`��S��[n���W�Յ?��%���ʲ|�}u��q;G���zår����%�x �6�WD-�:��׀�6���3]���q�^�)�e�D�p<3�c�3�<ŊG&{��>
W�7�F�>qr��;Խ�l��*d3�dw����(LF�[y��@-6������P��;@n��|�is�ʾ�;mrQ���6g���q��,�v�t:�UN�	��^�?}_n>c�*�Nb
������Qb�ҽ������<�@XW;Dc�,� �����;^w���q��kAԌiԶ}��i$�v�oŐL��0 Z�\����yu*_�ѬZ��$���UFق�k����p\��j�oP�9��]��w񤪙T�k&G+�Q`DnHw��s�T�6��
�����?����#[��=��[ C��V�"A�:�
�0��8��R<�PoM��t�t�~���9��d3���6[��E��5{��'�u�d|_��w��TI��8��Xl�ZT�O���8���&3TL����=7��̚8\���,�����k={��e�H����R�Z+Y����E;�*�Yl�%+��'aXk���'~�^.Q��vq*���X�ŐpW�c����\�:�v@ �����څ/�a�"ժ-,f1W���U����ec7ب�L�E���ݙ�ۍ���P��gt>�Y�	M��izgS��9SAۦAk�/^����k`���~�(�F�P�����>_Zo�D9� ��aSj���zz�b)O1P���-���S��G`�G2h���7�^�������>�74��K[��lR>���z�4�g�5&�o�ilM�-�W�l�b 1#�W�[}�HMb�]�@������K�ժQ@"/YqL�Ԇy6�����P��bVi@7�ܨ� [N\��Ljm��[T����I8��'U��Ɓ.t%R%�2�Ok�Pw�����&���>���5���J+G>1��/;#��r�;���&�����u� \���)=u�8�5#)�.��5-q�6[���z�C������;A4L�X����V��c:�+8�
=��~�v��!:R�HyV�ye!��x�{/��:H� / ��V0���?&����~ڛb�rQ�0��]�(�ܺ�ױa�j=ǜ�(C�%U�:d�O�n�I$����=#�[������U���-iˏۆ+����=�ʪ����Y��}�X1���鱀#��"�e��*��st�xF�ºՔ�̅����W&���t!Ъ�0����:R+�Ch֯��o��N2���ZA�#�D�3&ߘg��i�ydB;�޵Ch$MO�LB`L����R��/��#XC�V�#�F+�,2ū'�L#Q|\S,5��8����o?r��(��k��xl ��Q ��o��ii���(�|�8�Y`bu��JG�3�@U�Y�>�WD	���4@,��L����Y:4ߟ�Lˮ�;�0�	�`���]���vXlbu.&�%Fv_T��f�-�0�4ͩH�͍��Y�P܊���`�Q(oх��q4��a�R,��)�z
�BCt�-%����M�����Yۧe�R��͛���-�� o�'�V�'>��F\��HD�(�xA�xv!j�N�#��W�����g-����;���%2pHD�ߙm��b[ȋ��؀�
��$�OD�����C�= �l���?�[�PHR���9��3��aS�0�'݉�����%�y�JĜ5bF'�����g
���4?Ű�hN�50L5=ݢ�|��C�mA��fj,��m��u�[����k3""�-�S�(�@P��a1C�c4}��"~
U|V!+}��9���K��<�U�����;�. :�n>�������D�5�����8�Q4�m@��L��O���O���+�Rо-4�E[�;�b \�m����tm'm�|��������G9֋
�F�nK��2���-(O�~����4��F��Z�L"q|N��\���h?��]�37i'�����BzM]��B�$BA��IL�݁p��K>ô�*A�W��:/_\6V�	t������ѻܷ_Rm,Y^n���J�Q�^P�f��4:�KIl}~��'ˈ�=��>.���˝s��iKi�y��U'3���6��C^����q�\�\���q)V6A���t�sG.RR��K���p?�B���l���M��ni���[f�,t�J����Zō֩rt\��j��v�8�s_i�j,�R�P�8p,����PZMtW���
./F��(�ʋ2U�8u+Cx	��J�W�7/�U܊4PSOq��������O�^)��zQI E����h���1���tr���
�MhZ�2j��(�R�:��0.Z1�5{��v�˿8�k��6�nz�EkD�oZr�j���Ap'Xk�����M�1�)G�	�9���v�k?Y&{�������j�>X)���i�a1�ڗ���
' >��f�兖�|�	�P�]�a���r���l���Zb��F����)���/�ʄ�����jn�o��u���;�Ĩ�E�a����Gp�x����P����s��~�]�H~���'%|���M�2��Z�ʶ'�@�m�-fC
�3��-5}��vh�ƈ<i�2J:8r�F�U�;�hh5�"0��z�"��ԼS���Y�7}���HP"�Y:��rP2���Ѝ�eBYODl?E���9K���*GU���8��9�Z)L��V�yv5�� ��.&ԄU�Y `��)�gꊩS�\1��ͅ��D(�5�D���4y$����E��i�����@$&�5L��z���{�K7+��*)�2�B��'��Zq0E'�q]�O��p8C�����ķDK�wE��F)(y|���I��~7�QjoP)Y��'i���ΰ���4(.@;��i�B��?���	�Hϯ.5U���l�(��fI�8-�1Ϸ���l��eOf���Y���&:z.s����\�Y(@f!u����<��A�4�ރ�\��aU�U5w��"!��e� ���A�xh�o�8��\��T�^e�Q�x2`G떐8]�tK
:ũ��Ña��c�� Vu�	�t�*����2����.=M�*����~��Z�P'x�F+8���6W��e�	�-����mh�>+m�g�i,e�)��Nn��s�O���+yiDj��̐e��_����h9M��aİ	��f�[���{5B�m�4h�j?��m��L���͌IH7��+�y��8�y��p
[�ߖ���v��L�T���P��]Y7�\�Թ���I8����`�Fv]�cīu��4�e�>e,���p8��0*,��N���l�.!P��^�i2�k	T�xܷI�����2NGG�5~ń �/�}]^�'�a����Ȏ��>��F�j��5��5�RUT�"��pr+XT�6��>��u�j����xn�ȼH<ج� �g�ى�J�d+�4>�g�Rs`3]�??6�<��p�O]�3��
�g�u�U �<@�
���'��CKL	@D����[b��E�\�-(�O_�э;|�o�[������*9�O�}Zw�faЧG��PZ�b���"�8�ß@D
����8��o��bVrDT�@���RA%�nvBxxM���N�q�Ҡ1������w���dg�c|_���B֎<O��g,�tT����Dîn2 ��N��Uu�BhP'V�/�y��q��Xc<k��MS�A�2��o��8ւ/�F�L�"h�)�ԭ��ܪހeI!��4�2zk�Y��Ӱ��c;ƀ������2��Q�>��"=DUTQ�tk�}��q|�±^}�� ����6���	���:�+0�j�:�3)��{���s��͢b#׀D&/&E2�Wz��(�3���fPU��Hb�bg���.ST�����d�T���R1�e���^�J�^T.�zZ[R{������D������?e�R��hpϴ+j!�w�8�ȓ���s\l&c6P�j�-Lk�C�����?�U�u8�Nt�¥��1#b�m'G[�lg@9 �7��٪�s�<Rמ��W[�Q(�?p*���H�V�������<�1ܔKs�Dt�]j���-���6�R9�A�㈇#i�dO�����pd�^j���%�F�!H�	�+�x?�od�m�@�ȡ�Ԗ&z���I���$��ФśMn�-XM�b�Iј��k������6X�m������u_�P
/(�]��Q�c��n�T�[tz�_fj,��n���R���V�"����YgR%�Y�/UN��N�Y�G0����u�m}�-#ȢfGH��ǯ�+tY�-���as�3qV����ݲ�=�,����t��3��̔B@�\p�E�	�ݱ��P��z�������E��ҏ�h7�Mr�!��*K�2cm�U�s.l0���6M��Pff�o�x%.�O����Y�SqxFe:�Ro����ٍP����<ύ�������F<�)��{�3.�}�hW¥� �75��dp9¼��_��P�e��84��P����o�j���o��\��b��.�"�(9�mj^A"2p��&0��`�N��y���R#|v�	 G�/���F�ܿ8CΤ2�����C�]X��J>�z ���f�G̙w�J�;,hT#؃��%�q;�t1�?1��x�ZP*�^u��u|����U���� i��:!#����h��x�_U��T|�d��H5,AȜ*�*�迂0	ħ�t�O6?��O�����J�J�>ʾz>s��^D�׬��(xf�5X���o
��Y��Xw�z�ך`��|ʳ��ꄕ��2�+�Y��Z��I4����'^-:�x���&|��z�n$�3WӚ�.���n�A���>�ئ$���Ɂ1NS#�`n��LS��|�ޥ�}l� �Ԫ�/E�=���<`���|�y��4cOetк������A�Kˡz>�cI`*��z��]�~ݹ��E�,bK�n��Bewg�4��c���_�)"�7/���l�`1et0���>d�e�+%m߶8��@�� ^�Ә�����]�xҩ(��q(lп������]: 9�\�vl��^[^G�i�%k�Ra%�!�h*��m����D�گ&�*MZR[k}2� oLrŀ�^ԥ	%{�� �����x�a����N�D>q`V�A7��ٷD�)L{��tJ)� >xO	�m����p/��N�]M��Y���tB��F|��=Kq^��ץ|)���m��CK?���w�˺
�$���0F¹䗟��_p��A��ո9��w1�,�7|35�bV��OY|>-�c�1c�a�����K�#�G}�@�?����}Eo���|����]`*�^�"�T��wެ�6t|1��A�~%h@��|��jv������-��`�{�w��hV:3X$�T���d� ��v,:8Yw�e�ٱ=͙f�SJ�v��1qB��,n��nC[�m��*Q��Bz���Y������4 ���� �J%������f�i�:�nw���/uz����N_�U5n��IO���h>����lu��/��QZ�'��de�&���u������h�����)Q�=8[���Ip���xJ+����=��А���˫����Nm��p�����Z�Q�������lp�����w��z��'���j�����Ltá��\�lTB��w�xN��L[�0�t�X���C>|��6�y@i�ݣ����?��@��N�b�P@^V��nf���-�@0�_��O6�աs̲����lQȨ�;��1�x�W��;(��գ
P�$�ݍ�U)�C��-���a���ct�}�3��z�,-?��)�� ���%J6��ہC��2Xl��	����'R�k��<�)�f�u\�I\'a9pO@ͪ�L9�TYL��~���χ�K�hz�|��ګ߉-<t�V�k48�Td�o*/�x@K�q\�4�6<��J@�Ϛ�I(.<�NX�d��1��b_��3���ֵ�~��W#�ʉ>.	[�,�*�>2/�>ʺ��!��7��J;�|�1!Hpԟ��.�l��껙{�uAq�a��Y���[�Z�F��u�š�܅��A!w AH��%�(��EyPs}��Jܙ���A_5Uz������Z���KNK���yc�z�`d��$��9Bnn3;�\�u���5}A�����͛��1LY����S�����
�u�U�8��>���(M�e!�i��t�=6�O�m=���w���k�>sr���jGL�<H_O�jV%�����I�:I�3��p����
t3��<�<5�=W��`�<4�׹��j��~ڌ�U�$ٲ��f���`�U���BKd a���S;�Y�d�>��d��nV���uD����R�{���
�8�7���N��=�b�.�1L�:�W\�'2�f[�-֞E�<�m�A!�S\�3�[�&#�ߗ��,,��1oP��n��8s��m1��=^]F�����;�6wY8(o��VA�C��T6�y�)��<��V6�;�B�/���w��X�.��B��x�D�2�&��[J?��Z_�mP���{�e@���f�8��u"�����~6j.<�Ó�R+#��R�����KЂ
������	$O�K�|nvPj���|~�������r�)P%rUz�c�\+�[1z���ia?�^����#�!Ί)?A��ʣs �zH뮉*�D��H��q"�yj��*�7[Z�3�lf�v/�������ikb�O	���"�B�`N�<�$��Q�%���tڤ/4�mihd$i;��;�`z��!LU8�c�ǔ��9�=�˝^���V_^���4�U�s��?��.L<�1
�>e5�.t�}�es1
�u���1>V}+�%�cj���Y5	�< �*�i�-0�Lk^��|�p%d)�C��;E�z#��d �a�ϼ;�d�+}/MIa f�q��*6�?��%��,�ܰ��ٱ�����������3����C�s�������z��[���2z�}Gz�dM�(�o6i[!2��A9��.��8JY��Y��$�%c�v������h;��	��]bÈoj�ɢ�!��y�.2)3���t$@�U���Z���[��w5p�X����.&_�C������,t4�T�qHU_� �j$`� ������h�>U�p}z�{[SK6���=y�����կ�F�ׂ��R[�Wj�~ѵa��qr�t���	_�x�z�{Ly}s@Ŏ^����dHs -��(�Z���ڙ���xx�8^%M/��p�e���q�߼��v#`�d3�J�A�a��.}9�9�l�g'����/�.j����4�Y��b�巅����wW�$�we���B�ܰȶх����Ƙꈣ�7�~h��� )]9�ZSv� �iY"� �N�9�612fCg�bgD��B�8_�L/g��՗�o'��巵�*cЁ�_a�Ӯ�.�%��d�qH��9d��t!�a��Ƥ��A�V�O��2��Oq��&g���G�`�-;�:@1�y�Q@�E�eP�	%�5��i����^5�Mc%�:�
�Y0r�����A�_W63F){�6��y��'��!�(�f�奙XՍ$;�!��Џ��^/���V�I�l?�Z^c�A����k��Jy�Q���;�� �|�� �/)��!�#�	j+�{j��H���F'����ga����^�������pd���GӶW��G����Qa&9o�Uvi�� \y����e��p�2�kE�񻠑طR�*i!���b�
@Y�O)���18�����D� g��q~���섚�$�^M)���]`������RZa�S����ִ>��5������Gi�֐���h1�<�&��9,��š7���T�����e�>���@̞+A ��=6f�rw�c����z~��NYS�9�ċ�:*�p�2$�����.S�l\�$l[�λ|}�W9`7[�)'z7���ø�̝���`����U�EU������o�����y�l��P��ąS�GXw�$�-=A�K����d���]_Ƀ���ڹrq�e�P�����_�1�i��W9�Y�y����Pg9Y�����͒�a��	+��Ȫ���]�ʳ?T��@�����^���r���kt�i���l�P0�}V��)R��|��x+S�6����*Qf�	�ʳ����C��K+�6,Ӛy�Q�I��a���nvm�wY�!�\�'��;Ȯ�0�����'a��k���"+�k�r�)�Nx�w�@%՟��"��\�yG�Jj::&��|x]��Y~�ي<�a{�� ?�:�A�`�4.���ei��1�;�� �l!�����!���E`G�jWELa�����B�膾+�5��n��������e�-Fm�&��GO�a�b �ޞ56o˘.[��B�c0#����.�첈E�Ċ*�;(*X�8�?�*w��������O��䬏�wu2�K�pl���`Ϫ.O[�;<�7* ,a6i~:.��@�e�p��kU�۫|�7.���=�/$���6��|�>���I����u�Y�M���,��G�������O)�dV`��v���s����WE*��83�y�3��'�\+&��t3C�e8.��(CV9G9�V�Q�|��"�ss*������\2}��Nr1)�9�d�*�G���M(r��A˗��\�q�1�"EmK��F�[R�"�8�u�F�����b��پL�J����:�y�������vzP�fm�9�`�� �(��ԋ���a!�IQ�Ky��}�n�L�4��W#�qݒ���>FV��1۞��֕}� ��p�6��?ƺGf'L^�M��@i�j�E�b�̾���x�k�땝٠�b*�޼4z�̏��a�n�Ear��$:����0��"tr��ޥ�W��?�"˔_�bK�����%('�C��p¥s�mZkk�z>������m40N����E�c���f(tͽ�z}Pg5��N<��W/�͉t�o�y����C�,t�	���G�Z3ߌ�or�"jŎ�;����ř*�Pj)߭at��c�\u���T�����[yv$������0�?`Pf�6��/nK7�\����]�x�G��A�+���������d跷?iρ�XD�q��b]'oI���8ޫ�k=��'k�{Z��4���-�"K�͵b����M/ �dX�I+��b����Q*���_u�H��[��pA�4쒃�ᪧ�H���Ɔ��q�l���
�Q����٧��	��*5�@����x>��#��:�wx4>Z���2���:Y�(dy.��L����o���*b�Zj P�ځI�	̀/��ῐg��b�H�S�����d�&1��/=�o�̑F�Ä�I+���2{pT�#M�o��X#B��:8�sL��/YzL}_���+�Ź���M�1-8��M��>����R��\�������>��|
S/1Ė��Mk2�2�BP�^��d������b=ԝ��9R��Wո#�ܬԢ.#!�qg��&��E˻��K-k{���?ٳɿ����0�'Ni$�_q�`�P��(�b�����S���3��.���=Ć��J2{�ءع���j:�O�,!�7�SY�;UQ���@݂u�;�~
k��W�
i��,��Rʥ+1���olx�	v�6�_c��67L[�3�������`���M��{,aBŷa�#n�f?���\2(��k����-�fM����.[X;^�]u�����cܥ�n�F�ƥ-E�� ���������v}�����7��Su"}�A�K&UП�A�8�A�]�8�Xƪ���C�s�O^�jcZ�JY�gz"ټ�6��2sX����(�-r�]�c�C���r�4��&�"�scLA��of0w�!���J6F�t���5�2�鍉3p��5�a̒4���}2E���M��~j�&չeU��u'|`r65�[����ʊ�%"_����T��#�"��~�,�`�[�d��6v^A�)�֏8ꆯ�re�m҄4��dZ��	0�<�e0|%C��
Lc[�xk=�G>S���P�Al*ꚁw+�+�c�k�j���9�%�p�����<�x�)�3���*���ff�v.���A@�-�B�� ���.��=C���\�əP�gU�_��,>~ �Q��}n�+����)�ȵ��@��}zD��)`,ޚ��.��	0�5ԅc02� ɉ��ё0�*P���D}���+�4z]5�["5M)M��6
������\�>Ao�%*���{�*R�ovo^9��qܷ�/��y��\SL��j�Dp���.�d�KY�����G���+w�R�}��$V"�?D[�Nr4��7zOhi2c1	�Ɛ!12A�����:D%�_�aAp���Ί��!0$��ꞡ�޸�@��t�(q�G��|�O����!�� ��}��Ո���Tt�����A�RJ:-S6���/����V7�g�B�.ˑ1oC�!���R��\�A1���z~0�"
�j<��I�E�52�
�ہ���
���GP��Fu<��=�D(6�R7�����fg�d�-������OHc��s��u�'�홋�)�k�7'�~;�8�����o�|;��cې�Y�W�+��z��p�Nq`�c��%����:�-���Փ�1I��B��3��|���N+��V�5 Rl�l�LneʇY�UD�� 4�V�=�?C9]PJ���/��s��P��m|Q�o�$w[^��0fg�A��!z�$��;�@�}�V{���"�-O��vz6�Qh�V�p�S�_�T�u>���#���W��(�Q(76~���~"�p�\���K�|i9v�-U����Nc�#��	������lL[1W��{�v�D+���i疡آq���ʤ/v�1��j�8�J�:>ˤ�-m�#���Bv�)�L!�T�Y�]H(���@-׋F6��k
�}�, ���̭���[| �\�@�H�%��{m��\�?�L�	� ԀX3nq�Dv�c��92�(��T[��m��٨��"gDāF폪������zY�`��e�*^JӦ���Jɯ������4����N�q���������c�,M�:��ϱG�S��ו�|��
�'�����G~w�:��7ϻ�JJ� ��o
�L��5�L�:oC�D����s�+s�KlpӋ5Y�p@���xC�e��b��>�I*y1���2_�����������D��'xf�m�xe���4gt4���HX�N�߇8�v(j��w�\����撯u�Nڀ4~UO�ּ�_-@lX�9 �a
�!���XU�kQ�E5,WE�:�=��5��,�b�`����ɃB]�;ê���:��	��8e]
ˑ}"�^۵�}6�S��P�+������1��8�����[L�&'�I�0�N��g���3J���*)��v�b2uEVa�C�S ��T6�k�]�b��*�Ġ���c�)�qU��{��aj/{,`���9��v�[��SX�`��1�(��3+�p�3aٷ��o��
�g���:��dn��|��Bt�D�D� �jG.@3��`م�2IV$[�5=� Z��L���w�?�:#絊1v�o��
m�I��c6�7�P
�Y��7A�hP�.B�nk����H\�p��+MN>Ke�Z���X������C���9I����E��g�	 =�1���)�#B�[��0 �1�Wnl�|�"|H8ϟ�m�].+�W��Sk�?CF��O���l0^�Q�Xv�r�J_���F��P߭&q.��`�ε04�w���717)Sp��HI_��i�| G�}l���h��RP"�?��8h4؁/n�Y9G��,�+ˈ�ap��F���	�h���a��T����,� ?Y`������iұ��F���Ǡ�_��,].��b���G3��ݬ�K��p�����n��vTӲN*i=��������	�F/aOdv/�`K�����~QU%���`�׶����Z���7[�1�)��$F�Էz��⟩�����g'C�GN�YF���Ӵ�G�([�Jd�m�ۦ���K����]aF�J�t�,������E\�lZ��7h��#��Ɓp���:��q���~Ўh�
.�_��ŏ%!��E����1�#�oӕ.Fe�O$�D���%��z�_��e;����z��w�f{'ޯ'�&�;�^p<<Ȉ��p�~�#��*��D�o����3��{[v�	,f=����sK�S)$�D��I��=���+JDE�	1��WW�/�V��0��*j�8��;��.Ԛ��'t�3]��ڪbY0�i�c&>���u��ɳ�mE8�+��������DY�)���<7���h MȺ��ub�`ד, �U�����	_�
��Jĥ�~��o�3�4| 
̜����"��H�Jjx�?ǘA�[��K����9��i�;oK��(~gq������?��GO�w�B���Kp�[;��|�SH�:݋h2�
+��N�����fT��ښ UA9�B���?�vl�S�Ը����`�^a��5M	i+��/6}zv����2:�-����t>o��U�7��H/8�h�a8G�W�?t]�� N����"��-F�V�+�O�m`�d|���������������h�[���s7�<�[�c0���gYĊ/�WBq0 �s?SQb�Q׃Q^k�W<�l�݄�gAJ �A�4��D�4�-Ք��4.Ղ��h)u���i0hw&�*a��B��̾��|�O�m�mr����1H13��|6}�P-�}:���&��뮑�Ll�����
�RO�j��rg ]
�.��":�E��-�@8�N#�4�~�т������սY��X0��ȃ-�M,�v�_қЀ�N��MX<���)��w������N߼ Y_!�C]��7�b�DC��Y��"u�ss:�9|ךN���!<�3�r����	�	X��g��U��Rq� ؚ�5�n�h������H��iV��x9�B�Z���ҒL�X��"gQˌ�S�����?�OU�C��|o��`�$��Бq1�^���E����?Ls3k�߶���H�b� l��N�?g�u�1��JBJ�H= yGv�?�{O��F^��d���3�r�5ԇ�H�4��c�?�4a�3s} ���Z��̒4�rX�8�̂�M��)������/23��A�=�3X�����J����;��S2�`�{�&QW�t2�Am%\�u�.��m�QL��4�I��)�wRV�����(s���r��dJ:�=pY���~��p�*�XӍP����r�Y���U=�c5]�
���8�^ʩ�S�OK�����R$�/r�ԟ��	R�h��a:�%������DI�7L�T< ��?��b�;��>��	3׀�-�R������P�}��C�!*VR	l93���SC�R	�Sc=�h:O�5Oq�!���`�l�^����64�{�'.l�bm4���.�ɖ���/^���!i�_��S�\� �p[
5�����q�va�b�F1��B�t�R��ըк�R�!�|9p������;��T�ԣ`A�e�#��(;���HF���1�����/T�ޔ�7���w@Ҡ�j�R�9�<Τm�a�y��\���I5�+��w0:�M�<4<yފ��eXV0C1 �V�|�ݜ����j >!�����Dp��{�":9p��M�o�a����y3��$�s�<�'�t��gF����~vDr8LA�g��L�ƞ$�|��78�}�=����,��||��ؐMh��G��۰=�벪���d$L�� +�3C9U,Y�~^�i�ae^[eov���pB��%R��F��[�d�՜zd��%��+�o�G�h�P���LN��4 ~׌bk�򑝒+�|���q� ���zc�G��cp�PK�X���#.�r�Tw��4��7�	���/>73��2bt����mW�f"Qˋ��T~��G����5�Íu[����@�S�K+֚(H�tٶu�p��;:°窢H$���h�s`Ik�w^��A R���M+>�!	��`�X��n7�)H1�{[��tWO�[����C�P�*��4]_��z����@��=�����'������k��@۴[�	��Y�_��KaWZ����B�
;_=��N,OT�����ӛ���fi��`D �����q��$%�6CI���Y�d�}GI)|�������%�P��������
R�(����}�Y��̻,�g4ؚ�����X�е�V;��;V�p>�Q$���x�����M�e>®��t����K�"�~�k:�1̐��,���ӧ��E�7�o[��.�;��6d^�ɭn�d�'�4ۊWv�)a��[�q�g���)*6w�}_b���4D�~/�.�0��I���[R�}U�Sv�(�����P�ZnZv�H�qXtM����h�'��.�/e�s���.	�3?E��H�`��#�M,fK5�R�-�R�^ֈl�vL�"p'[�I ���<�;��s>p�Io�}d*��B�R/F�gæ�щ=S�l*dJF]^o��J��Q)��u[�*�0�h71ebLA����f ?$ᛚ�)u�~�B?��M�Uܳ�)��M5��}�<��#�����J�9�����6Y"�ew�8�:S�Wm�/��+\�s�jl�x(�&�6ƞ;`��e�
Q;J>O�_��L�
(��?����8kI�
q}Q[DE1�=�8/J�R����܇��'����7�&���=|��-8I��8J���]���"��$�ho���3
��wa�� ��^������I�(�X�`�M��O�ãn墙�lNE���Y�kj13hl�th&�l��ǜ�C�w�#R��Hv==*��]��bs<y����>��R<�ޒ���SD,�����@�Cs.��5�h���X$�A�ݽ�R*�����*dn"���Yʮ�9�'���؄�������`��Sݰ����"�G�oyp��3TzC�CY`hm7�j�NʐgDw/l��F�8��aM����ߘ$�����i�9UυT{@.�k�o(��eę9WI��179�~Ɠ
�
|_O8)e���|�����þ���I�ui��9)�����l�Z �U*���ș﫠�/4]��rR��%��������G�6��NA�y����W�Hy���'��8�9�^��C���k�_�~m�^��\�ڒ!�çX.��(�?���(��	>�g��#�A�B�!U��k�z��'�-�̏h�:"���Vn�u�qȯȥdN�g"W�@k���I��Ο�9@jl;�i��2���7�x���k{��"�S� D��3~��������%�;��t%�w����s��u�������c�M�C)xt|{sr��Ο�.��*g�	�_���t�TB@Zٴ��	&���l9وLn�k��E�uh�C�-��/N����y�&n؞E5���փ�z�Yb���4�a+�`���n��P8!M��y�ڏ��ܗ�-���&w50���h̹�����b̳�})�T��op��t�*g󕌽X�Q��n�>"�����٬�sq�*�sG������b�Q���Z��z�2X��Ҹ�� �o�,@SRq���9��i��!�i�ؙ�10��\P62q�^�8"

��b��7,`,��c�EhL��+S��[��:�>?4��g[�k�U��ZKمC��9D�j�8�r��ܼP���/	�Hƃ�2 V7�Sly��־�aF���+����j�4�*����;��z���=?��H��� �j䌪�u�eiI��-���%�sR�IK�s3?i�ng�ݣܛP.��}��6��N9+?��,�V9���%B��)e0��w��%dl�f���T���T?�z\&�a���ʂ�H��SS����M�27�*��@V��t\�PH�][t���};�Q5�	�E@~x�� ��;̧�g�j^R"-�V㘦�ܟLN����\8Ŕ:A��nzU�`�J�_Ұ�(#l@�� s�r
������E2Z^oѧ��T�ܪ�A��Sex�ߵmH_7X�i���`�V=��@\X+�λqy�������� ψR,K!E՝N�B�b�vx��,#{1��Q��3,�J�6:�K.*�xq�ӝeX�;Q��/W�k�d�)�'H(-a'�ɠ�5��4�>+0IY�o{;P��lĉ�t3��m���	s���-�����`2��&7�ɩ�"8�i���c^p�e��* �2m4��K���Lsp�V.��V����{��`��+�
�P�#��O�rL*a[�.�@�O�ȩ��-�i㞃�`o^9��%�OB��h�&t�-�,��T�)*��B�4�*���B�{�쵎��n�.���{ܚgz�bn�:~B��	��D2�ǍL��a>�#L9z�'zAC��A����Oa)��w�@�������l��:�9;uA�!���U�t���q�@WZ�n��C�oE�e+�C���D�2f���I̱U� ݸ��ɳTKS�S0 wĔ�mQW�Ky(t"ȱ�Gn���:�jNmP��M;��N���kH��26���5D{
���@�f�-�D���v�=�%��[����(2)ȑ�D�E�����nd�܈k�lyr������6�h�o_�י����=zf
`t�ie?)�1$�gY%ԋ�|eˀ��	oNծ�#������uY����MyĬ]�hbKjə�A]�7?ڭ�^p�۹2�f�aU����H�\�����J���+#���]W�� d��ڊxeL���J�@Kq�[t~_�d�a���6�I��dT�JT덆����w�fPOB�����U	҃�6v]����r?�~�i�*s�熲>ҝ���2���D��G��2����A��{|%�Q�z�¦���f`|�鲦B>u�%މ/�5uz��ڍ�H^�}��cb��ܯ= h�׾/'<�U�9:���ku�B�	��[u� ��.)���M����R9y��|�V���B0DH9`���H�T-���d���&ki�?5q'���gZ�)9S^�9��g;Q��Y�8�18ޫŕ�5�ʢF��x�֛	��{B�,�bG�G0���.\c�i�-�&�����a��ǎ%s
!�ɫR�>>+���v_Q\�}U��~�ߊ~�+c���3KAL��/��,�p�r�� R��!�`j/����"Ib��9��G#G�be�v�[`��t~,�jW#�9d���-��0:ik���6��	���.��<&OVȗ2���4��l:
�W_C���;��B٣r�A�����C-�!�h8ݤ �}����)�a�1��Gg�h	ܡ��k��F=�gAA�o�Zw����=K�\����X3�t��Y�j]����g���wT�7��X�q���F\MO��C�O�M?�C��	Y[B!ZL{ɾ��6$��nwI|uwGZdfgڨ��fWZ����Wd�|�������y5�Q0O�����W M��x���>����M�u$��v��7$�T�U�JF����ߠ�L�,j�����R��j �	��	��B��Rim�N����ڠ��2��viVi.lf>L.�3:�u���@8C���c
��>��/�\��>ۙ	�P�</���{8�H�r���X�ֶ'՝���#�G�KӶg7(C�H��E�,Π���jK!.������r
�lv�=W�M����At;%��}۵��^�2y��m@6���� �s��"l���Γ���}/�7#	�	5؜m�xV��v��B�B��'΅~M3w��U\��ڋ(>	�Z�I1S�й�|���l�'swk��%��Z����+z_��6�"�ڔ��v}�-}��IO��$�Q_�����Q�H��5�sMfQC��1:��js���x���u�
.�GT���� B��_�}E�?��F���Y�4���ޜ��lt/1��v5>Y�L�I��*���Y��ijܾǴ4G+<U��1�z*��L��0>#cQ�b#�ؾ�d�o�b���]�ܫ�U�Ro�AzW�U�^U!�֗E�ˇ�69w��Z!ϝNq}0hZ0��N������e'�J���$����o��NɶN+�E�ɻzHw�'��?t@�4�f,u~�[Gm�K@��ƽ�0ڒ)��^v���Z�YS�-��xO�/��:?>A��~z�Z�c��y"K���V��ȖUyW]��Z�
�N%w�9�=�����?��п��i^m�����e7��R��ŭ���*%3>;��\�;x���)q�%{��{� Y�<6$EQ=���Ck?�ho=d]?v�IF���Ɯݸ��ٱ�s����	�2 �����x/v��laJOB㎀�_�sU񚽪Pk�2��c
䡻9�b����^��I����<p�!u�n
Z�tm�Zx�k����%�����
���Y[�Ψ��L3����d(~� � |�|U�|^@�?�x�W�b�q���|~��m\_�ᆶ�����55�#,�P;mrg�ՌrB&ڍˉa�y���m�t�+�1m���$�Z~�0%$wN��~Z����«��$����\绖�4 �l� ���g�A������br�S
�6|��#���qN *E�"�I's��?ޝ�V�)H5-
W����'V�h 'N���r
}jl�F�ݽ}�7��d�c�	ro���bÂw�I���I���b;=i�*0�2*�M��`5Pk9��2�<8���$7����� �֯�,�3����P�z��o�d�s�
�;�Q��6����z�]1��i�$�QM�o~�>,�^Q��/D����X�:	AK��Q֦���#�e�} ���&o��#�v���FEx�~����o�S���VyY���w{��w�O�]y�X�ϸ;[���_�@�6@�=:yH hL~AQ��(�����뚒��+���:a�UGzZ�gE�0&ɪl6�#)�l��g�E ��/�/U$��s>[ �4�[S�CY�r�a�V.�U�	h�C����\�R�r���؃*e[�@V����|D��F?4J�j�H��5�����j��l������{f�~n�+�e�޶R�Q�k_�#��옾��y1Sdێ�Ba����عc�lC�y⟬P_����B[�&[�\[��vt Fij�'$?N
NN@@�q��|���f�w!TV��Q7�Ν��ٵJ�����W7��%S�h���*������[���ǹn�T��=���~���0�y����:�B���'�U {����!* ���.&��a`-M���K�Y��znY2�{4�Op��mt��;1�괻��OO��&f>�*/���[��i�'��;X;c1f��g,5r�B���A6i(4���3U�s�,6����S�?T�i|�u�T��(� �x�Q��=�Ys>Z�7	&=�D��|��S0�g�PFy���q�ޘ��L�(a�e6������4�H��B#.d��f�'3���%�9�P����v�A��c�2��Z�"5�2���C�iIX����x߫�5���xӀ�)��qc zM�E�W�����R��2�%�x~e:Yg?�}ljs�����*�/��hm���G1�3��/��`R#���Ƀ-IC�RL��z��$��	�S���$a֣K��=�a���t�a��pS)��w�׶�XM,Ə�VASM���/�J�*w��ՓF�ĕ[�G	D�� hyX}G�Q�)9L̇o����A�E���5r^X��0�Y>���R�ɂW�q7¥���6;�J���x�"��l=�����z�U_�m#�*��'�O������0���9�%�+�~�O��m")<th��ۥ��ؓ�iJe�邁ӛ�]�h���E&�_�(��Mm?ȕ�Jm!W�y�p�A���2�j�m�H�;������}"#�O�P5) ��w�9l�
zD�?\#X
cy[YB�+�����ܼL6�u�H��f �o��{z�i�Y_"�-$J���e����S�f�@D �c������WG˴����04j��`3ⶎ8Yk)����f5�S�N2Ej�>B�0��1������3�쯔w*5�!�B�rIc�gg��W�1�5B���̃�Ӑ�Z��.Xf�X7R�V��o'P7���Td�5�y~oǢln��řp:�H!���
���E�*�I@ʷ<���X�^�=cDa Av�]rB�W���\�<�f��r��i�޹�NPɩL�э�<�����uIw4w3#�=��J��{�(�h��"[^��[T6z�5~~_o�`��h_IF���,Z(�yb��Lf&���o��Qn��^��g���I����;"�=ſ��&���n)��d�]ӄ��޸���]��5i&�-�ÒQa�	҉+J��ީ�DeW���E�w�ӌ������"�
�1�|�m�P�L˪aJ���2s�7F���)L�Z�9b9S�=
-�ΏcE��8T�ٽ:�#���ԕRT	xY����5����۵���v�����w{�?�(��h����f3��t�4x���f��0���zr]u�������r�$���a�	W���w��W�%�mne�#�f�1B��q6�;��1�A��
�_1����8Ĵ�_K[���c��`�Q�<0%\
�����Z�7�)GLamڥ��^@�}��.w������p�xk��\��֨v���ѵ�Ȝ�yW�E�W�9��^1%1�X�3����mk2�� `צv��K�ƞT���N�߱Ԟ%��A�Rq��*�9~�-p9�W�f�Pa7�{T/���b��@ӗ�.򔋂]�Q�U�
�/����F��#�
�I���GzHyX��c��:������<�SN�Z틶:��03�㺸@�R��-O�~�����T�%�ʃ��yj7�,�.�����y��h��Xx���@�W]��o�D�̿T�tL#eӼ�4E��T���)��S�,�\�����Xz��yҜ1K����W�%5@��*:�N�0��]&�M0)#�~L���-�-�Z�2�����v���Eg����2Zi:?�z1�6����sz�SHW��<�>�����h��-x�+z���D���oO(SZ
KlŐ��T$ɠ�)���V3絠nڿ`ҤO�<)"�j�yeȪ�J���rd����څjoz?ϒG"��&� ��.	rI�E��{6|�J�n���;�kY���۠r)�"~���q�3��N�̤����H���0�-i�pDl����(���1?3�0x\k�*��{D-t���ͥU*kU5_�;�-~{�J�$[@W���{弳���s�����eV��eg�z�G��7+�q�=;.�_ ����Y�`x' ?|�nr���W����g06z,�C*�:(��87��C�^�PrX�1�!��
��D�#��=x�Ώ��ĩ����N�>̟��9+�(�CC�f�h»�RE��l�0lk�$'8�R��2 �i/�m��54��%;����cnd��Dl��|:�	�rHW�j-HX]x�^t�bpl��@ 9�Kz[_uuȜ�$gB���������l5�#ħ!įO�Q����X����0��!	,�`t`�f�[7�?���� �|�����w�~��!f�#�wGn��d��a?� ���^J��18��ʒ�O�d����1,�%�X%�~s�$ A�0?�3�ຼ��0O�e�fo>�§�i6��H���Al�K�㼡@��t�F�����	�.K����{gU�" "�/�|��1�ă_F�2"��y0yjp�иLg��ȷ�d�Ou@q4v�����Rԅ�7��%^aT߫x���a|6f�)=��j�=�h%
��@C�˨s�����܎7&��h,R 3��@Oz�J�H�Y����%����u���˝+�_O����\��������ͯ��h3�OXS	/�\Y��U���������Z��O6�ˡ�,�.]l�t�m�@��L���o�@-�q`7��T}#<�L�]Tۤ��i��H;�H��A��Yi5��~7h<�f!fc�ӂ�"2cp���$���>����V�jy�bhyK�pM�B`V�p�Gn*�gv~���Tm���LϺ��F}��X��q������|/Z_YL���?F"#�i��V������$�B؄��;�L� U6k��UnE�CVHUd�?�4�pؕ-\s�2ؘe�^�a��f��ʒCؤ��9�H��⻙��lro���{��:J|N����$���*���'lzlg=�x��&}O��H{�ޭ�]�d��������2�i/�X��5�v���j��]��I�{IS37og�T���[��\iO^�s�xn*�J�7�n�����34˘cW�f�P�W�N���m'�(J��	}�}j.�M�]MHo��V�&튈Qf�5v�D}� t���xh݁�p��d����z|,j�{�|����m����Lzy�ˑ��E���P�޳������_3?����[*E㌘͍���7-uIu����mӥ�����Ko7^h/�� �)��Ep!5(y1���o���:IQ�N��$�?�nƸ������!�#�yY~�V"�w�����1�����_��L�x"��V��'~:��q�6T���!�-	3W�r�.2h,efT,�:U��ʳ��n��k�&6	{B��ן®iS�V�!���m�ޔ��ϣUE��h���hC���5h��m6;F��|�j�d�����\�ۅ*���ev���+��*A,�BJj�m�{e���B�Z E哃?ӹ�%ڶ������:K��\�z%~67�Q&gl{��m��Q��F�������d�2���_w���p~4y2cJa""�Du1�؜p�,��p��d�� �1�#�:&�F�7���4:��o�e5�� �"8�Cg|�D����l֥v�r��*���}R�rɯDJ�hGD��I�}��!Px��R�rM�j-�Y�>Ǆ�;%oX�ݟ �(����5�����9&o�e�	Cj��q. ���O������![Ǖ\�R%�!��v�dߞ��@
��=8�V�}]�ť�K��*G[Z��k6?r�����2��P�'�� �R�g�^S/�Ӣ��o>K���~ߛPZ��kS��d��|`��L\==o���
���+C��
"���C^�Ƃ[f��&aa�/�MBU�:�ջ��*n	� �&�jV��?LFb��R��怨#�;gM)�,��\쟋�~'�f��|��͚���s=�H�\��!1�/���W��1����>Ɖg����_c	Da��#*���܊gZ�U81��	Ļ�ߟ��n�顴��8��(�?�Uo�9�AT1'�膌��r/+}W��U�����	v�����E׻_�zYʱ�n�W���.g}^4��O�f�= ���݄AII����*��������%@L��6��W�������h/���x��=�n��2˯��i�K��P��B̰*�zہ��@�v`G���ѣ�&p�5�ד���1����苑����ɩ �^�k���Dz(����fb�o���@>�S���z8��D��%��.6�p�N��½�Թ)@>�n=����B�nW�rc>ũ�5G��6�l��l�|a��c��߁�~ T��o�S+�U��_'U��HV���:@��-I�EZ�&���.���j�)bA?����˧<"E(8�v�ܧ���?.R:�v/JN�^m�Z!X�V$��@��
�,=:�m�y�'4.[ع�ԘpNgR�h�{p�����Y�j�u��7��#a��h��A��E�ǭw�r�h��p<�b�X��dW���w5���f%��ݍ��ֹ���̫����V@)u|��g��� sM)� �Q�4�S�M2k������j��hF�������88� .��j����D��XS'�そ�W�D��.���)�9w�i�4�q�5��<9�S1���xE�9��?J���Ei��ϭ2ʺ��I�EL���z'��x(���1j�EL�ӅE�7�9\�2��ib�I+����`��/�/��9�2\.���[m(���e��<�ظ��k�D�i���t*_�����B4�s��7�f�u��`d���2K����P�.b�|ai9�6���>�D���@�w]��pZ�G�1e�n���"����j7U؏�	������)�Y{7YA91�l��Mz��n��3��x�.��i��n�� %8�<�������\�6�����?�#﷖��G�#��ΖLq��P@!Yg���H��MK�e�+�h`mT>+���y���A��*���Ⅳ��<1Uc������b�Rˀ���Ȇ�6tqP�G��u�?NYyf�q�++U �~��v+8���_^��B���;[�<R���U�A<�
[�N�˖?�B��}�T���vRr�(:s��A�L�]��(���w��!��C`��Z[=��{~_�ӎ9l��H1K	��TعA��KE����ںh(W8e�zų���`$��n^�䘛�3<����{��Z�G��6r������FH:V�(af�s>�}A`-��YQOz8=�Lή���1��W��;�r��u�C\�2�/�Һp*��r%ˍ]��n�������c��a�!L��M5p�K8��9+ ,^�'I�Kn�d�E�I���i������մ�y�C��B�_�������C��C�����ʷ�ƻ�Q8v���5H���Z�R3����H����;~�.!�*��]͈�L�OqC��YjFd��K+J�Tf��b��͆� �؄Y�:\�`��xr`��H���f����M���n@�+�ml�N
�y�ku�b}�<W� �EԀT���(R�Ύ���,�
�^m�!}��[�YKT�n���S�d�h�.��i)lxj��^ج´�~�C	��=<B�L8�ڌ�J�PG�	vN�L�I�����;FbD�i�hUA1�ʦ/;x�$�ڰ���k2���$����y��"�g��/ḿר ����ts���`D0h<*�(?����`�6�S�*He�r��b� �_A�=������O-�
a"��jXL��gW ҩ%oCχ��wc���V-Io�K�c�~�o�%R*]�OGt���zл��d4G�^���yUvS�e��xh��Z	�B�l� sT�s���a�� ��Hj��c�P϶�},��L� �:+b�Mp�:�-�Ф��N������K[�m�B��_��\<�[��XۃƝm���&Y�W\bq�?Qe/ݱ��t`bH10ٲ�����,q����Jb��X�%B�*���	BpW�-�S�E6�Z�7�*J8�W�rM��t����,eJ{�qa�N��)J��!w����r�.�]����Em��o��,����n[��� �=ߘU�0�Q���f��m'җ	��ZLd�!<H~<��q���L�0%��g�j�?�{{������Ct/��))�Xb�j��lA�2�1��N�SI�G� WY����Pa5>'�g���:i���{I���|.� �oO@�l�D��'<@R�Q3d(�y�uo�T�Q%H�p��S6ti�t�8���@�	f�+���'M�FB����edp��#Z�R��@o]�;�bBN(��O&�zD_�br;���5n��AQ>��4o��oL�7�Y������B��00㻦<>:J�X��{ȶC��/tj���ت�f��w��S,��眤Bܙ(�u�[n��q��$���Y�=Gd�JZ�0�����}4�O� f�ML��@Ʈ��И�gK���J+p����KQ�)�x�B+�-��*�l#��٠�vV����a��il���(�8���s,爐fX9��0ߨ�L��z�_�@����7�<�9��]b'&�%�qQ���ΩȎG]�cj����,�e9�<X�^HX�Rz�uP��-��k��6�[�=Dvu���"�;p���9��5ܑL�!�N_)s��3�^���cg��_��/��g�;��aB�����+��_�3vA��"&b[�"�V�弁)ѡ�2��%q˞{�
��N�|r1�(n<�-����vWh\��9	i�60Ž��dvXF�� {R��z4U�������Sy����e@�j��`T�>}5\�|�G�)�W�ۙ��Pyc��h������(#eX%kE��]u&�Y,��������XV��_���t>�qsD�iF~����ˊ�##J��k��[�M.l��@��!��u��
�8�gFD�Qe�׼w眞a��1��K���2�̰���h"pNR��������$}J׹��Yv�~��m�Q������-�뗜d��8P���[?y5 \~��� ���<��h�I����oм���8y�\_vy�D�K�9A���#2��۱�Azb�KD1l��Ǣv�.�8p�{�΋/�I6�Y�٘�Bq%�D��f�$-���X������HO]q��u��?��	�Q���T��m�jm�2x�@8x|?(t��L�:�3�ޡ��=J����Br��(�Pp���)�i��$�Р�l���@+K�z�zk���j"�I��Ok��Ƒ��0�chr ^ ��bt��-��f�N�1��p��٦�6��Vܵ��b�{�Z*�H�2�|~���ʾ�+`/+��wy#j��c���#�"���`UC��!���V96>�����c��BP{e�dU��D�C
d6�Ga���ۄ�����[IJɲ ���v������x}�?�U?�n���$�Pt��C�F-(Ѣ�Eoэ�A�3G4��m��,L#����`d*��K�>y"�EoX��O�r�AE)��-�,� @&
�Ū ��\�K�m3-gm"��	�a��.�A�8[�S�H��i��l%�b���z�T����e�7�L@lx�'�|l��)K����n�Л�E����y��Q�~-�,��R/5FqIi�P:XO������D4�g�6Ḧ́�x�����f,�^Ge%����%���(����s�I���1)����h3>���p��f鄇���c���f���,M�eŊ�]�7��jI6H�sn�`h.�,eMMc���1��1����Y{I�G*7�� ����Л��H���9����*�prOZ�o{��n�AS��fyo.�*��n��Tx���6�!zcH&8�yؒ4�6o���ߧ�����8���/na�p�->b�-Z�_e�m�s��9����Cv�=��r���0P�����P����6,ދ�Rދ�hf�{d0��� J���guE�l�
���Rp7�.�����fSd�u+�8d����bi���ލǁ*gw��/5�$@�͢����k9����ʡ
'��� �T��M�q�I��6X�L�Ҟ�G���G�']r���0��v*�Օ�ck�HbV��Lv9g�o	�2��B�X�-D��' ���y�sRh|y�=tt�ߪ�D��XCu|P�4����I_nY�E:t�8AM�Uz�n҆�>샥C<1����%{��sV�i;�����`��e��9��.�9���2C�E��S�5�Ҕ�o�R���I��Y��^%U�}Yޯ�z͚�8�V��=�ΑFN�����(�t��L�]Ww��sJ��;���n*����F�R���D)$�kX�[�j�@+���'F|�fN���M����S�����G�gX���5��n���RQÝ�s����FcB���D�T1����MC��Ʒ��X�G�� ��R�``�j�C�uh�NJH��S?�,�>�`-����%�ENl�ά�i����/���q���E�HT����8�r�Ӛ��#?kj��_:)̧s4���5�\��^��f���H-4Q4��2!��D���唟5 �	SB��T��:S5U[��ˑ2����,`�&�;7�|n0�#�%�y`�n"��/z�OX\�Z�Ik���z%{����vd����Mm��8�7��N0��2�͟�J-�=˪��h���2^4о��I���+*R��g�.�v#��&�3B0��7M70�3��c���oQY�����.ў��CR����otJu�#�\�����Sn�6Q��Ӑ7�(-8��+��|	��-P*o��2n�(�\NJԂ��fc~&f�G�I��^ə���'�-.��ƺ	�i3��B-$5��8o��Zi//Rh�%��p��?ֹdЋ��2|h�	�^ډX�O}��C_���A�C�?��G�֞��]|�@�w�k�h��q��l�����t ��uX��Q;Ϳ3���ٌ�H#������KM9�g3�y�|���f�V"ALZT�X@d(�MK����ʌ��s���خ̈́�P��k'C��؂�e\�ܖ�_��6Q�y ��L�&#�b`��6� 
�R���7���.�g�(t�tEC���&gBH��Q��E��G���J���,7I6�y�ٟs�1C�Q�T��[�_cw�=�k/e����42:IT���׀(0#2�k��M�i���ɖQ�Kye���i�Y�V�<�cCB��J��q��Y�5��tv�E��'\tq�C1ڴ�q6֮��'kܚ]�rK�N��t��硥���ꕂP���)j	��FzV!�ti7�ne����o�g1���b8ᓿ��8��}m�/p�%��uSeb}���
C(v��o��c�g[p�کs�8blv�y~J�{�I�@��hΦ�3��@�S��;��N�uE�

�u�3�I�W��pȅ��,����xy�n�Φ�ka^�g�L���L!>����ٔ��+q]R@T�Q�qPV��ŀ1�)�I��h��|iM�	.v�l�����Ԃƚ���+x�3# o�r�qI����F~��*Y�C2�l:_X:2]�����m���ۛ��^G2��`2�|��[�'�կ7SyKN��g����Z�r��.Qy�HRϝ���qt��%��Ou�5�_l!�^sm�6�Q{��B8F��q8t���T�F�#�.�P�~�� -��o��.��xLkFS\���Ɗ�����"����.��.�w�b"/��� ��:z����؂�F�Z6P�'b�yQ����I��GC*�aײ|����%��Y.l&���H��EE�"��2�d�����|7DD�2@�� ���x���05j6Kc�ֻJ1Z��q�8N}��8d��.�|��9=�Sd��]Q/�s�`	=��b���(�r�%\!w��$�=�S]��/=%�|��\�� ��G���9b3J�v(N��pJ��������X ���n��d
�q��/5�pZ�BK��f1ǆ1J�7R��7��H$M�c�X&iň:���g�a>�H�/��ۃ�ﳼY:�2ӱ�6q�M��%�ɨg��r^�z�?}�7���Jt�ŹQ���~��C!���q�.����;uP)וs�t��+'����tgߐa�i�w:�{Y��&�����C��P���l4�l�nc6�-FsC�Q��+O��d���q�6�@��KOU�Y�5=�4�)��:%:L>�]c��}�J����l��4;�+]��H}W%jIɍV��a*��mߑ�S=h�\�9��S��E��5�i����K%���� �ꕑI� "ѿ�#��u݈��}P��]y�N�������5g��7o+�4�`���O�wPi��:q�N �*n0�C��`H������՗�thP���^e)Q�Ų���ը�W� :=#�]��x>d���"��>��!��Di��$���W��z�e�x��<�8�������� �\��۹������VL)llv& 
�����E5�Y<j�;Y0Ѫ���X��"���Wc9<�_Fϰ�����8\C�������kn����6"��z�L�Y�~*ό�o�U�1��I��Z�_s�����O<����W�D�;|�m�o>w���=�v2�S?�#�/])Q-fZ.��&7+'�a��|��M�Р�d�N���$;����� ��Et����!f�\�J-��y�OG2��SYY}�q &(��#�r�|���'���ڇ�0ܴ��Pr8��=���KO�<��C^����k��������7���[$y���B�C
6��3�M����1@����I[�)H>��$a��eH�s����7�-�b6�h�����}O��C񽉞�Q>fe^v,z�!��}N��5��E���������O��V��3{O� �(����1l���5'aY��{�*f�4��$�>�\�R��)B?Jx�g�oo#��cB�y��U��6I}彔�8�������I:��}6,D��\n��E�K(VXe�Y�N!P����/�̓�t7����_��m�m��~C	�� @M]�:�Ʃ5! �R��C-���<mO6�U�mY��&��Ej�#Y��o��X��Y�2B�rn	M� p�0g��1�ϔ�����6@�=8�_��,�u�qZf�A���^���(�%�����%q�j�Z?�%-�>��D��sF-���y;�]a�˄a�@�U�6��德o޿��e�ȍ����ܹw��!Qc��/�	H}T=�����N���x�1raڌn�7B,8���	�j��py�VY�]���ot2�Fʸ�v�<�Q�h-����
f֒���@:��O��\�2v�련v�X��s ����=1@����.�jp��JۤzlC���J��p�� �[���;�y9�UV�+�y<���#;i�y���.�q����5��ۮ�� �dlY����ی�,�M�)�bh���U��c��X����Cm_�q--һ��
��݂F�:T�vt�H� /_v	�ǋ�a�rb�i�c�g�7�2#A���`-KMx#9y�D�,(T�>�Z�f��a|��R�?J��B[�B��^���P�H�C�A3s����{�O��c�(b��`Z�_��U7¢>���J3��`��>�F�2��۹Tl<�������Ҡ�\Q�*=�L�Yx�`��]}%� �v.#��.U ul��KR?N+Il �+5~��`x+���h���k$
��{6����k�2����,�V3F�.|��?� �x���AQ�!/���?�#]�.#�Tg�דr����Oi��
���R|��Q���%�c���jFI�=�Nx֠|y���W�D�#z��+8�a7:��g9�gЅ]�W��v��A5� �Zub�PL�*9H<3Ix��l������&�|�o�/�+��;6r4N�A]����C9�5���Γ;U�e(y2 K�QΥ�h��6�'Ω�/�*q��c��}�u�R�p[��a�����\Ǵ�[^8�0HD���&�Y2��5�
�`��/x/�LҾˋ���F�)�A����J���)a��ںwG�l��_��C�N������P�w�� �tI��OA����Ժ���෽�.Hu[���5u)�P�a����$y���E =�_Lm�ԧ6.��r<��!�Y��y߆�g:�K!}��w���l]]հ���{_������F!Jb*�ɳ��Ch\��o��`��ڝ��pk�ט��udх��.�n���L��Lޡ?��ϵE�Ѳo羓��8v|�}�8z���C��vN�]��gaX�����c{\S�r�B���}�
(_�3�� �0���J;;����vRu�Ao�5����G�����-6C��5&�B5�)�����]���U��%b
��ыUڀ�W�!����^�o����(�[�m���fp���mgx&���|�gomT��n봢Y�]��,�pz�3vwKQ�d�lIcP���͢�S2�_lY:��Q��*���}�=�*mB���k
��-��89ΞC�"�{�jH�Y���e��vZ*�����/b�k�Bo9���c���f�4��MLƶS��_�=���U�D�� o�.�F�Ǻ��D��QL����$�%���I��h3�F;օ�Kw\���ݡ�}E.��4�S��+�X��\G�O��z��.:��v�$*v^�t&�r�'Ǐ�dȪ?\����@��Eg0��4R Q.�x�lf�e�jK����H���P#�{83���2���ͅ��~&�P�C�坽�П{{Q�޳�9�HQ!�D�haW���o�^�ں��i��s�Q��.�Y���a���-��z�X�}��2�1_����Gg8�ՙ�t#,{�8�;����W�����M)�t����Ӿq��bS�Y?h,�Zk`�{*��c�Y�����G[]���vM��œ�gf�.�}w�7����&TZ`2r(�� ����ｗJ�M`�@��կ�ũQ�v}p����[f�:
��{:9~��ԅ�CP��q�t(^�Q2&]��3?j�����5����ڨ�S((gȐ�}�V�#�1�:.��8�զ�*Ы(��b��-͟�����O@R=�鲚���CrDҼ.e�H��@�y��� :QXn����u�ĩ}����L)^�1�,���6]x��W1b`�_�M����h�'�����e���bf>�*wY@����D���O����t*��W�A��ڨ_���	햧{#=��[0V���%#���ra�a�^�q\���+���6���_勘~��m��i5߂h�L,ԙ�2d����坑(&�k�4@�N��D
츿4)�߀Н��L���Fw�}.���<�����-+�c跡]z� ?r�����8j5ݖD���컛��Ӓ��p�ȸ��	
J)s�)�ˋԏ�94ʺ���E�,���[=���s��a��6jǷ�O~3���?X(W����p$�^�a4g-B
��a���;��*�K������-�	m>Aal�l��:P5��1\�;�Fu�ͅ���=PS��z{�	���?�� eK���4f6���1�.e��p�?��늱%�f;{�y��u.������<�5�<?�|�n��I�����X˟.��٬��R�S��|�"��P���H�Z(d�~%1�����}�8ZI�������na���K����)�}�{�4ϭ�DX��z��2�7��}O9xj��T�_낦Hh߶j3�WO\z@����E���Ɛ���|l͹`vB:�?�"~^�,xJ��-8F5�,�}uo��~���S���Z��7���u�Wv%k�s���c�n�E�|}�5��q����߸��%�)�/G�t�C��͔7��""�OxZ�sr�b�ՄR���N�4�ͿTJ�R���Ő�sK�UEog�?tq��w65��h�tx]>}�c��"��3�N����r�:���,�P/���Ų�jB��/>�6hsj~e;�L͠>}~oal�]*�n������w���fǸ˟���K�V�L�\��z�����&3F���}B�:��ڵ�^�X�|��Z�E���`�u�ԗ���,f,�k҂�V�A����C�~)ۉ��V�(ɿ�b�Ӯ�����ng�a[(;��<��,B�3�xy�wp�Ǹ]����BA�.x!k�ڥG��W��au<)&��XC`��XC~N�i?��L3��a��!��I�邖��,��`���5�]u&���з>���f�*����g����cǆ��h��R)R��0���W��W	�XW�Ĩ����=d�b�\P)��r��� V�S�V
��v8,��_)L���q%�Fy��9��k.�J�,�u�[O��؆K/֧�$���}�?%����v�'��LE�\9��<���y�g�\G9��]�Z�V�K��-����#�6JGRk� ��N�l�55��Zq�֤Ƹ�⠰�_K�"��� ���������
�Ƣ��V�x�H`5u�dѐ�g��7U]�m����;�).����5�e�nr�3��Z��Ч�~n�R�ݎ��N���V�d4��p��$��Q�]��Y�^ .�ϙ
I�F��KS�������%��gf�_�lW���F���m9e��u�g�`�o�X,؋XO�/�I�>�\��� 5 ��}�;�|��E~������?}e��iS}�p��,"l)Pph�v�;9�O��6�߱�2�r�鸴H��a�w��74C;���"gϑ7�D�>/���t}�� Vӯ$I�d\p$�ȥX;�F�C�Sw\���0����B]���ΤB���Z־\���WB��r(Οy,�R�������Mt����Q�[$\����y7�ފ�f�%�."�ē��&K����e}&
�Σj�J��!C�O���C��}P%}�c)z!�:x3���7qf5��g����0����ǟ��&��FӦ�WMz��3O#�Z� ]�͒B�R��)�KI�����B����U> �Ѹ�o���\�6J,d��E��'I��Ĵ[v\�� o��v��%���F~;eY��zso^�Ͽ�W	ۼ�A�4��m"��y�Ņt2	�XT�5{�ޙU����C�-�G�j�8[�IuA�<\wV�p�\��cբ���؋���G�\]}��W�v�w���Z�
`��٫SfG?�K<��Q�]H���3IIj���}M�#���dTv�����f��z-�7Q%H�֐�z�-�|�;1F�[�M4}'�A���1A[��!�)?�f�<�	ѿ��궘�`/%�EV��(�����39��pod���uCQc�0�b'�W�����w��Y[���=�|Bt#���K`>���=���X�ฌ�k��K�'����2.ǹ����N�I�x�%d:��yB5��&@&'����aJ����ؠ̅8�+�p}-,ZFsV��`�'%������G�ѐw��4�C��d��d`��&
���U��s4%�u$}��V�Wv,�^����`�S�Pv�?�Gs ����1X�Q�!x�# D[��S���Q���M��ݱx��6c�s�
����tD��&�%Ϲs'npt�6���=��&m��ŧ�n)i� V� <،JFt$k5���	�1=3���(�-䚳�kt?�@��B�Y�b����5�r��	2�k��-> ��%����slfv�����e�aÂ��5�Gf�P�G`�h qP?� �Ѭ�h�� <��A�g�E������:
���:8�پ](�L��bM����Ao�������!+o��+e&߯ŧg�z`�$_,=_JӺ��G+���c����Ը�K5���+j��{d�sYky/W	��M��"P��B�@�R��	���ԯ��<y >st��0	��ճ�Ӫr��%r�e�!Ĥ�p��	r�q���>��M���uN$��e��G� �"�S�H��9�\q�1��o����|�-�"�{���B��c�n 0�G]�*F��:���n��L���`���N3����
son�}�]8�=@�Ky�4���U7	�^sev����y��ܼ)�>��O|�慎O_��
�g�jPv�	َ0O?�T*սt�؂��{��|̧�����S��eTRu!9��
�Ġ�����
���X/�6��o�h�T@
EN�
��
�H��\UM�S�sC:h�-|ܫ��p�\��M�������3�F:A��VDm�W[�0K�8���Oz�[{oe���3�tUp�#T`c)��-½̋e#{TQk�:3�����~���CO#�D�v�-�B"���k*/���cL؁8��doFk��(&oK��Mʋ�Y�~!�������[�_����P�/H,?,9���*q�
���Z�g` ���T�8/��b"+�ܷhn~XO,!�/�#g��#�xfYf�j��� �%�x��Sv���L
�9�To�&�� 3�,��[r�����T�m�8 /E�k�W�u���.�g.��~���"����w+�;��EK��~�&�;e_�b#e' �H�%��
���9lԱ��{������kC��J<�G�� lp��,a�:&>m��_[g����rf��-�]]�g�A�燙m-�:>�eqo3������X}ċӦ%����c�
Z��@��o�jf����;��t��˅�_TӦ WҋlӃ���ÎK	�!�P5V�,�N9x��\�Uo�����7��T�E�sDp��H��7�wL�/��Z�0#g︙y�0����o��(�v����q�b���������	ӗK�k.�� �S��A,�fՒ����諪fd?��y�&���/Xxy.%�;7T	��q���p��ym�ߔ�|��f���|�C�����n�EV
�-^&��f��Dijɛbx�ܪ�p�d��Fg�o��^L�mG�"�'n�ܬ�UٝT޽���t���<FP&�Б�Θ� k �%����;2�D@%~�F�IӰ��s�q�2.��gv;r6���,���ƚA���d
�@�<�� �Q�zW�e���S�#��۾��ap��`i�|E���
}Cs����ޱ]�����p��Vȣ�	���s@���nI�����ma�~��������L�	th�~^��G?��"sǬ���%�0�C�C߱`��*K�GͲ���Q�LB��zo�^�Q��[�#_�"Y�k�`��u�E$���D��!��r9��\8�[ؑ+���6�Z�֚_�Hz�_�Z�O^��,p��Y�%��Tq�Oݾ� ���#?�r\A���57}	�����"e���榙IX�x�`v�Rp(8�x���j����離v70Cq8;z�I�a!��ަ-�cq���d�u�k�#u8��6�i����������v���	T�^����-��� t{���]rTt@���6w˱߇�wHi����Q�u˫ë�#�HP�`��Y�N0�j����Y�0qčV!i��W�!"8ݽ��	�؎rE������B�H��O�g&^͏��8#���n�K`�V\f�L�i�a\C�Vd�-P�4}��T�\�5�x�J��+�𶿺���l��f�cB�!-v��[��7ʜ���K�Ə����$��|����y�������ح���oS��	�x��(B�{�/dmku��a�B)<�� ���hbr�v�Y�u��,����5VϹƪz,ӑ=+?"��y�;s�^�-�&��;�(�.T�[;�|H��)D�(0�;bYށ
v�&�5~?ɟ�|����&J�;A?�d�Ix�����\ld�0j�Y��_rK�\����[�\5T%��vRT���xc�%i�i�e'�$LY�4?�.���r�DX�b|(Ӝ#_��	��0U��^.A3Q$���sC�Z��c�������D5p�K��q��;�
nȐ�\�B).HN�ȣ���E�8!�ή��)���v.δ9:��"q��|�X�嘼3�e:"b�[PY8���p'�iPR�c}NI��de��W:�*��al'=�!�n����:�"��B�S������]�3�J�Jp��IX)h_oL cA�,(;��@�kD'��O��,(m�A�A��q���~h��p��p���,ꩋ�Ͻ|h8�M3�0&�2�{�xߩ5F��ß+Oc��EK��F�z$JNY�;s*\#�����G���Srn�Z]���T����<? �&7�J`�oY�V�"dW�� �����:�`��[^�8��e���-���1��ף���&��Vr=bRPd�Ib���Sk�x�I��ܑ<0'�U��;�?^g�����q��MR�v�����0;�݉R&
�gp@�^�˛�*���R�gG�d:��Н�N�"�	�}?���
L��v%�Č7���d��P��5,����mۻ{��� �R*�,���W�ᲊk��5���#���r�m�M���f��t}�������@�9� �i����XGV���)� p~�6
���2&������]LG|qC50H�W�@��k���+H��K����~��2u!;���~3ͬa�L:���-m�5)ӂ3��Xo�ѷ���V���ʎU��P�8�WxoQë>���S{���jX�]6؈��R�W��!�QZ�a-���>��������ϭY����<�K��P2�/�������;�JX��~	Fj���
�5-'�8k�{XNK�mĶni@�G�\أ`�A���l�j��0y!	�����鳝Q���ib<8�݋��J�`m��r|��/��0����Ԅ�?A��#b��%b��_P�am�*�u���b}��ȩlR�E?�\�3pM�(9{�ߚv��`��g�थ��㓺C�$^���s���f�0Fi���j���,:/y<��ͱ��o_������_|72��!�'� H?����3��X�k�Y�:�)���4�yƧ���C\��v�9�)q�?H�b�@�j�<���㥡!���Ϙ��-�as&�ʯ=?Q�Lᬦ��ds��O7^��eu�����+�W �fO��V-���ф�@=)r�E0>�O�@�=6�E[ ��[Z_.���a�,i*���mm�����$ Ƕm�g�Uޠd+t�<�[_+��ymy�=?P7o�2��זf�s�28����<��SO9��d�p�c�n��=<6s�A'Uќ�?�X���o��"�}��E�������G���t�}�P(����|63/�	���o���E�f�KU���<P��c��f������Ρ#9M5Vؓ���zo��Po��P���w�7'��7A�|̯�1���6iM{^9�-\C��̚C���k.�	��0!�t|���Y*<��t������/)4J���g}��9��9'	�U;�Y��C�L� ڕ���jZ,�μ���1ʎ}LGBͷ:��j����|l��w\��,�P&����s��~��T��k'����y�Уd�Ÿ�L%�y��I�1q�u�@s'Î�`U����w~	�{ZH_���N�Sj�֕�K�؃úKl�$xU��--
��'*�����<�\m�� ;k�� ,��%�D?Ͼ* U�Dǖ��?��k\���1��"	S��űfe�ዬ&<�U�A4׸���.��<HO_mۣ�%�9f��X�U��|".B�uZ��:D��[���h%"b�8�}����=�SA���K����-dz�_�Z��E�ʴ�Mྥt-��MpN�
�v����~��	�
V�"�&W\3��TG�ڕ\��VZ�a1��lM{#Lz�� )Ե�ʻ�
�|��&��5e�:�s�_�;��+�>�R��@���A��n�M�!.i���h�4��%��㕛evi�\e�:~�\���E�E�"4ӟt:">XX�Ǽ9�0ˑu���$����E�l�-��G��p�MF��Y����꾘���Mβ�HE�?(��"ȴ���E��-�ޡv��F��Q��h�t��{�{;��7� ��}NH��� �^��]Iyn��%�m3���䧑���\>��DOv�nM���`�:a�-3��2�p���� �����:�+!�+�H��O�x8��y��eW�c��==��8"s��>Nx�n���9�&X0'Ybe���"��r��;���K�.CbbcHy�*f����ݫ��4��	�0q����n�Ğ�;;q>�6	˞z-m&���=@��%���"l��'�N�7_�A��O��R}��](Mc��2'�n�x��GUo���bb[v�^�A�h+�6#i3@A:����zz�u1<�)���"�i�r��	�1#�g�Zj��Tȡ~S[y��V2�K������Zp���4�����-;9+��xm�Vej�w�Ess�GaK��^T)h��Z���C&�07�İT_�rH�V��߉w���X1�6F��ډ�
�Є��q�D_|����V+}��W�ǯ23f!��[B��x�I7
�p�;�s"�l e���9p�k�h�:~B]`��]����i�J��3λ	p�k�N�F��L^'�d��}��F`,�[���<��*,�KJ���idb��0f�.���M?��ʒ��K
Y��v���Eg�u{�lD��5�Eߋ$%���΋k�f�ه��6�蓤J�]O[�g��̴L��e`�@76�<��_9y�)�����Eԯ�� �CA�����X���M����>dk6.e��2L}�5�>�Ê�VAӎN�:͍2���Jj���S-���$�μ�v��7o����@v���Ȧm��.Q̆85���;�ڮ�=�y�$��A�P_6:e����rm��9"�섦�]`X��]����f U�O���-�W�{c!��q��y0��dn�#��f/�c�wy牁U6|���Ǚ�C�9t����Xt�ao�`c���rV�F�U��NA��׀e
�u|_��2�?ȑ'�b)�Ƃ8G�0;��%���/���Y����=	���~rK�Δ�}ARn�c��șs�1�
H�4��PI�g��Y�p��� R�]#��Mc�Q
m���ū�7+�HN�&g���m+�f��dYoƅ����V���R�W�j�VNnx�a�n���γ��e/�n�M�%D�bAݚ
>W�|(IkP�L&ғy�X�ݽ�W��'k���bA���뤌>��vÙ�_�J�w��q�aA���P+{>����J?�E�IK�:Ar����F��ϲ;�f��X��i�s�j|��{^�?�D�:��L7�l���"V�]x�Ke���l���TϴS؝d)i7�U`�v;�ǧ��f���7�׾�;����Z�>^{�}k���B淂"A���nA��Ga��!q��=Ò#���@:ҥ���xS�F����"+-�a��	��t`���~����H�Jdp��>"�+	ā�h3Pi*=*�L�(K�f��ۄC�C;�I�vL.ˉ��8���=a6Z�;wPm�7�^��=ޛ��Xs�H*M�vuKa�L�*s\�jVn�V�#t+�g�s��\2��|�?GS�7���x���2'�S�$�%��7-��5�jވ a�T��0�h��MK�2ZC����6L��%��$D�xR��n�c�YHs��j���l��m ��/��AQ���B��=�޺PL�Jt���U�`�|����^���󝄄f�Qt��ѧ��������-s$��e�jVXd.���ՁF
�6/$P�jCi:W��ԩ���m����M	3�OZk�F6�Ԩ6�{S���2j�BWg���!ܭ����F�_q�W	�K�B�:��)���DJo�6����������P�Y�_��l��<[a.���K�s�c9�L�1MG�蕨��ނ������#G�c6��>�r���/e�L8,ڻ{���i�ؖs�X��і�@9�+�8N|S舥�?���u[��<)F*�b͟��ԗ��1�u,�3�@*-�=|Q��+��J���Tq��0����t�aQ�t��˝����0�,�����30-�2|�03$Tu֨bW�Q���,�Oz��+�hi��q�����pcAMş�憳U
���͐��n7��a�; �t�bVI��a�~�NF�N���(�"��$J3:Y�@��!(:;����A/l��} ��LC�L~`:�MNq�H$/j'ܵY�d`(�۠��o9�5�����DZ"��D��`��7���NTZS�j�ˮZ�n�1�n�(Rh�ѱn2��5 ��K�s�(�� �X��5��TϠ:������P%��~�f��&	���OFw���d#�g���Lv��1����ŏp�J�i� �xnJXG���R��%���QݙWT@3�u�PlR	8 ϠG���F�eK�-�����-*��=.�F<g�wsXr��\!�r5���Օ��5��٩4i90�=��H�	�)>~%1��ݸ���4�{���j��l�D֚�e�d�a<p�k���C���r�#����W�iu��3R�ET�H���6/�n�K[[���`�*�2��XW�^R3U@jݼ:aQ����Vp+|��ƍ�jZ���h�ez,&$DlԟX~��G;_�x�1~d�&}e	�a܏֪.�&�>���������M��W�cL�Ȥ�ʺ�"$�ˬ���8hU�H�Q{v49	���[�	zv�D��&��϶� �/;�(��yd�Z�:���H�|����nB�@�C��t�D%~�$�aP!8��S��{u�t���y�%��6'���b�4'85r��#"�gc�Jn�K��7��[�F��u���TJ�A
Uc�kF��b�B�M)t,2�,�޷�#i���$6���:�X-���.���x��fB� ���.��8{3n<��^"�*;
)c ��,#�nHE��^d�jT;���߱��	\p�a�]���@�>�p�Р�	p�7O���Ž?d�EQ���#�@�(�'5���?����P������������X��Ťv�-�����=���a�g�j��R����@��ߞ$f�����c!J9fe����Il��7�L�,���H�Ö�w�c,���z�~��
��	_�{������u.�4�Z��0�	�H���K��,i���/%W��T���R1�3fVͳ�HZ9ll&���HBr�$�:q�����MA>(ffw�z�!b�lm��7��&*�L7lr[`=���^B��+�a����� +�v�!0v�H���O[����Vv]�r���=֔�ˁ�s�^p<� �t�j���Uc��?%���ʲB���'�\��Zs�tb�p!�GO���S$8��1�X���P*-��Gq�ǜ���Q�ֆ����@��M���4����:=Ëz� ��1�|�=�8���ꢲcf���m�L���4O�'�����	����fK�k0I�0U�9Tp�	��0�����T˳�>�F��e��ġ/����2U����|����kj��xęd����Y���jY���Bx>~��L��q�<��	�8��yli��k	܎}��ZRg+"%������fO����#~='jy�������l�Q�Pߓ�e��rޚ����VQM�.��E��wb�Kq8������ �:���h��o���o�0b�̵�c�N�lB�N�u��G�	�R�~
��Vx�N>%�����p���6s�*�5}A� /vz���3��ܙ�	�i�⳸�dj�gc��^0%����p�w/jbkR���=Gk�f �W�	��lw��c�>ts����p�t�U�"P����%8.E>�.� ��{x��y2���6Kh�[����RG=��[�'k)GKX�0z�P*�+/X�º�M�_>f@X��D�\�����hvrL5�(_�����L�C��b�B6l�}�N?|�"~V"�z��B��U�KU"m N���̆/�{�葁��Wt�Y�	�,eZ���H���ohlu�`���E?�M��tݣ�F������؁ί�!ЇCb��!����5����5���qv�mC��UG)��d���f�l���整�h��f�c�}%�����GE�[���[_3�aQ@���6(�o��{/���yf|ș����IdȮp��\6Lta�ж��vj���X1_���Q�gX�oU4q��=������<@y����)�Q1�D��F׽�]���h%�ٌ�~��,�bd�r[l	�\��z�������/Y��h%�*��#*H��ݰu�ݫ�i�G$d~"�;�vx�1&=��x�s�4�)��$b�^1���G�kZ��j%���N�ݫ���L׍ �}m�m�P�δ�#5֏�.�#�Z�#Bb�nǅV���t�\�����7��:�5(��v �J����]Ö�@h��Bjb�8�F�G�)&g5�N'Ѩ�]>A"Iq�#j���
�?~ �<vw2?�ڞ���e�A����5j��$�oe�G,�l��׃.��D�(T(�U���~�ՁM��T�K��#�UиnD�������b��zT�=�A!r�L��v4^G���ow�k�dƺ���@F/�gQ$���g��lƫ-)}��p���.�g���In�y�=�~�}~�̪�ִ�v��-����@/Ac;|"� I3:�-EGj*���0 �����k[MQZQ�M{b�����{��os�N۽+�xjB�;�n'	��X���ة�e���`-h��8��#�nՌ����h��)E	�����}8�8��\�6ᗝD�yG��&�\N����;�c�e�\4-����s`��ѯ�����C>�&�ĩ��76a����|N<^��qw�����Qg,�`�s�E��{��k�BvI�(\v�;����ʾ�F�Z���q|�i5��>�;�<�d��/JJi|1ƿ�x������6"�ߴ˼Wq�Y@|-���|��A�ъ�/��0��{�� �h����Uyk(2!B�˨��	×�[�������_)�p�%8�J�SJ�p�8+�RJ��{��~�i-�B!���g�n�Z�*�ZH�ٮ#Z���I6@��h�^�L�w�k�5��1L9�h�ct����c�{+h�q�U��)V'�<;"�:c�Uv�4����`t�Lo1�`ȕ�a�TҾ �7�yu|����1I:���+����(&�^�w�QE�j׃�tM&���ߙ�%G��QD&���G`R���@o)IkC Y���.�� 0������Rۢ62B��6�7���������}Y��|4.����M�S����[>����6Ś���n�ߛ1�p8�"��<�o�ʔ�A�g��d������^�<`�=��J/xX�]�m{��3���Ց�eln������,r�.\I��?,ԯ�xKU	����ߕ���X���O)̩��Jwxwa��	�
^#q����������&�`�)!ӈ�E񻯳RK�Ӊ,���M�H��mg�;�=�q{Ax`G�x�iX�w+��#�X�v�x�m�MOX��:K�v��s^G+�
��:��o��e	l���� G��!������B�Wv���w���.0E`��hZ�(��m���m%3���&��80~�5�Q���ܤ�lN8�A0ǼN�;���/)����d&:���FPLb���ؗr��/�E�ѱ6��ʕ�����m tҪ�:��L|A$W�����vA��3�8��7%�!�0����d�t������h'�8���b�Dj���=N�b�L23�_p�������_B6�ߪ-���)b�������Ҍ�?=�f��,X9���V"�7��N��_#"l� �]��D5��oSP�_��Z@`ϲ����a�L�S��/�j�i�L�0W�ΣNݭ���.�D���w#4���e���+?�_ecG-�uB�!�wi����,XA��W`��X����f��hxO`O���V�7L�b���t����@.;�R��om��lN�t��_NQ��D+v�:��B 7Hy���)�yq�MH��c���M
MJu4�_˭�@1�9X�n���.\M��_3�����ٿ��O��4�oY�}��0��D�]~���%E9�M|g��	��h&8˹�7H7��=�5�T�x��1����B��1�A�\�5�W@W7�E��ՎO�����A}ܕ*������o�BZ��XюÍ�^���V�~x!)e�\e6{pw��VzS1��o�F#�-j�OL�߃b;�°rP�	���E�(H]��O���W��}�֥�|VIG���%�����l%uG�������+��W}����*A�[��,��ӂ}��1���5�|�+z9@���ac���)XL�Ό�#�c4��E�dp!�����t����A��p�9{���I*�x{e�1�!�x;YB-��� d>��+,�n:X8}���8l�'����Y'�,���&y5^u��?~ctj�~}�,=�R���,A
ReR����2c��q�[m/2�/�D�V%1�b��>O�ʻ_:����f��y��ְ�U#��w�+��� &h��� A$3�{�Py��(E��� ��X|,��j���z��<�����P�ET�uXu��ڿC��	Y(A�����+��4����0���!�sf��.2z�/AI�B�=�,'O�!����;������6ܵo���>��.{���5W8_�뺽�������t��̛�{c1D���G�XRo�q?\ȗ���!9?;_ɻX�g��� '�+e��-A��]U�3���+��u��\���m�����/�ą�ⱷ�}���{�?Cˌ�4��0t� pwt��G���0��fi;�a+	&�3[�� ,"��~l yC���F�D�
�{��0��{g^��D"�r�=L��;T>k$qE�g���n�N�}�u�v�r�Ĝe�T+��)]�FAb������	}����{���3	�8�|�A�(������R!#�Q�Ȃ����MO_�����g5Sx����I��H�J��F�[��O4y�88��f�͆ �^��{�q9?Z}@c[������B��.���mܸ3t� E�tN7�`�_���a�yy�R�9���cʶ>V��)��T��̧(f�@Æ5�Q�@�HG�J<rN���]�>=<��}�,��,��/��UF+m�:�N퐢cǢG� �����L��{-f=�I=�BT��bY��m���F�����P��ŏ�6���e��䷤c�"��D0��V8`��f�-90bTb9�1s�_,������w
�H�����fm�p�1@���H|�~VǗ�[�"Fˏ�UT�L�Ȑ]�o���~����ޛ���Z����X\ �3 ס7r��4�<��jܫ}�F�h~�~����2̑+q���3�ɂ�l��i�*�-�U������BRY���F��! �ߕ&/�g��w��"�;7E�k�f�>�䕕�0�X�1`��V��g���������Š\�z��֓#UmǨ�Y���,0 ��Ueg&e�1<A�`��b��pV	�}8d����3)�e �ZP��M�6���Tg�����bwx���L
\�V�2]��(��H=�����?�n(U��;N�yUc͆;q��(>�l��Q`��}"?�� ��p����=�ȏ\�&r�����D;�Z�?�����<'7�2C���"�$V���#�#��ڸ����k���0�m;�q<�+;��:r�� ���:�a�&�	痬�<R;kF7����2�̼ 5�WW��ٗO[/O�g�J���$��ޟДVY�����L�K���9HԘ(�ش�)\b3�|⹘پX�z0��Η&@)U�;!�WA�.���%{��F.�Bx՜��Х���Ğ�����$v}[�
n�뚉Y����L�3TwZ_��$Nxj&�y�i�)Spwi%P�,�����k��6�U�}羴r�Ґ�K	⑷+��`�t�?��N'l�yv���o�v�w�z�g��׈��A��!1&�F;،j�>��n��(`�ygN�!MeͨR��"X��T3��`�^g}�S��K5��P�z�쒲46��'�bCv_�8���q�j-|~����C1�@V7+�IaoQ�,8<�i���X��yBz�W}��YqÏ�S��sl�豱�Y:��+��u����_���4�ޜϬ��y~��X��f
�?"Sa�m;��E:��{N�f�\�KZm�������F/�:7��#��
� �6�-��P0r'B<>\�;E�����c��$��&�x�-�ζ�a3|J� ���5��;a�A�aV�$hX���%�Iʎ��*4U�	#�-����E���S����m;�4��y}�S�����+�D>)�OHR���BC��?@���?e]|+�ZI�Z"��1��v���������D8 ��0����+�SXy�8���Rw������栚��p+����Π��[�|�G\�o�T�����V��"�-Zokj���+v�!��A�����3�c�[�B�!�F󼪀����fz�j>�W$�F������9�O�(v�B��#����$ۑ�$����?@��eV�A���#:s���յ棐d��9�6,�)OPW��$��A��E���G��H�cJ�WA�A8{�$�s_@-,��b4�Ißj�Ml���Ϙ���Y��$�N�����Ȭ�P��|��f,�tL������Rg��L�3��B����i��1@�05g����g���͡��������X�pSR�Ն�����P��bᎸM�&�{"v0�b�&�qbU�Kly�ڈc�"��'�Y�j�&�b/���}���/$)��]����-�\���i,��h4�)_V�Ѹ^���P죐^�)��$E䀓��X,�B�T:���+�X�=�N,�>� k���T;�}²�$���P�.��*ׯ��`�V����K���c��~e�p8��<}�6���3{mNى����^1�4�Qg�E�[	�.id=�+P��"�ɿoW��,�-�������o�1�S�*��%��tZ�\�A{��=�E�����;f�n��C�����5�qꄖeV:�����)ʉj�����4`�u	7�� �a��x.�M�*oi�83��� ]���PzW��=���D�fK�ap����Cgr�J�����i��}��7-�Lv����������[ J]>�g�l��E4�E���z ���E��.��zx)ʚ��"�|�ww@�qE���W����e8~�dEO�!��یS�'p��W�8�jc�uf�63j�j�S�����<�=����{M����"Xf�	h%���� ���L��RjI�h{�IE���n�C���g��5���/�{��Y�S�d4��SV�VR�������KwZ</�b�Rp���c�$}K'˳�!9�7n�u�W����*j*ڍd�Ĵ�CD��2铎gО҇�z[�dR�[n4j�Sd��{�\ Y��n>��2�$�㥐�,�S��	�4����Sg���l�Rmr�w���B�&yƏT=V���;2q�1_�$���qG� ���l��q�[Qſae�j~�W��������Ĩ)&�rS g��|܀��ʹ�g�P���Z~_���SR��O0���2^�.d����.a�v��/w����v���J���� ؞��V+)*���I����'^zB�����G�	˅X�r<�6����?�B�Qb�6�z�S����C�M~��Ş/���7υ\���T�~�2��g�/L�̮�i�d�g^�"Q	PZ/�Z�!��H�s��b�J���-�ۛ�V�5-󌚚��F1N� [��W�'\W�$�1�N�Mmg�W��jC	�g��ޚֺ��6����9�6V�DQE(�j��>��S�,�s���k�F�:#���č,�_��"�F����4�iC��K�\VLBa���h�B��FX撳�- Dp�g2���r�TiA\n�b��&�Q�n{ N�v;�F���[�A0�1��p)�g��emXr�o\\ ��C��_%�f#���f��)�*�/e�!�H��>���-:��Fi�@%�pI�D�<�s4�w[�j��ۉ��(Jl����Y��n!���RiR�T-�͑�J,���3?*.�=*�F/�tƲn�4*7�j��~�"�op��zpx�����~��2����v��!��{Z�j�%���J�\^;�{��'��=Cy�Wd�a��.�L��L/����@�^-、4�=R/y��D�~���?�˶��yR���=��]�[�C}fc��V����*���+������� \x5`�J��%2�5��3ErY�ٟYm���*�����'^���b�
� �;N��O	�\���"\�>�9���m���_[��n�J��hfNѝ��n��R|V���eDW�I�l�T��5*��x����c|(7�ɢra�'B+�z~���T}�"V~k�����O�-�`��I��W����"@E����j%��ޏ�ǶD��R���9�n<�l��R�l��F�%)%�hG=��Q>.�6݈Ȃ��uZ���>�q��?��F^�:����_)��`��Ν#�V��!ߦ���q�Y�ii.�K��6�F a��j�Jn�a��>�:k�(��IA,�[ä�	Gܻ �1g9�ܬvX�~�PF�Oi/.�Ԥ3�k� )�Ik&LB����2V���W:%��y�Rv{ʢ?+v:���{g�I����DJW��_$�"��om��ڄ��S�fyq?�����b��@�v�ұ�?n��������*��v�_+rH�>�0^[xw%��%� �s\�N������~ޒ�ؐNe�9�p�{T�	�SS���$$6�J���������3��<.�:^�܆�t��ą�vO6�#�#�>��q��,�F��<���RY4�o�C����`��س�sʠɔ��Qx��U�� ���~�h�=rA�����4�	e��P�dK��a���G��ˈ���BX�9w�SK�3�� s`*�|*;N��}�J6�m�3	p��X��?�rH"0�*��G�~��C�6輳ew�6(?b85���7G*}%��}y�ۨ��=	�\�|��oAM��8�~�K9�E���0"��ǥ��RpCP��iR�Ȃ��C��2���ͧ���+�_xj�oq��(�/� �`_˺�� ֖|�
֥�� R.@:��ԙE�z��B.����di��9��h�PK��-����1�J��/v�����E���r�L�T"OߓgQ=X��s�5�{�#��`���̲*)��g]Et4wg~�
�
a�c��+��\�R�{Z����߹_�� �ؗJ�}���=ҡ��8#Ԟ�",������dVZ��4kZ8G�:q1�6y?cB��iN��:������q�Z~i��{����j_�&�G9�g�#G��C��q�Sx���l�C8��u��)���������d�.�1!�nU�v**g�a�ҷ�]-�Ƚ��H)Ù�OȘT����ϲ"��DYZ:+��ެ}�y�J�Ԣ�����]�����\Xna���� ~	j�/l @�QT��a��r4�­���0d	nOg���AM��u�*,��S�N@,�%���X���u?���=�it�s7˲2��w�݋˱�Jt�H���(�@j�q��1��@m����'�{o��sj"�p ��Y��@��h�z��Ȝ�F6l:a�E2Nnr�F-'�n��Hd\%Ϙځ����zzײT�������t�f�u.}i�wg$T,���e�斚���Gǳ����67U����Xݤ��p*��!1��#� �A��7��/0�:)QKN��7`�� o�|2��ce�� �ǩՈ�$v�#��}�0o)۠�o�0���_����jP
��N�h� ��`�� F:�:om��v���p�<e����U�Y�,�b�����Q*Le��j�J"^�ۊi
^ꠥmDͱ�>�c�+Λ�'::��}�$��C)o���F:>���gm�?��H�e��Z!\.��M�6��^�#��t�**B���
� S>��I^�H�c���{��%�x�{�p�F���_Q����3��-�����F��`��(����m{|��=�1b�������Y��j���őF��[I|-bA�T���K��%�yB��I�pT((���l.�擷?n�/#VMt�YZ���o�:���E]<T�o+���P���������T_洩��/����Y�"��i�w��������Q`�ny�5��!�Rd��-�Tv�ٖ�Q�� ���4��"�e��'K�J��`�9�u�U��n6&�E��q���/qv��C���L�CdRu��(�Kl=%䈎��&��W_)�^\���5�?��T`5-ϐ�?���j�����j$=�o����6��狳��'����5�e2�z���-l��ng�@'y}.�H�js�A/T�`˫���Gy�s��;�hv"�vrP(�/�ž~/���O_9o�"�-j�{�?�L�n�&Iw�mZ�a�$u�%-�3��V��fB��}��E����5�xH���]i�g	(�PTh���(ɋ,he�B�w_�{HMAA�y�m��n�Q9�;�ں��2�;���D�M!�:!h�9P=B�s�a��L����[he��W�6�fHs�f��-`�j�>��A!Xz��Z�{R��T����cH$�`�H9�=�y	�ȅzVg#;����{�Ŧ���>�� ?����k!��!&�;��������������:%�$��,ƫ����ެA�Kc���������^��$+�[
�|�>閿��>�~9�?A��â�	�� -Y�"&�`s-6C?1V�m�ZZ�VQc4��\V�@6�{��p���j!���������nĸ��'ι[^^'�lE~��l���UvE}����݊/_�50P���D��!�+�o��+����X6z��H�(�f�Z��=��F�aV�rrAߕ!�� �����Q�_U�$ϕ ��>1�z�j6�ƹ�s��aS�������������̱ͤRk�}~�V����K��l|ԓ
>��R�o���o��}iw�x;V-jlј�'kI~��`��3wQ5",��d��Y�R:�Q2@�f�aΒ��C��`�ٿ��J�/_~u,4�n3D�B)��on���{&Ȇ�^[4�X��tw6h�e��>��T��_�C@��O�prf������,��U�Pj|->z��-T(�jbR�H���AԪ�_Kc��sa����n^4z��plbZ>�`�vjX��u%g$����(p� �&�w�)|����n%s�m�y�w���\D=�-I����O�b�Ş���$]�ޥI+E���|��P�	T�,O�����m��+P0�=wՔ��j�6i
�������C%4�p����F����srn�2�E���%ӹ���Ƅa.�z��B؁�詮n?z�[GOTOȔ��U�sxY@�ժW�3�	�R==��?w�a<A��WP��T�>�͡3U�d�*kTd�^�S��d|쬷>�na|���F��(��ٲ� �fS�)�}��+1Ը��i�>�E��>e�f�_[�`6ά�gÖ�����x�k����j��2�A�vfTA�aT��������@�DVD�N?��a��H�T�lVٔ���9TN�Z�WD}�3ʉ����p��D0c�u.7�6��9-*v��z�#uzF3�^p����uğmI{v����Mn���t�3��<a�O�oي/�:_U��M����-���ĳ�#�lE^��WJ�J��l�_nR����T���>*"�LKPw�T��<���h{Wŧs��+Bf�����Gn�P�[&w<�e-b=�W�a��+shMe��������w�ݔ� �*�L��ѻh�@\�QOtj�����"�|�[z������R'�1|p��
|Z�	F}�h-΋+�Ƹ�~4שN�?���~T����z`?p?��b�A�����LM�6�lxR��3//EsM���2>���f�&��ڪs��o�2qԢx����˘י�Ȉu���<�C��۲b� ����
��:��H(Ȏ�=T�5�W,̋w�^3<��Q��t������g����Qx��	��u�v��-���}y��r�|�����0�7j���"0������Q�m�\���}
��W�>�9oIoO��~Vgm�"�����XgQ�����K�L�v�mT�?�9�һ8��fĂ,���1&��p+�P1��ktZ=����YH����هUc��w��u�C�`L�M�}(����O�ك�����h%n�����\�i��H{��&q��MXw����g.p���Y'�}���i�S&p��U���m�ҵ�>�BP#��,�?u���Ai�,W1$f���R,(��b|)ѵ�@�
�;Ȳ�&�U�=��z�0{�)NFd����&�D�xw�r�,�����˹���#R��&	Й���!���
��Qqؤ��v����$�u��� 7��3���g����u��[�ֶ�?F�W�<`�E�q=�6	>��ҩ�S�-N<n�Ax��܍�T(ܱA���XB��Yg<���H�����e�s]���z��j�<A�@~�Z�2�uqg���p�����Al7_lQ��j"��d��<��s0W}5�h�hZ�hu�E��Hj��0n1ki��U�픮k�o�+�?u8}�ȕߙ�X�K�l�J��:���ܮ�Z�����ntİ7�Hjf�Z@�{ꠢ^D����W�I(	�l����_�]�	�n�d�E^��){r�E�o>�����j��V�s�51�v�݌'Qh"U=&�gOĭ�bnmfJ�$�jcK���X}O���!����ZC���x�(����ni ̍UV⇝~��Y8,���"9�\=��:�ȝW �3{ؾf/�����||��uNY���C�i��3W�$ؾ��z�"8"Ὠ#-���b�n?�X"կAc"x䌂$�)a�էA����ބ�[�����5!rZD�I���F�Xɋ*�s�O�6�x7Jǅk�����[c0���;)&���G1vX���~>�m`���:�e�N OK#�Y�z��
$.+=��uJ���N]1�0v���r�h�����L�߱k��:r���r|HR��.'_v@����j }��= *��.&az�6��<
~�}W��Ntf�b��LN�_����S�r�^ ������^<'Z�V-�6V�B�l��B����e�?u��8����ģ.�K��I�E���=*�����8/4@0�t����u욈:��Bm���9lcFRZ�L�"�|���t� �����~�  Gx�D� 7�5TB|�IJ}JO���@�{���C��I��jR�r:`���.\�p�ʱf�ׁ����
A0Y��� q�"g��^5g3��4��	�g��V����+(��ϳG{��ʌ�a�%q��{���g�yV��n�p��3�J ��p�C�mN׶��o�0��y�:)%a�4MRI����K7��Z�7��$�~<���}�ݥ4��D���ᯯ�/�/*�ŚD!��&Y��wM5 �d�L�8$�rǫkV��5;/)���P�?�:ON����-��f�J��#�8��~l5�a�K{2|!��s��3!''{ns�7��[��ΑAݚq��U��q)
U܃��7��tBN��	�q��\���ôr�Ǌ~@a2�Y|��h�H�}�]��Y	��^�a���1�<X�r�N��=d�~����
��X�eϠྑ�z�#>�n��sɦ+�9��!W�vW�%}Nl��V��+|��㚖��~ȫ�OK 5����r��]8������@1��m {ed���kp��G��~�?i/,�<B	yd<Y��k�m1�efY�����B8cRq�w���KJC�!���C7���&J��{^m�;���b��!ޘ�&�R�]b�L?�����c�Ђ�@ ʐ�2�k�������p�H�6��&Xf`p��+�P�$���a1/~�x�v���;��4�/1��M�3y'NOy����	׋�%���L6��.ރa���XU����d���y�)s'�H4��8��ӿ���*w�`0CC�j�[�.�_�
�e�Z���KtX��Z��|��z�.�3SK�G��z'�A��f_Ba��p���Ù���`��S���Yx��Q�ѐ�� p�A;���j���?�Y�N����h�A[��Z�4��z��F=�̺��K�g���:�P�H�h׬�l�n%����:�T�S�t�2�S��cI�����ށ��E,&�ؤ�։G�x�{����k-���ci�;�`z��B���mdq�K�=,Z)�3���t�b⦟7��J1:j��;M�J�)������mƱ��h$�)ݨY�R��F�g!���k8���qk��j�h�V5�'�rb^�pT"�"-�f�$�m�%K��ʪ�8Q1\�8����_WgW���*�0U�`C��/A�?S��	�x�2J�� J��Gz��廽mF�H5_�8��.S�!�_�v�(N�y8���.�n�3�b���W1���t6MFS�S@_O�֖��B�ǑPBr��o

���7"���1x'�8�W;z]�M�͡��f*�e�'�"���?+�	W�S�U��X'�JKt�	��_���8yFݹ�Q��'�l/�ۇN	O�7A7^gr;��A�Ֆ����s9j#��M3W�4g� 5����G��zAf8e]�`���d�4bz0�R~��}k�~.����e��p�A�p1���h��o[����,����|:ڷ�E����褽�h�y]���|:�����/���6���ݏ �����𢡄&��9s�����c�"ĺ8r���ڒ~28y��v�����?�O2����y����l)h�n�t��ۖ��ۈ��M]��d堫�V��gw-܃��wD�dsh�@��\�!rh*::
! ��=ٖ�
�H�_,�T�n��8k��paςQ
UY��;^���Zl ����Zf$���xi��Κ`�W輹�3����ř�/Du���̺�k��H�=Q��8�_���>�U�zl"ȧ��ܯ�p��(i��f���%x���m���L����L�ymU�f��;�_,�e�nSM�R"P�`�M"���=�cDZ.8���|�`)���r6�j�5}Uf͚�A���M������+&&Wײ%l|`lZ�TA�!����g�3#�0�������Kƣv<�!�� ���i��\mH�!O����$��"J��D�J��-˷�	L���a��5��f�g�������L	�y���RЁTxF�OQ|��=;;$��y�����������<lNC�V!?H�m-���}7�lJ%ڠݿӒ��ܫ�S��,�8WP��kw�g����#�W^� |��
��M��P�J&��X���3��~;�!���d�����3��� US)-V�#y�s�Y��ٔ��}}���pq�.�v�������h��1��@I���Ma���d/7�{�`�ϺYԇ�������V�k�`q2�q���h)�S�7".�����J������L���D�c��f��FO�j���_iԖ�h<#��º����O.O��丗o�E}K)W��B�f|BS ��J[ n�^����Bՙ��3f��rd�Ǆ~��yc�?��
�l;�ObQ�`�gx�G��	�d����K�P G��	�./�]�n(�D�َd� �^0S�ϴ�����@'�X���S����#)Q��O��@��4i���� `�(&�:ݿ�ɉN��Y�����:�bd2�r�I�2��#���ᏻ'��AyA�Nq|v(ΐk6��C	>4�m�Cco!Ofo�}����N~�i S��a�i��3�����6�_Qh�eո���D(\=�2ח����ы��T�`��v�-+3~#�!�YkG�c�g6@8
 jۣTF&[�7�	S�7J<��Ny2�[�>^�O�k1�¾��&p !3~�t��§�p8���?�����%��-qv���u������T�5ፌ!��:�����:�Ε��;
(�ލ�aӲ�dHV����E6/��N��B�H@�R��o(�ې��C�4^����JF�`^版'���*3Z�(n�e���(�<���\���jv�
d��xr�d%&��/^�f��ku`�_f�>;'R��V���[[�PJâ���V��ݻ��O��R~�l�K_B$tH+�m��`��ڨ���o���RI~���ɮ_��
rQ���#)oR���O/��U��
v�"�/3#}yl+S��.��I������W���|��N�J�	���V��-�Q�Ubq��
Qn\��������R��4i�8��_�Ȉ79,:�y;�M�mr���85���D&F��`PB���:��.:;�}�6�i���|���z�B����E��kn��/_&������9�::
#Q�NicP�<1�֮6>'d��0���4 ~\"?���r�սx�.@��0~�BU�kWF3	\S�2���Kɜ.��T5�=�"�Qi{�r-�P�m�F��= D��>����iޅ �
����ֳ�y.����C�aӗ\�� ��iP����W�ت��<�b�$��%��0r���k��rQ��+�w���W�J����p+�e9S����P��d"W���On`�"!p�U_K J8ߍ���~V��8RL�	T0c���I�M��!p�X/�+���:1�V�;�괦?$h��{
˳��L&�0j�1�O��l7�����*D$���.ܬt^��bؒ�N�?��b��5('j���_�Y�K[
WTMb���L����m'����}P$�e��J(7��8cC�SdY�"YMʾȬJ���OY���y�@\s=���K�\�����F�鵙)�b����C�$)��>��g���	|����R��_���A4v6O�9�=�Tp#3���a7EN���P�=F_d�z���|���Տ��Ы�N���u�{�?�X!�:	 o�{�z�w��5kT-F��Tଥ��1bf���ȳ�Q�J�}3"3H(��Tۥ��2fve��ީ��J�yC���7	)]��"�0��&�`:�TہAfRͥ{�%�y���bxe�9MZ�������PAsO��4*Z�iB����l�=��%��g({�٘0�aF�ByK��=rh��$�e�`��׿"�!�;CXf��z�If��}�����K��AC�GI�A^n/�#�u���,W�s�f� �U_%sIu�h��*�6�����xƛFi��4}A�F���I���-����e��-}�mn��RwA����%�f�9�f��(!�x��`�g�e>�ؘ�v�·��|&��zq_�JEX"M��H��04�ltR�a���a��Z���UTj1)-��7����8�20��V�}�W�z�4��$9������'�*��@���Ԉ�_�#���q��F���J�,J�j�K�	����9����VlboC<����t���'��w����U����rֆtq���p�%���h(٩H�	/B��u���|���clء�l�+�Շ1�E�I>���{DJ�1#�:���������~��<�m�y�(�r[�݊�p��Z\��|��
GD�X�,^�W��;���s���w��6��Af�Vm㿋?�Ŕ�a
R����[���"b�]9�.���.5���6��Lb�О�����"��W҆!,q��O��w�E��k��i�_Hv�*}��#�q�7�2f��;oO��\-�f}}����(S��9|q�N3�K�Ƃ���+ڒ���s7r������:.J�F � /6}`,��j���S�ұ��eQ�J�Ө��@`�ϝ
m�ǀt�VW�9���u`R=�7룝�.�q��Wh������cH5ET�m0[\�	��4Y�@$*��[jm�t�\��v�+��#�SLK�>c��Wx��xl��y�D� |����M��,q�������7�d�f-��2����B�T*�����̵��0�W����#�;�j�v�(%�}u�:�j�E���	b��#��nVfs#�w��Y�E3��=V�/he?PA�7-/e�2!5��B1XW(x���R�L8�h*�WC�T��y�8��	����'|U�5�,�uu��ݶ��9�`�֞,\:?7�$�Am# ٯ��r3��QHdR���-܅�r�Ug���ї�1<��t�YJ:)*���v)�5W���ztTw�R����oϑ�g)���_��{���ԙ,C��N���Z߈��:0��V5�)&�o��vt`I�%q��Ɛ��zY˓1���-��	 �I��Q?��6)��l�q�X�O�#� ��'z̦1g��ЪN�Q��z�}Ԅ�
}��ڙ�G&�0�գ��},N��5���D8G��~��B�#�p���ӥ��z�����vWr�R(F��k	�$�hd^�5�w��)(O ���B�JRG���D�9��HxH`���v��~,�ڦf�,�[�+���;����'�¤!b%�Ŧ#��!�v���.����Ց=�Ï_MK�㯿
0Ʈ��oo�E�%Թ!r��:�JQ�D^�\���̑�*�D}Zqڢ?�%#_�˾Բ(j�i�]��~���j>Bi�t��T���=���X���i`
�J&��y���F#]�����$p��.zy�:���\�?��'��O"��8��Cq �c hԕ��\όO@�u�K�4���g¼�0MF��S�2�:�c�JY%��7�,!I�^ڍR8lȘ!��6�0�id�����P�8���Y�A��q������F�������}F�e��H��}n����du�6(?�ڿ$@5Gy��{oS������VC{\�^���AU��IA�ǚ�6���:O�.5��u�cƹ����w�'Р(�����v��=����d��R�*�ڦ��MU��~��b�\�ŋ�~�40i��{-ʝ��~�l���GU'=RE��:�[�V���v�B8�B�e�p�Fe����Y�� y4j=7Un�d��u�x������oǣ������V1ٕI���*l��X�Jx�L(�(��ݳ!�����w��n[�Y�?��|�<��6Z
*�.��f��W��6h���_w0����ٰ���Y��÷�O5����>��D�~���J�U�0ȝZY��{��HǨ7q{�#,Y%�}��!���w�@�0���%��*I��@�׬'o��1�+�@�V��1�cf�%+��tD���Z؆��������Qu���������%�b¿K8yx!P�,�b7���F#ͶLh�7�#|	~���cH����z�&q�JI���W�TJ� ��RA�>Ow��:���&_o#�b9�� ����A�#_�f�ܢ���R�(��p����y��c�1qzF�"�T����S�����7�j�ل��}���Ie���%M��L%6��t���4ѩ1چ&��B�s��m!����*bi�����]f	�H=)MN�����q���ӊ��!�ً���x�c��]��.o��ou�T�>�0�?����wJ+Zs��F�E�[�R���u:����L��_��H&�2͜r_<S�*����#\��wb�f�=��?�g����(� �1���H��&[�׼�����-��������X��y:f5z����"�a;�"���5	]��ޞ��Px�'ϓZ�r����P�#�4���-�DOgz4y�6@����-7~?=jy�$U���V� ��W&� ة�)N%�[�g��t�}�lb�qG��ku���K�������r�Po�
�.�z�PW�9�r��y�F��&i�a׆�jb,�3��_L=����aѾW�F��/4�W��K`�Ku7l5�T�i��}nEq��ڒ�yc�c*��"lK�@ϲ+�!�SO�:��
�����(T��"�<��z�ʽ�·La����3�l��� 
i�V� �D�|ݴNGe�^e�4Դ�������5X�oR%�*"w�	�8g�W%}��xU�k�c~�^$��)��+�>��Mx� Q%�}�/���~����kVF�m�i&�K`42,�0�۸{S<��h����7�]V�.O�8��t͌Qj�ѧ�?�`��iu�>�RJO�>RŴ��kvZ�ZWW�ۧ�
`�wh����ג4T�j�@c���4���*8e{�P��Y#8,"ɜ$�I�3�=�^[��^�b�'_]�@~rJHI��NUI:�`��ƕ��$B r`Q���A����!:��p6R��������b�_��+�&Ope�K��hPa�,����?>� hM"zj�%O�֚t�R�i��K �,@$.��V9�n���I{������J�xS1t2��}͵�Ï�;\���Ϊ5%ϯ���t��ez�&D�R�`/��x�՝���U��M���bm����t$�I��X��<�#�8ȩ������̖*���!9kR�(Mr��
~?���0�"����mU+�����̡�iy���5�DԐ<��q'����s$)��J�r.o��0�j]�ŹD��Fr�>��I;��ٟq��&��:*䯭˥�����:aި-(�-w��1
��PIL��n���2�Ne_yw.���L��d,ߋ#��h��zZn�.�����5��uV����]���4W�G0�K���*�����4��ţ���p�4��^� h�p�N� �=dp�=�U�B�����Wɨ�,�ʁ�㝄0W_0��1L��}��9�n-�{ĴO�/O�a�n[y�!Myz�B͹k����T��܏��Z���Mx,��첋$�~�w���������9�zn%�ǯ�rmtcB�f�k���M@]�^�]ܓ�j8Y�@�����.uT��&�[JF��a���L]�K�!��ɪ��_ME��;��]��	���~a������L0�%X>���)F��o>�N(�V�XqhfM�{r1�ņQ���1�wUe�6����S2PP��F�d��g(�?�
s�&A��]��u+H����6�@�L�{R�H����3<�Tn_�S"*nx�de(������7�J����������#7���t[��#����%O���q$y�a���#����GD�Kς�sd��jm��_8C�z]�
��X��b�0�����9(S���
&ȝ�%�>� jK��0���= �0-z;��fEK3]B@�D�l䗈�E��!h�.���멉�A�P?adQM{j�Ep&����DK�`���&W���c���5�K:�m�6�f<[�>�ߩC{]z��/0U����?p��_���u��&��8[���'�Mc�g��"A��C���RL�����8pp��)�)��(vu�,d&R$�ܶ���{�����h�-K����`�~���_��(4�n������C,�b����c��ByW�3���������;nh�2���ĺ �NKᒖ8$)�ޙ����.	�0P�/9!�����	�7����k��)�m�2R���վ.'��b&���q6�$ e��ϡ`&oa�)LT�[N�9���3c�b�J��[���4E��ϓ9s'�b���zQzyը��j+M��Ui�x5�2(3k�>mh��S@4l�A�U'3.�*+�Q7�9��|:�,�<B7!6֕��a��k�KQI�\�y1�3bg �
"(��m�Eͻ�24�����E}��`m)}��c�n���SN�_���u�X�u��\�\Ƥm����QB�ȸr#5шh�/^a|��בt�ҪLq�]mdɑ@:���\�^�Ki��R�x2<��G;>#�x֮��(ď%̘�hB��v/��2hF�44��u"+�A�?�z�f�bd����뙆[g`�$�D��WaLG/�|Η��v,����U��o��@��y����q�:�ٕ*�\~Îv�����]��u6��*}A�D�%<�*�O�6�rH�C?�0RI��,0�[�vZT��lf�k
�-��2FINh|�ɉ��tG�x�sh	𳯖�7��e�K�����sA�R���E�-�T���+: ��bw;X���9֭B�f���v���Gq'���]�*2)r>�GbH�R�!��G�aP����������P�z��N�PR/���� ��sMA<`�x���Z*s����-?O�r�@2�1��KI�e���C�'�)��76�n����sKD��q>�J$9��g��uv�Zm;����'�n��t�IlR�b�
���w��ޖ�:��H�.?�����<l*n�[�Q��4�]l�y?��4���I�u5���_�>��")��Y
`�S����[�<�] �l+���.� L��}I���{B�?"�F��B`>��{9K����V<cͣ0��?Πe�3^�#����R�.Xh��g��oZ�'A�ٖXV�4Jݳ��ۿ�t��:f�@��ɕ(-Ҕ����>]�SF���d�S�7�8"9LY�׆R�y}Z��..�!���jRtp�FZ1I�	�f��z.ysjf�r��ڰ}�6�ѐ��&�h��;�Ѯ!��Hv��SD|�0o�|��bW��-]I���t��� ����W�R��&�Y~q��1-�rV�/�(e=�z��$J��׸�W����G(D��`�3�`S�S�ma�?0J���#�N�Oe�0 �mtTm�oU0�"��pD�v�1R�p������l���� ���X������4	��VV2�֌叴\���\n*v��a�'�É�tSHH�y�:��;7�H#k���6�W����#p����׌X���/��'M?=�7���o������� 9�%�����!	��[8�~9��3�yJ`a�D\O	�/�J�&��3��~��(*����J�\�0%°�7����� apD%�"26Ud���&��:e�Sý�;������:��h�k��p�R� �a�]��x�=�*.�-F7n�	I\kL˳x|"���oj��xz�@�nX�%`�y�̈́��5��=$��r_��A��q(^�|����F���������r֕:������+n}{C�w"	�2�4 ����"@<�3G��|�}w:��/OG=q�6�Wꍄ� t&�l'y�L�I�����$���O����m��;��|��8ۚwԮ��J<��_�\?k-��E)\��цe"������[O׈6m� 1܆vb
�h"%T��o�����$(Z�q�3��b�̳پ ��sm9��d�j�)�G7�Y��pc6@	H�T�wˠ����̾�h'mǬ�N+1
�����a5�1�}�E��[�Y?O��O�KI�������f8,�S���|��0�ݕ�,S��ؓV�Et��D c�#�A��?zj�����$o��/�J������F�p��^Gh�ޟ� Pܕ������y�c>��zJ�i��K��t�]D3����p�h�;u/��AT���N
���9 ���x��� _�^��c^�|�LU)s:�-r4z=|
��GsG"Q�+vL�cear�L�<y�ȿW�W�d��{�.��xN�NzY�ٛ;��9*��� �=�|a���Ip&a�'�l	�s-p�I�'xo1�nk|/�h�t�I�fmq��bRW7	�xi�;��:� z�J�+�eY�����R�|"	����%ֻ�Bq�8s�]�� E�V��~EQ��*��唶 �8�lg��؟�Bh}�=���Sʻ�Yi6�����	���f�CwX���])sU�v�q�+�<��Ӛ ���&�HRAz wT4�mn��Q o��)��+�oDoޤ�k�"$�/rT��_m�=1�}d��Hi9�Ĕ�ϵi��{^m���xͮ�� ���Q�9{ǽ��]��_'�ж�4d�bv|��gCCH4 Y�3�s66Q����r%�I{F`�]���!H0�Vk!;�,��:b�`���d}� 315�`W�*B�xud��,�ZV�/�|������N�+��E^	�xz�!���L��8]�E4ǁ?�����:|�D�?�G��V�L-��,���kW"1��z�K:�b٩I@��ϣ�kh[�3=�1^�>%
я%^�R�.�WE�722t�$]I>d�=�rՇ43XlU*� ?[-�qI����	p��b�YoL�.���w�����m�UГC�_l����Ѓ�M��HI���/E��=m~�XgE�^*}����˻��b*�0~9�#�>������ebn�:m$��9�mMQ�Z�@մ��CS }��22ʯ��Ժ��2H�4��9��ӊ.:=�����J���95m=�����;A��0��%,m�O�V#0V%;w�Td�M�Wʋ;Vfl�V[m�wH��+�I�9:������	�͗�9�R2� \?a�t*�}�J\��
�W����T�n�w�zy-jw������ѡ?����N�4��-�N�jOKb
�����ǀo�5Y��!��	� I�o�T�]M���v�A:8��bI���-���ssb+tP�|\�*ˌejc�un���Q��h�vnHZ��x��y_]CL%�"9�4��^�_D�V���Zk��C4(|{AŬ�y8~��_�r�.�O�T.���F�|z�d������ᥒ�x�L�Yщ��D|��o�����uȬ��u�kwMe��,ɣ@�-Z�@ڴ|=�Go�O���S0� �
=��ݒ�Nh��$��آ��q���W��ӵ�m�@Ъ�H����8��[��x��jq�C���~����{�]�Mׅ]wCa~&��/uJ��uu� EBv�bs�RΈ�C��ؕ�Į;�N�qR�?A�6,6@u��]�o��!uAH<m�p�c:��F�����Z�|^��_0����XV°����r����I�{�����i�UT�"�1W���A��A�q\]$g@b��B ����4������5	TM�)4�NJP��%��TJ�p�`��˄z��_-A��Y�Z0&����
�Ey�C����k?���iyy�J��#�Q[ ��E/l�j�\`h�ޭ�)���>�9��2����)4���t�
M/�(S��toZ 5F�b=�������(c�hP4�O0��:%��)�g:�*�hG�\�"Ŧ�����"��;]f|Id��{"޻���MBt�h��� 5�C��N��ꚦ��LA��̣v��k)��±�r�Z'�d;��ik�f�oX�n��n�"1����Nu
���� ��A7�l��)���5! $�_�{�\����>�,���M0��:0�h�f�ra�����<�i�f���5��n����Qa�9ON��Fɖ�� �c'`�^�[��0RM�}۷)��Ii�5��b6kRdL.�M�����.m�W��L;}��R/"�����P��@\��hd,M�.�q�a���w��/�5-F�M6����Rp�A��*�#(@*�ˀ.��~4oV�!��Ǉ<J��BdJ2�t��5l��J�<��_⁝Tv��VĸU���C�]}��צ�Aic�@�Vҹ�����}!��G0KGRӪ_�I,��Rj��a��#��C=�����%I�M�z���D��
�E�fQa�*���<$-̺0��N�����:y�<㢹%*�v��/m`C3$h��
��\*`�8�otI藕
-|r�='>M-���4{x���E�Q]`7�ekcX�Ow�CX���Z�yR�� �'���Z���:X�!��'�����P�!$���S�xl��p
�1���3�=���*K�<��eS��{b<jp�x>�A�#�R��{ZQ�f���/k��E��=��&�mx�J�v�#}��+ӌ8R58�ɴ��n�	jD�����*�v�knUqL��1|�Ö�I���@,��Y�E�gm��h��N��a<M�Ej�%�D��(5��2��� rK{X�Y)>�b�����Q�c7 v9�Q`m%�lV2d R��7>�a�!���!�Hohކ�֕<�P�&�4������Ӟ�p�V�EC8�����$��~&p']n��q#I�J��S5���W`��aϢ��{�#�`�������T<�`����:��o���P����3p�'e����8_l�52Y��+�L�����f'��\��pZ��&O)�l$9Y���G!�jY������r.��4f�KL�vo@�;�Y��0T�p��W1f�3;"� G�~�}W�	�a% 9�_��k;D�c��,�YV�صY	���&n?��]<���5Ov�&3]Rg����/��G����4�Mk+��D���u���XҠ�P);H�� p��Oxd٩�ݦv��������=�t�+��u*�МhE؀Y���y�/5��1��$i,#)�ʜI�nK)k��K#R�_�&a����}�%�V������V��㽝w����i_��kс�`�� 5iX���붊����/d�Cl� l}`�$���XWjt>�1�#z���t�^�|��f��pSo�j�NBk�}c�����d�>�c'�բc�3��JG T�-��ٽ�`�l�RF�,E�J¥c�[ЊnH���+S�K|F���Ꭱ����.�{��	�q��zԯP!J!�a�ӌ���x�NTId�+�a �KZ�{B�������EW�
۾�]��c5�PNF�(Rr�?,�Z�Q���Q�l�Lf���j>�ʆ,�-�!_`M��U�x&�Zo>e�m�8�G1c� q�7��:B�	]0�<<Ɉ��jm�~U�#I�aT��0C ि���-��N�vM��;z5:'NZ�<�hyqm3����-#�EJ�pq'>��͒wŖTm)�v�e�n�p ��Q�)0����/���a��Q(7�v�j#�Ez0�AZ+(F��
H��F���Kq^8/*�՗��_:��󍴗���m�ԽM��Q:J"d�wOl'C�\=?#�i/�`a���܃@3vI�Z�B��^(7w�͘k4�!���m�I��7��*HUg�w�Q���l$��݉���/��tVKw:�G��ص着�~�7�܉�3s	T���`���z�"����Z�m/^w�tt1ʹm<���&���B���7�-��
�����-�53T>���<��L��p]c�]*'�eꙀ+F�٢�J~c�28�`���)�� XJ,$�MT��G���`�!8����m��ȿۺ���Ϫ�y����Q�o7K�x���rP���y-F���+yZ�`=�&x��9���V+���ߵAF)����YC�qⷁR_�f���Y�.�V�D�1)i�Z�<z))��Io�T9_�"- S�Ե���$�m�Z�O�R�̴zY���`&er�����_���Sҡ'�f	@�2sH\��_,	'�mj'����^���VBQ���~s:>�H��!Q	� ם��Ȃ$�8����464�д=���R�O�	�%�4���3{�cb�l�N����F���D��@�Nk���������h)��@��x�W�%��l�s��sn�q�$�_�y�jv������or�vC(S0
A�����/0�4[�vc]�l_��l�����i,�c�Qb����(G֜i^0�6HL�-�_��d���^�K��Ϧz 䎖��Pa�Z�U-J�ry@W�?����T�~O���t����#�۳/�P�������T�K����Ey7@e��o��$(7`����#��Ed��F���L��pQ]��ߟé_kcu�&��}�U	�
gָ��=�t�c�♨��-�������k��E��vU����9�������m�q���'&:�����U�O�ݣ���R6�?o��԰qQ��tȳ]���A����b�t��럤�86���sܭ>��f�M��X��L�ɢf��v/q�BDވ�@�8�5�u��?���VD���F��=d���&cEZ�Ë����d�>�ôb�ᢰ�g�z�2�lks�Jr��s�+}�$����h�t�3���P��y�<���xZ��#j���u�E� �e�͉񘲪n��A3݈ye�cE��������BS��ҧ�I5�6��{'V���:��ަ�Ձ����B��'�'�{�w9ؐ��O�镂XP���E�$j�>�p갚��T��:���	�6�`��N�Tt�/����T�m���A(uj�J�������\���Pt|	��~U�V�u�1�8=2�Ch����pA�6�ìRx��%�fWŚ{.��3��6�$#�ѢOh!h3���B
J!����BK3�<VY��_�E�q�JH�W9i��M<�����ho_�W�GR�jT�8�Fte�V:�����V11H1Z�|-��50�{Z(}�z+�H@��_���h�֣0�����R�rmޥ���L����D>d�[w/�!!�WR���I��[�Q�!��S$�F��m�+zi-��%��Ő�c�qa��"���76�H���P�>3�a�dtD
U�lz�m~�F�U<��|��;�C�N�*(W���3��l�͍�� "�>7L	�H���gv�z��t
+��̸}���k�n����[�NWX� (C�-}��ʞ8D��Z�P��|���P�sjQ{��kc}np�~V������sˡY���w��o/]@���a�+�]FL QE��t��HZ�l42F�����1U���M�x������f��Y'��hP<_��0�ww��h�XQH����>�ɔ�����B(y�%��}8�_��-(�"�d�խ~	Ƹ��p�6�?����U����L�Ȑ����k��W ˡ�m��W��x����-�%+����)3-�Xq���3 `���iQ|�n���e��P�<�4
��x����a�`T�m�����n3ݷ�̈N/VV4����&?�7�f�^Q����g��~��]�9�	Ww�6BL��k���(�A�N>j�[,��j�W�`E�Ӽ6��=
UXP��uF=�=y��d���x����h�[�^�s�t���Kf}y���WkG1@�M��#��c6z����~!)]�u�m���!�y|x���ȡq�>o��I�B��Y�-��K	�w������*��K�ub�aRy����_�je���J��/)�l<�ʼ�4�g�������y�l���y��&[T�Cx��{UW$��\T&=��Ӛp��![��T�7"8�9W��,��-Z'V�e��8�(8�ҋ����~��u�.��0-Abg��o���e�p��j�Q0��&�vz����=ۈ��F� �eI�,W=�N�J���N<��6�~n<��X +p��fi��vEV1d�|�#����vz��q�P8;}���eNI�%�r��R5tcU@�2�Z+���9J�6�RN1vN���*��??�:Y�/�S��,�� "t�?b�&�o��z�㯑B .x:Z�����{6_)G2�����2׃�%%F�+8�7)"Q@�-(����R������A��� Ģ�K&q�Y�;�Ą���U�s.��7���Tt5�<0z1���^Jc�d�yU�e-^��k�~tY.�\ix�Q܁�Cu_�`�?~ʨ�J�8�&�;dH�g�bޢ)�*y8_��/@w�S�]o썔�Bj@���?�n����V�u�D�w�i�#>�ӻ_�FY�)����5�����	����e5"����?�Qvx$ym.��UA�n8L\�m!�*E�vk�8�*�)%�.b(Q���F҇�K�BUae��'kdΪ�ņWp���w�����6c�m�����ϻv�I��� ^ ���*��(����c���D��lA�e����p�I҂wĵ�$��i��T�xϣ6m�eזV=B>�A�H��^�v��,od��i�n����_�'�C6KGȚ�#�Ǆ<� ��Qh`�$�g/��Q	/l�I=��e������(�p�u�CB��±7;	�IJ`�fǑ�X�1�vJ��n��.�0���D�WB����=�b��M�!�+k�+��i���������{�혦T�Y��b�!D� �#}�Н�{���8u�!֥��5�pߠJ�&_�'���I`�����+�e aO�u"]���M�d0ƽ��'�������#��Qm���|[-Y��\�r�s�,��e�����j; �37��3�+�Rɚ����#߾O�ɿ��r�:�̨�Oa�H�� ��h�IZ-�{s��گ}���AWEܗ����,>�TM�&IKj�����6 �������Ĺ���5�r��H��xة������Z(�qT���զ��Q��[6=(tL�#ŗ䗱���?͝�Q����RԪ��/���pF��̻�^��N�+ ���>�H+�p�`��Y�T3嚱Cx+��֩�̯?4�܉��rP�&��Ug��;G�I�p��1r):�E%�a�^��5)���2ݲ����;t%7��A�Ĉ��3��>E�^h���p@U�<ބ�p9j�P*�B��J�R�hM��p8e9<���n�I<��">�Q��w ��w�QƯ����2�d���) �^�xc����8�OO����������-��{���}�x�j�7\$8bEII����0���T���f����=��W��\��n�Kd����ٗ�	���\]�Q�oTKs�z������Dk�l�ݝn��'q]�Q��=��������Wz�kz6�O��uU8�>���tZP~�&I�*@�łx���'�Qy�?��B�p�S���������fO�I���s�������8��;��-Oލf�׈ё0	�D�k��Z��zL�����/-yJ�<�,H*�����ivH�ug�v��U4M�F�V�?T�c�N��	�-Rߐ4��6%~��J*�zB�IE5M�z�v-K�$2��T��=@��1P@@5��ȵ�^@�{�u���S���;��'�­w*�����Ć.���y����II�d�GU���v<|ݦ�~��L��"ɒ;eBt�Z��|V5r�����27�#}6���DA?�D�v�-	9�-��i��#6�g�����C�� U�,��n��tz������RdD� ��׈����-���y�$x��ypЏ������r�-@�	�gasT!���f!ǉ�ET]�!w�P�=R��D���x��9�!\��2�v?@��i�v�';=���< �n���	���z��6��\+a��|Qa$�ןB�ͻ����ܬ��Ռ IDP}�HC��Ex���/z�"�:��/���J���}a�����v��>�5����.ab����?ˏ��l��8��4��)ibk	���؞��o|h�/�{�vR��dɨf�2ۺP��em���鐖Y$
5�B���t0v��TVb�WU�6W�������� ���W���
�=���/
������~%߇�gr[���i	ӛ�~�Y����}F1]�e��Ɉ�?:[j�}��Є���B:y�u����v�a\{�1��F���.H}��y�m3upn#WG�Vb��/�������ѐ��Ҹf��ωS���YO��b�y&��
�����5�1���R#C�!�s*[�A5��5P��������Π�+Z1Q�igJ��\YK���Dg�?bX�Z���o�َ��/��hl7��d~k~Z���EtC4� �T#=6��c���EC�{�'����8>GGO3s���� Veԣg+�Ư�&�н��s�n0��^`�2^�.0����!_94�+7)n>������m6s���d��9dw0��f�W��h��Q��I�l�!��qݽ�F
��w\�J'4�|C�7�7���g0z6-��k��Nv%�\�F�r�� �</.Ӿ�����Mi `pB�̽�31�?x����cXz���Zd:��9&s�o�4Új�hC	�%v�т��+{�ǳt�>͚��i�]	%=�c7U:4�.�Ȝ��f�U��$ڑ��FK��b��>�,�`���H��s�q�^O�� �W�����QK	
�J�>���F�jm4�M�;�X��}u�3������J�<qF��o�*�6��wW3"��~�L�	hA�k����0ӯ����@X�oS�L�d0I]���[.�v��!q&��2��U��m�?HTf蘵��_SCr�΂��w�s�S�	�_My��.�.9OP�"�Q�6ů�d�is��5:s �)SP�13b�����l��3���������|�r�x?K�Rs�4��G�$��	��o�ǡ	Hv����0� �%���ǚX�0��ZH۞��ڳ6*�pG6����@��(x�zi���"��+�V�c���t�K�����4���A��7�&��*^{�ǉ7�76�B�*���֋��H˝n�m7�'�/�H��G*�M�]t�����G��#h��-Q[bv�xu�����Z0
5�ǿ��g�F���^�M�[ZB
�rn:ԗwy�fp����/�KwDP�IK?�8~`���y-�X���1-J�k'�Zo4L7�?��"$3��ޟ��݊cER��1^S���,�Ĺ䵚8�y%vK���o��2�����ڿE�Wf�w��*ަ�ܧ'��BSe2��4�{N���M�d�&�(����^�����jR��=N�g��o�:D����q����`�g!~}%'�Q����2�͟�h/C�n�u���hpCٓ��RK��i]�,�5��FM77�����)�̎^{w0Iu�G�(��73���C���g�jmg �8����Bo�"\>/��h5_�$�C�[����${%��rF�^�)�v�D�"�_��))�����f4����B@Gu�yN(4(��+6�����i�a2#˜Sc�f� �bU�?�E�oS�Ԁ��X)���Oe�&�!��9B�K�x;�}��e�L��do�E�E.�ࢆȑٹJ=	{�C��K{��=�������n�N/z�^�8�����$ &�<�٠�3�M�-Srz�X��s.G��V{EQ�򱉧VV ��'��x9Z�J"`�zf+J��l���_n7kkMe\_��G������]I;�I��C4)S�\~E�M��('��bP�R*�7m$偠̪����N�s���nz1�|�Ѣ�}�j*���n~1�e�ҿ�Wc�@K�dfq,�ş�<0�;��z	��������D?�R~��b��zf�����3�V߱=o�@ �(U�
'@�@%���-w�	���9��u��d�;�����lʕɰ����3o�;���<g&c��L����<>EJ��7����R�MLߨ����-�Zq;��������5�ٛ�
]����wV���h ���
n7�,���`=�̤<���1��Q{�E��ZF���T�y�h�a�Q;�8�Q�3��o㘀/��37��M(2WP�\�Hd9_f2��S�f�G�h�T�?0p��#ޮ�mCN�P��w8g��#�A`lx�!w����B���[7�<���ޫ�Bض�)0��� !]�H̲h�y��}{�	̯�y��:#�=֠m=�}�>j�V X�b/����s��	�wi�9mdnl7��������*T6��_4�^���(ۧ]���	Z��I�`�8VT!���8-���lR�#bw6�ӛ�8��az$��L�잒x�`H���FT���C(��|D9�[k%�'	��C���7�0�h����|�^��	�o�$�@A�6� ���T��=������V;�*>���S�h���g�*Oz�,.-��َ����`�h�	٧�貅v�>nL-�goh�op�C�f R<c��j�H��_�*�4��IԾ�tR�h�JE'-�*��q�F*�lT�/R�a���ן�wC��� ��J���|�;pK75�;��L�g7�}���"����_0@7���
�L����RFſ>��@P\��Y�Y&���
o�
�6w��
!�a�I]0=����`i���0�/��v^(ʚ�)ɍ�K�{�;><O�]�o���<Vj�l�$�W�	��#D#�J�)K���V��N�$�XU��3KT���Y����UL(P<j�~���iG�}=��*^q����o����k���c������>h�T ���,����ifhUh�0"��:�I�!]6�8�q�`�5�P���1Z;h<+�4��	�/]G<���4�ʫ%v'D*g$Q�}nő���v{ە��EU�� l�5��u?�i�v-��ʙ��N�^ ���÷;��v�HBLw��p����ά�Q����z�}�u#C�ƶx��N@�F,��p���7&�+I��g�TXq6%�l#�?�׫!v��7��ox���v�d���AYTBMuB�`K�������":�&|TE�f���ޙKV=��wƏ���A0%tS�J���!y��8^H.��[�N������C?,xB�O�
wvz��&i���~Vc�wP ~���
����L !vZ,�Ж���"u=�Ǵ�p7�'5<Dx�*n��؜��s�Z����<����ǅ��\���W�O��K����ư�1J;X|,/3��{n���rh�?Ǩ����i�>	�y��<�8u��rS��k{)ʝ3�Oh�nԱj�o+i�W�lK� Ψ`%��0~��:�\�>E�s��72C!E��U�7���C��fO�h#Hj,���.)GSp�t{<>|���&�����|U�3:���dA���Nkr�MM�ܫ�Oǟ�e�m^\���7�n+�6�L�A�����jZC�\���+�ڱ˾�o���WgE�?��T�����q�q�#T��M}-U�w�FƋv�����u�y
�O�r�ez'fn=�,h��H���I$���>��g�xD4�	QuLbot"�&z����h�Y@5p �ì��w`:�f���H���e��ܑ��h�M�l�}�5���ٿ�-�����O��ػ�0��,U��]���P�S�:Q��vuW��:�Jm�xGbQA��`����J�C�/������	z��IY���^zsO�<� �7���_�Y(�Ln��'�����c���
$v�"������a�>L�\�<1�&V`G�ō^�M����G�z�i�u�p��vr��$ېt���
W�Bl�wA����Z�E��mk5�J%��6�DC��42Y�^��--��<�M��p�\�$9�iW?�յ����t��/�AC1�B�1��@�+2"aѽ�Ԃ�9�7��A8���as�4}Q��	���{�t��E��ʤ���a�)2���BF�h�K
Eb��u�[�D�u3�z䦧�/�2כ�2n/aq���2.��W�X����@�N�&:��4r�+x#1Y2��C��9��Й�8'�0�?ao���$���Z�K��Ќ�h��m�nꉴ�{���m`�o4�I���5`S���p����37u��O���9����af��)�����Y���p�v��f�U�����O����i��L�	�mQt �O��P�v=t�=�ҌNN�%uZxz8ω��>H���wڸW(�>�ŅDx�	Q��� S�߿o��;�*��Ң�7DT�[��gÐ;!���;��D���	������պ�,	�.�8�@?�����U��(4Z[�����l����}�.|`�v��@����p	m�!�Y���*К�,y 