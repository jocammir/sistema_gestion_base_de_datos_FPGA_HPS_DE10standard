��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��ᕫ��H��gq�f}���+����c��0�7�*�y�HXH�+��Y�Ar�#�<�k���bu�-��.���O�;����b���7pE+�������v@��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T幫$��7��`��$��l���MvZ2���"k��n�����ƚ�B�$GaY��5PFJ|T3�la c&�}`�Т�;��l�ݫ�F�.Jܩ�<�l��l�<�޿cJ؛FR���d�\Z�9NK#�Hj�#������H��(%`�Ǒ��T��:��&kd����'�'���V���
�z��Z��pGs(TS�e\���3�(�^UЏ�:�MS�|2ua9������������c.����]|��ާ�Ǖ4C�?ԠKS�:a� v�9oU����Zlxu�&E�\�Q���}���Ν�fS�#A�f*�
������l/^�//��D��_������>\���ɛ4e[_�n�Q5���YI�#9��٩ZZ:��#�kn��/���1Y�u�<f&�r#��/��}R~_���:��ܛ%��T,��9��zN���3h+�o��3d"j�Ym/�Do��)�A�p�Sy��}��-$��
���-9���ͪ���Q�&9i(�I��-���<�����=ox��m��ờR/R�K��%X����	�����wxv�]�\µ@OK�P�fFo��G4�l�g����<�� ����_lS@g�� �o��X����#עRQ��!��Ԣ/���yN�c�z�y��Z�"��{���[�x�nsg������b�H6%r9�"�8�w����*�[U|�T��k�����a�E��"� �F�/�ݛ��HSƢ�