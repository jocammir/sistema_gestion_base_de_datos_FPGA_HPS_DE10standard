��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0���p�?�gu:���@�6h� !�8��%cq�xQG��!ϙy-a���|�"���[AoH�r[س�[2W��o�\���]D�4�hwx&�Im����<�v�i�Ź��,�u���x���F�)��ƞ`�D�<�7�1j����I���C����M��<�4j���
��U�ɗ��Q�rA0ַ	�$ �:��h����3ۼ5��i��ӅD/I�͈ k @���ᐠ͝P4�ym�	̈́+�v�)`WF� "���j�4����=C)��q8%��Ջ�n�y�5��U�bz��kGG��b�2�&����C(�g4���ɝ ��wt��O��S���B��Z�p�³��OQ�@?}eq$�aB�*�� ��X���K �m  �BvET�^�}d�dA�!^��3���K>.n��f��!\�l��M�3�� �G ����%��kh͠U�Mq��v��Kl�eSd�7�
B?���K+yK
u� {�)�e`�B�{�����v��}�YXhw��͢�ȧ7o\)�g�6�r0�g/�����?1f����cw϶�O�ˑ��of��y(��&��
q&�&$U�z|ſ���ȘT��ܑ �SjҦ�8��K��#]1�}�M�[�V7]�᪤��s��͢6�;Ν�'�����5�(Q�?�H�@.#���P�uG�!h�)[�� �}���/�wm�Ф3k�T򶌈������G/���p�u�_� ���g2�^JC^ф(�N��U�a\�h��������?΢��e��؏��-�SdI6j]���3CbG�MG`h��,~��:4�XlH���Oi����r��������9K�`�����sQ}��8{��'����pn�D���vI�,�c
Oi�UC)"��by/�����8��5 OLwE��4@�:���N�FE�2_;X�*X����.��:�N�V��S���5���}2]�&T�|���}�r�s�%��ؾձ�A���֩p��/W�\���z����h���B���������?�O`�q�T`E�R!!S!�.e��&�A��8�K�$s�y�V��r���������p�����ao���Q_�)�%���Y��^{@��\����>��D��hߋrܧ��&#�*5"-w���+-%{ɸ�-*�@ݮ���Ao`�1�`lMeBoN�z��BPew"����ֻ@�L/���\�s��|6)]i|�s���U���+�ِ�9����۬����*�&��Ns\j`�A�3������2ŷ�&a��G�jb�7�o����� ����P(��r���2`� ��q=S
����
�Khe)o��е64�a�Y��*���Z\��_�G�;��pC����(��(ڙ$� ")���%��6����0O�Q�rc7]�V��V��HK1=��3�>�`2l�P%�w8�Y��,0��:����& z^Bv��`��K1<A��+���*�A*��h1����o�&;�)vNQ����|���
t"�ԉ��4`[�N��/+�-�<��SHڢ�����Ǟ?�ȓ�1��d�WwZ.�^ ��VL1If�#�񈠧|j�Z@%�(6]�.�E����t��t.��7<)�9��Z@\�`��@г����J ,+��i��Bc�)�H_:0�a-���¶k#�n�Y�ݔ�|6U�1p��A�B���]:)e(D��\�"G�1~�'�7���'IPR���n�N�f�����v�Z���a��Ul9eϚ'�y��� [��S4�N�|���p8�MGEEW#�4����1Po��6�,>�>�t��h��# ����F�_/���o�>nW|%�P����*Okr�B�D���A���4=���D��A�(�t�6׹\�۶H�3�D&�m�%����*�1ʶ5W��B5<d]�!����T�[}_�� �1ڴ%�8�=�i��u���ռXꋜ�>:�v�A>�=�˾�"�V1b�(ؖ-����=��K����g��y�����#�a�_�n�2뒄�*�ڇ�Z]�9��	^%q[,C��)aT�rOL�>f���t�<�/b��]�Yj�L�8�D��E�)��@>b@4|R�b���^����p��u��n�N%���>
ǳ��	�`�S� &�SK�1M�H�W���J�?�����~�@>����}��'�k�P����Kҫ�d��#3a��:���*n��I#��άL�6�_e&Ls���;�	dc�w+�/?�!�fo�<��K��/G:~R���g�1����߯�,�G4�2p4�^�;�ދr�x�\�0y_q�-5[y;ゾ��MGd�k)��B��q���O�0Y��%bn�������KF���H��OhR����������H�`����� ��%�D��x�-v�%8�W��.]�&[�UC��j��zt���[ؽM2�����+\?H��V梒s}�;H4&��؍�#����n�r"�o����="@�}�����V'󧎋�GkU4���ԇC(�����U.�t�a�l�p��vϨ�Lj���Td�
��Å'��<P~�*#H?<2�G&M�&75�>�U盺�������k)^�P���/�`��g4ø� ���+l���(����ڶ')9��b�#��8�i�Z��ɳ�8x+!n�u��O_T<K���	U|�6<c�z��o=c}s��!��n�}~�{����eV�o[s}�3Ҽ�ǡ����Q���ռ"��1'��M�jXR��������Ԕ���{�-�͖uJ����TL�H����E�O�0���8U�*�>XS89n�N�9�ݫi��G�2:&a���~��	s��oz���e���\y��lV�V�*��u���FC�������A�QS�j���hT*�Ez�d[�
�����R����:la]ǃ�-Ŀ���\�U�k?��<]��.@��q�c�y��]q�ߎx��J��e���߻��W�h�"��=p��	/,��z�z�I�X#uB��md_�y�\m���KP�g#���1��V����>T�����5f���V�<��_׶<<ʔ#��I�Q��\
C����}
E���t�@�b���k�<
KFY��q�fU�OG@�zV���e_� �]'9Z��ú�X:aO�gL�^�k؂�Ih�R�� �{�B$�O��7��8x��@� ؒ"��2�]� (M:�Z�I�n��8�d�X6Se�&ܮ�v���=2Ui��p�T!J� �h�2�'��a~������N%�%���*���'�c��@/�:��g������
i���!͓����k���(u !Ӽ��-�V����e���mAs��//�K�%�Zv�^��~Lf3���-�����C�噷�$�OXN��zX�i�9�)T ^QʢW� �z%%�!iz�v�3�4?1�7��=��)ag���CJ���by��
��Z��<�b�"��P��6O}�ޏp=�\{��~�$3�p�ӫ�UR8Ζ:th$4�2u9�r��������s�.�侴�k-�-j7��wC�E�xM��.��3��W�A�*\j��AJn"���s��܃��������0��փĢJ�h��C��	*�x9'=i��;��!��P�$١ FJ�D1R���PA\��8��N����N�lG�ⓤ���Hk��M���g��o4{+�n��d]� ���!�?��6#�rD�1R���\�o7����C)����C`mS `��ˎLɠ@<�0�8'�Ԯ��#Y=�p�|>j���T�U\G�Cy����?�XQ�y*����_�S�V`�r�P9}y�X��0���M�7h�ɞýD"Dž��h�n�5�q��˪Mm��`)�`D��YvJP�v=�k�GR��������g��]�M�B�1x7K��&c�ح鼒w����;oG�TGG1������_�v]�λ�8D�z�N���z<Vf��&J@�Q��0��C��N�)21����3�ijl��j#r���G�"�O�z^��B<*�W�dQ,��@�Q�}�a-Q�em!��Ţ[��l�" v�����.JϾ .>3�'I0��o|E�u����ь��i�g�Y�{�S���Q�d�L��
z䐥�Uw�KW�P���P�svR�Z�T�5��f�] =�Q��a7���Z��jwه�!B���6H��  �D���h��/���U�����Q�P��b��:��k_$K�A����M����]=���)�"��Ǯ�QE.�B̖I#��z����-	J��<�;�*�x:�m)4���x 9�K+ �ҫ���^��?�R���/���<�#�b�Η�eIl�t[O�W�<jSV-�<�H)՛�+�`,�Ye�k��Kk�Ld���h�����{6*� �5�5k�Ϥ�߽G�Ñ{�{���Z��Cs�_(�N��<t���&d���=��i��ɺEWp�l��Yi[g0=�I�JyUw��.i�|�!	�o�b�>r��a4W�s��\����ᳵ�|.�s"745���oI�M���{�4��"�
�3MZ��ᩗi.�����"�0�<e%+���i��>R��S���CS���+��ٔ��b�9�؏O�iv>2 g�'%�Y�mk�5f�-�<�'%��\�"-��1m��T�.0���ޫ�Q�,JS��V�K��@t������ɲ����@+jc�?	s+>N1�s�3މ��2���AȻ#.f-�9q��F��-��0��*���<�h����V����b���6�X��J#�_�%Zk�VL��<��>g��kb��ԛق���!��Tĕ7�d�����KT>as�^�l��a]�X�4g�I�o4�0� �5�����Pzs�\_�cS�?i\��i�g(�%�d� �,�8F�9<�'���>�h�������^��� ���GFHx����C�dM�e�`>�+ "�d��U����@�JO)�.|yB6��q�Y7+n9H�a�ڳ�)�ƉK����fȇ�[�3�V� n�n���Ɩ��t#�՝�c��i��A��,�jI(lps�qfc�]��,P��ٮ�^�ǐ}ڪ޼��Bb�z�&��=���L�Į  f�d��z$�@�w��~`a>�Drl6Ny
�ؼ�	�,�6i(z���bo�rY�%ѳj�cU�9Hݒ�RLin���� ��MV)S�E�A"��}J
�7/�:� KT�GB�K�E��Y.��ҚR�;,���FN"p|~O
�Pg�3�\*�0.ߺ�2�ϯ��[�~@�G"��&0��(UkjS�C}�긏ݠVܒ��C.bM�;�(/S�ki���vߡ-�>�&K?�(��hiSgBd���6��&��9���s�����6q4
0�\ u�c~oK�Tn<�&�ѧ3��ND�]��=���I
E�Eǯ�7�7\�1=څ�ցu�
+o����4�5 1^�[8=��88ϓ`��^Ue��G�heJ��qg�ZJ-���g.�P� P� �5�oM�m( �=�3��lo�.�PU���s�aR-�S�r,&��1�>W >�ӿ��+�rg��^�Y����<)��^>θT�� rl�@2=K\9s�A��!��f��/ݤ��`e�O���o���g�B@݆<��1�i�A�ԩ�����mڞt�d��5�%�$	ƲE�d*�sJ!T�JI���#H�'§2����ң0�<���z��;0��J��,�!���k�� P./�����?�a�3��e
A��R�z�U�Qc5��2��E�(\�1� K!o�����8�h��%�(8ڀ�8���;�
x��	+������Vzt��ᾓ�K��l�T[}h���԰�4�8�ٜ����g����o����
���R�Z+�����;3���#g"N>�ou��1�P,����;6z9��d�s�S����N�/gc,{�2�3�ӌ��$�戃Zpt�z���"�@�r�U,YΏ(T�n>)d]�Z;������{���x�/��P�o����C*qy�����v5��N(�R�]��+kt[_�'�Ɍ)3��?-|�v �l���۞�lEC�!��h�,�Q��G��*b�~�;�(vR"�I�wn���5�رX�_���W�L����/�q��� ;X��={ڊ��D���N����!��zO �LEc��A���o�bȄ�����0ʎ )�ą-۱���pH���p��P�@_/��Pk��Ra�1'�DT\C3���$0�D�����Pd6�c�eRI�Av��
�����d�Z F�%R����?2�L%�(�y�'0!+�I��&�H�҃D9uUEV����?�B��1x1�b?�	�O��]c��I�95���%�bKG���4�QJUjY��R��)����"�M�ܱ� ��t����NXm-k�v�O#��g3�a��A��Vs��攰��xB�zN�0���=}[�`���}���3
�mE0�^���`2��&us�S�2�vD����A�\�� ��ɫ}`�NI�G���c��|�y ��&2t�@�U�7jW��¤Jj�]ҧ���@i��ԈE���LN�ELm��hZ.M�ɽ��U��z���?E
�u'3ʒ?B.!gkBQ_G-�>�c;�����%p�����
r��Ǹ���Q��2g�m�ey�
5un�e�%��и��k���M�����@�3��m�]���A]!vX�R�:r$�'�6����
�Ο(���ښ�;���+[���.W�,�#�7����`+��,L�Cz��`9��?�Ո��\�I���JL���ӆl���$�g'��B;	����c���{�O�#fp�J�N�ZE���!����|@ŶVK���U��$��g9}>�#�exv�j�u�ｧ�����=��ٮ���x�>��$u$����q�<�T趗B�㉞=A�ƻ7�b�C%t�˓L��%{�#���e�����8��q֍{*m�����ZG�}�&�JN� 4���K���eG��"vG��1~iX�A�PxAe���⤦��a�
U�Јr�U��_W�@9��=�xsۭ�-؊I������=�<tI+&ic7�At����8ެ��m���"3�Y��ٚV�p�	�.1(�������}$�m�j�y3�j�yubD��wĨ��f�1cOmX'`�����|��Z1�4}�-�j��Hdf��3 �hD��(��yM�z'�0"���&�
�U̼�S�w�t��goUF	�j����l�3���W����>*���d���2y���q̢�*���x��Qa��+�!��k��!f,�qohS~jg�[�?n�h&��*}�X�&R���F_�C5*�����S�c
h�A�O�M��
I3�P��:�ӖD��	�� |%f��?t:܇H;���	d\�]`��p����ΰ'�|,�2���������yc�zt���Y��/�� ���;�i�K����L���Lk��<Xl�K�xx���e����J(�M��%4s=l^�eF�����R�FX	A��ǽ�لņcۭ�@M�&�m��\'��҄@�OG:�A�7�G�`u����Ħ}�_N�߅74$u{�f�����W�{���qtj��rr�):����+X�Y�Ւ��:vK~or2jt�+R�,�,�� �U�)�ƨ'�K�g����b`��e�A1Z%�����̷6@
c@��ú���<���u��㾉�]�`C����9�[6��)r3Ȼ���'�g'2�'��8e2��,��$�����Y�^_{�� (G�J���~}��:��4R�A8�[jD���a��e���uL�]��wN�3U�0����l����[d�~O~RҍҔS�=.��1�7��` ��S�E�[,���Kꤹ�z�G-@ӹ]{oPJ�Դc�� t��fT ���b���1�v\&��/�7ﾍ��%� ze^�g��S�l�ӂ�%�@^3�K�`]��ֆJ�;�_�e4���D�)����.*J���c�]�c�D{y�( ��)޻]�����V��q�����<����_��6���U}U�d�\��LC�����
ɲ���_Cg�_�H���HӍ�*��\�Ax9֎q�ԝ���=�-���B�r<j��w���
���������T��xM>Fg1�;��.���d{�q����6J��ww뙩���,�~?��}��.� Ď,���#-�֫�#̙�
�o/�KY"�FˠL��f���cv��z�(�{�Í��l&�G�(��q'��"����J���j�����-o0۲B��� �>d?|�����	ZS�B��Sz�fZ(bD�/ɱ5Fn�$���K~��+�b�W�m/�A4]r@��]]��K�p���\���a�H��M��6��uF|��ޑ�_F�����T�F&��5 +���v�h�!a&�B���@�hR�Ⲵ"�{�����9V��X�B�=%��F�#�C�+� �"��l�=�ވ��L�&7(��������n�c裎�a��؈��O_��H2O���ܸâk�k�c��#d�;����EZp[�7kp�G�Κi')i5�r<�]�)�$i��|Y�w�p����HZ�e��;uw���?�)߰���!b�Q<�����vm�]�8�2�Ko�	ʮ�(j����~'�+�#���c 3S1Z\��7��[���O���M����t���S���i��A:7^�Sp����s���i�P@�V�.�	sADk~1d��Iw�����Aķ&��t��L���l�@�;�AY��?��(�J�����9�2���*������d�@��DgS@׍l��ٳ����1Ӹ��aSE[�U+f�� F�u9�`����Yk���}��;�10���7���+�&+N}��ۂ:cR!��f$R�$�ȭo>u�1n�a���������1o�b>��f��c�I�:�X�����8����G��
�rB��WpjY�����1+����PK���ʳ�쭗����"�Ε��\�T�̦S���EDhp?mT�-�[�G�\I	L=R��$,Naя��H����u���\.�G���Nzc��6����X����z=NS%-ð쭻�9nA��8u�)��+�^ס:��)�f�d}��B�������ÆQ@��R��7p�]ugjY`j�H����|;��o�<k�����
���'a�5o��)�� ��ç��xg����L4��lT�a���l^����IW�)nA�*=��o�9�b���A��G��n�0��ӧ��N��$ftϪ���]�����o@l��zّ͔��Vž�EQ����=�@�k�q��|���g�҈�� ����kN�,�*���x�Mӥ?�i|Y�7>�
 ��1?����AR?���C�S��~��G�O�	Ӧ9�w~Vlt��v��[�#�j�^��{��C��(t�8�ƒ�+���3���{��,]3�ƙ�Hޛz����֯Wbk���X���z�$��!����i.�Ln셈g�T���`/�[l���~`�c�k���4�<{��x]���y�l���� �.;XĘ����"��y���{����4�ٜ0���/[q*'5���p���v�+�A���F'�=e�!yf��P��20���Qd�{�����/�~t�fq'f�&]�^@pM�vP������r���#��u"i��h0�.��(:KCd{a�s��=�Ket��V��m�x����!��{��AT,Hn��t�؃&�_���}���)�ʽ%�E�B��0�?S�BQ�w���6�����b�����_�5�����&f�z2�֟��<4�[�rUI�F6j��Sa�D�/�׷.���׈�K�*�1���eL���
c���z�F�p|d1�\qH�_�t��ņ`n�}��Y�S?ϵ;�_�eG���U���X�! ~��[j�	�5<w>��1�:��㢯�rqq��w��P @�2q���Q�)�k�]"�œ�P�>ؘu#�Afg�SЃ+����1��?֮>�i�dmg��W�}(��t'�P�����!�˙>sg5U���\X�"*�yi�S6��%G���؋<��+�Ϯa��<�hѳ��\�$�y�[۝!]��*},��%�����8�@\�2�w�^������^F������A��\:��:�S��>��V�`����ٖ���hp����x�'���b��.P!@�-�C�5(��YT�p�����C�gf.@B-�p��/5\�5|I3��[J��"_�ze����}�F�h'D�h�,��b�]Cך"x�j�F�V��m�פ��Z�*��F�
�E��ȀZ��Ȼ�B$�ĀJ�NO���Ǩ���i�n�_7����*�9��g<f��6�,�?�jhxǔ������-5��������TZ��  ���l�r:�-��i׋�uwI`A1\~�ndc���-�L�-;Kl;"Lf�x	�8�B��Ȋ�se Ꭳn�Uc���Tf��~��PsV�Ä���E��s�4�5P��;�"Z��-z#��)w��D��87	��bH"a�zzu�Ct�*x�%E>5M�
vy6�Y�>t)�(ʈ��@o���A�F.1W\!��H>ъ�Q���9 JcL�}�2_�,���BY�����Ӭ:oc ���2��N�]
��(zzZ�0"G�o�>�ZU�����ļڰ8�X/ݐAr
�&�0d�D g�q�V����߀��Ғ�"R��7yD~��3FQ)�8+�W���"��eS����Μa!��O�"v��~���A��
����ݤ�H�6J  *+�X���r@�=0Wd��6�J"2*��/�B��7x0���k;�G�ʥ:w�Rm���b��T�9��E�)�u&�5�~{��`4 �S`�˺��k�!p�%���7N���?磳A+]�-X����
���X�e_��/NV�t��"q�5S�1@7��ݏ�eӾ��ً��Lޤz[�~�݉1�+a 3�X�!����S�9�a��Uq�p��$�\��<M��Ť��2���Ӽ�> y}�׮O�Pi�]T|������|��}af�}}��o��_n.�]���=%�
^���EeRq�>�H��ɔ�O�a׍Y��Rw�}(�'������図�;�EsSbc������`8���πPȟ���׬�bDV��~{A̱$zht<-M	;s�m��|��	w�S�d��3m�/�x� �`��#�\��� (L����,����#���k��>I}D�t�W�.��0����c��W3�L
}dOື?�5p�(�9YCN�p�$A�0o<8>^�d�YV��D�e@q����š!\"~�杘��@y������&�#0O��Ҫ<�+�> ����Jn�����.�4ЛFT�E���*;>�[v�W�<}-��i� ]MOe���*7�l0b1�\�R���}b������N�P��5�5s��m� �Ϝ�2���	F��1}=��g���m0/��D}��u��-����ޠ(��)�K��5%}�@�v}��^?E�?��R��VE�l��a{#]�{P:0 F/�ٛ��%ޥ!OK���z�6�0��:�Y�D�m1���P��#�]3"��*W�϶��n��u��.���خ����� �lßX��8%��Mir<r�N�ș�|} u� /���iv��丶��}���ע�u��Þ���p�Za�D���lY$ܐ8Y���H����X���.�nH
�	H����$[P#ҳˢ.��\5���Ϊ[�ɥQۥ	gN12�N������Wc��xt4�`B���S/�Eڕ<���}h�����Agz��������]�����BeB/�����
�e�t^�Օؘ��)�}ZeF�+�;rW-��y7�}���C ������I׏$	��=4EșY[R��N�j��)��7暈t���b�+,���8���l����`-#1�ϕ'���t�|�%�E�e1x�U%rE,	�Rr7�w�j�{k���@�+�JY���}p"=}~�lAF��|���:�Vm� aūy�=��IQ!�Pw"�[X�t�Y�)�����~�Y�Fg!��^�0�R�4<�`��Rw��e)>RUGM��U��O~?3�PL��	�r��K	��T��h��d�%e8���W��fvI�:�"@#�d���Z�v���	�֜oש؄9�\��	|�@�v!���Ŏ8̺������S�p��s���.��z���E�!��� N7G6ܶͼs̚��8Q�`��QG�[)���>8W63��;>]���J����b�6m���z/岐�p�;āe����[��J�����5 4���%��&z�
s�$�A���U@��'��(�Gg#=�ϼ���{Y�@���-�VbA8��e.sf	i]�xN��ǿ�C�(Np�т��S��˶@Af]�<�m Sh�S�����s��y)���ā�z��G*2S8�=�#�t|�]Lw~%&��h7i�K!�O^Q�d�=��ߠ�����	�ډu��?1�BA��ĳ�>jg�V_?�n��H
�����$�׮O�h/��j�"V����]����Z��jBG}�I��+4Fe�>�H��J2,�IVҥ��sh�Oi���A��Ψt/)|P��H]��_K%IP١�7%�~#*�BB����d�r&�9�A��9m�����*-����&�IB�nMS�!2��@�Y2�����������m��N�r�5JGK7��9SG.�)�y)8�yBJ�8c�ͅ�xbԋ�� r����͖���4�Ձ�.i$b�h�����S�=9%����s�kg�nv�c8��!�B���m�q-�;��vl6�/H�Nn�Kܒg�n�'�e�k&3�򝿫�e�OO���xi~c[�nr��@��> ���ݚXצ���˸U�������:�����9m���L����0�2�-��1~.�_`��2J����y���t�f�8\N����Zκ9� ���0��ƣ*,�_並&����`�WoR�Κ�O$������[����h�ltXTهN�?� n��X}�]���'�5~�Ck�����w�9m4.�_�x&���z�υ������c���F X�_Gt����2����ȵ�h'd����=:�i�vL�B{�"�Z�FCc��:%�����ֻ��.�2�%U��:����u1O���Z��Z�K�P���H�����5ZGsTL��F*������ɳ��'lp �v}Sd�����һ��;�E9��� ټ߹��o�N��N���"Q�[[�xTzԚM���4��,�`8G,f����"C��)��<���5%P����h;�����c���Zߡ����O�NX!ג �ay��̖��^E($d�|]Ѧ���U�!�����|�Y���&����ә�(
��Yv|���?pltQ��5�]�����ej9q"�∨>�uu�hR���.l5�3%4�P� 1����20j�Pv��W���QV��:@��ϳ�?p2��%ܐ��jr�$f @fNy��$8�h���[AVI��l��w�̛�pœ�3���#y�������������Nk���ȍ�G$���m���Y�]���8^(,|ez���ޟ��}���zzW�`5h��]Â�ٍ��	�Jzj���ӝsk��ڰ2M{�G���zo}�r���dkR��U��IN�ؑ��8\\UӬ�cK�����HkAOs�	ɵI�ğ�bͤ���PI�nVt��g�gMM�P�e�)��ߥ2��e4�e��=�)�k�L(E� '���[bރ�)�N���js�EQ�J�u�28�����?�Db�1�3��j;��Y`�����}��>��8�0���e���A'f�:U��ͯ!�`^��4��N8Ă�`�b#)�"�U30V��;hD�,�_�ݸP:��bt����aә�$M�ս�5!� Vsf���g��j��v��䧡�^%����� ��CR��P�H�P��|k�Hq%��*�z�h?��r�n�#����� 핁cc>w�ߠ�,�^[��*9 �$�J2J�W?��uD�����ц{���u喔1\�I�uɜ�ߝR��*����[*q �P��\	~����0��]��S�r@�U� ��K�l���p�2��3|����h��AT�ҿ��"_z�Sl���C��p�zN�T�1�}�5����xp���R$�Р�����6�|[��d�<{����l�]���-c��R�N�̳]�b�/텥-O���V�ÊB����o�E� ��~][y{��/dcO!����HM8��Ϟ�zE�YI�cg�F�<�vg�#v$�K{�D�Z��t��z�Oa�B״�M����j(y���6�jt�V3D�0��l�A"k-�mb���}x��[�,"g�m���Uxm="�_�*o9n�Cn"�0>�hz�7r;�har�<�n��|ߤ�K쐡4�R�ш�В��.,��͈���zW�	?��&9��X/[)�DN��.�g�hY���H���g�t�-%�\JOe���ʖh�2S��ǣ.��q�9����wb��Ɣ�ྔ^�ط��L/$\Pf�c�7��{�n�b�JqU��Z�X�N5�Q��W@�����������"4pd�����2=��א|��YG���9R���R��#\]��
˥�����CT�C��5�%��C��[L�s���d��},�!��("ě�G1����Y�	B�#0��"�t[K��O.9�/��q���/N����蠁AOH�} 3�<Ƙ��������H'l�_eͻVxX1?^{��_��k�������1��y�m���u%�6�۽��h9M�m��o	���P�Zi㹁p��<B��["u�C�m	�F�.�EG�����7��E�J�;��D��_��5� 81ڳ&�"��.[nlw��u�:�o���p���*��'(�j��6�\�k�Io_`2�K�Ě�L�̳x�wr.�@��'��%�5�՜}Ҧ7�	�B�. lﰨ�l�٥�Z����O��������5��G�Lr��Ui��z\�J�v���]�ܯ�P����q3<? �IO��g{�A�܅�Nv�y2�|���O��m��zwMW�X|(���iƔ�I�Ř�gS&B�6��(!x��U5��6;����Ǧ+��"���'&��`�n;��A���ل"C�x4�kc��݄gLwa�ܽ�{�dQ�{�Ju��}�oA��%,ӗ�HaMV���~��o��t<�Vt����_!f��@�1ΖC���@J���Q�ш��Oi�s��A��n4���Б�>8�u�W�hU�U.J�-�Ȱ��̼|7	�@E}��XYrA5������Y�0�!�_
��CL�|�="���7D�n���Y�o���P�(�a��#�9���A���6L���,s�T���ttEl
�<�V�����T���*+�$$�2��6���ف9�ZC9�R䊝baE}��=悆eߙP�!�>7���@���ء���xu;�]E�웭��i4P�����q/���c��~8����ym��}��+Y*���P[��к�y)�}�`l��#��E�Ƿ�g)1��
N�Q�����/v�e�L�c\<d��)�6v�|�"� z�<힩��l�ķ��I���@�,����X�5=�k�>��mE��y,��˷l��X����)]Ħ j5z���)]���o9�������H�u�m�&]E� W!��Vc����r��x�
�8���H���%�R��cX�K������/�\}����4i�9�����<���K�O����ه������,��~��a���Ǖ��2�?�J���UuS�ϋջVБ���"z�h`�a.>E��;�a:���ù�r�}O5������#��8�%M��X��~.��s��>,�۩��AmC�s��m�iD��k���^]���
�}�6@��@ v��p0s��������jG;�5��#zW�����Yy��ըV�UM�qP����	z[W툹�_&�p;�e��*?�	j6��0�S�qs5㱏�$�JL��/��;#�\����v�����l5\~.7�d{��/9"~����	OSм��'B��.�=1�]?�۱E���]L`�^��}ݑ�W�#�����f�d�l7����s�S��'��\���)_�N�(_|4�:���'=�h��S�u7K�S?�����i�uh�3j�ҬH�ɲ�_D���� �i9*���oj�X�w��;=���X��X�J���s��Y�\�2���;"u��"拧+����^|�z�\e����5$����@�q�sM}����B}K���Rhp�`�Ay��y�!_�����w�qx�Y?M�,�	��
WL6�7JI.S� �h����� �͒������ \0��5b�!?;�߃uH#�E�J�����]�Z�f1���;���������+$�D�+�f�}6�i����UVȍ��#��{$@�c^u�'7ڧ2QjRi3+p�9@�:�o��8������m�H���R��M}$�gq�6
(�(/1\��ᴦ�5X R�j�� �)��g�ǖ@�0�/� ���5�U/	ap�+k�wf�u�S�a]�}��S���Q��UE.;�3+Jݦ|.�,:W�9O؀�D����jZQC���m���#���ԥ�F*a�ޥ���/���� ��s]�5�T�P�ғF�o�%#~���F*i�a�����x��SB��1 ����-T	��"���H֣��Z/�"q��(��4�t�N�����}H7};�g�GQ3��N:�/9E#��A���3א�=i�(�L���JoQ�
tƮO��+
C8�'�[� z�r��SV��@��1�a�p��B���I'C���n�$��)�]�����^�/���9�M��V$z
���
�%G��ӊ�MܒN"��K�+�ԕ����7_ń^mCn���;��q+����?F�:�L	�h��)e׻��uh�<{tor�Z����Ew=�A-l>1zn�?-���EC��Mx��/cS*�E�8����,�B�U�6�L���˖6�䲴=��ln|��zβ �K�O~Z�S�O��Gꑣ�c�':��1i�&8(,�84�Y�O� �P��&���'l��t��l��1��go1w]W���w��oDBi�F�
{�u!�Ng���O�~�F|��ȍ�ȼ�4朽��]]{������ð��&��<&�~����
�-y;��P/�ú���ƚx�B���󎑉�U����6I�H�����(m������,�و�m_�\��?v���vw��>XK7�-��Z5��-)��	��̽��ݻ6*������/����ɗs%%2c����׊� V��M����}%6��<�f����L(��n��ڑ;��U~uD,]���A�Q3��*�X�O�5E�Ga����Ӫ#L�5�܈�C��Kv�Qv�}V��+�^(2�Z����?4�V�v�wg. ���Ux~�P�QF���=����*R�i��SS��烔���!����܃�u��bё�QI�'�L���=���T�9X,N���������@ȝ�aD�*�X>�@z.�"&���⇬�4�"�ƦϒQ�lz����@!�el�M��Z�0�F�DHw	a�7{�j�=�H���u��7�K�1�X{&ݝP�K����$��&BёF��k�Ҏ�	��e�wn��hp�����0^��}���[���kO�H�UM��w��\����zg	Iľ?������g�x���~hR��R��~��'ӭ�!�{���0���1��\������G+�*��2�C��t�RB2�v�^�8L�����0I���t�+:lZ�:��g����+��}C�?k�H����j#�.U�&�ëu1�3����%�.�oǶQ:5��qpHħ�nj~�Ȥ!
,6��BD�o��P��K�����㛺D�I��|dLb�AG�D�s��+�,�䡴�������-��{,ךeo_*���,�ʒ���FEPq�y�AX��v��V�����rcM�Z�N�:���r������5�{|d�+p ^v���+U��X-];H.���r~N�ޗ����*����4��eQZ��V�!����*뜋��f+;_WZ�-��&d���Pm�ɇZ�����ws�	���f�&H���]R����f�\��p�%q	�J�$�I���򢿟�����z0M�����?J��I�f�}"�k;';qƜ����wq=����E�\����W���mqѫ�"8�ϓM*�-�?�3�����X�̖�SȦTv��P/�*��<��8���;f�s>��;���L�[]������o;"�h��ݙ������/���bN�V�붚��Fǧ�e4�7&u��& �,�}m�$+`�4<ޝ���ޤ0
� d�'�J`����n6U*�֮Jw��J�7��� �j��³�h4hJ��x_��]�A�zV���kRm�_��!����0�2fX�u���9�'�m��	�}��YE�R�6z�z��7��J���M\���J�Hc�@uZ��bV+Ԥ�`��ǭO���0�1��}���H��[X.h���g-课N(�HB��x�B�m2�Ee)���c�7�Re�Z3G��#��ԏ���,�e� ����h��}�$�`n��[�"*��d���h��iW�����bH�x���j�A��lb��{Kb#0��H~5��n�����u�����+kY��1x�)~� =	�~��Ǡ!�@QV��hO��yEp�`׊���ǫ����FY��g�+��$eV	�`Hob�K`�T�wH�L<pS�i5|��6T���x�?"�^]:�q$����9tM�ҕ�Z��p%���"w떽�n�oy��q!N� wI�l��)z�_1������h�Țx�k�,�q��pLp�u�����9�O�5��,��B��h��p�#����a�����ɶ4s~U�8`�zw9Hv_���<`�%�U��Qs�7}o��O`M3���<\���w)�� ��="~m���78t�[.5E�M"��ҽ &i��x�i�L]�k��6���������x�%���I
W�ml�]���xj�Z�6En~��B��U��O��陸*yd�Tg
4k�JU�jf|����=���dFM3bM��ǫ�p�s�h6Ȅx����q=�E�^�������F
t���|3���>�`��̦�E,��L�R��h;���Cc�XIh�6�˺��ɓ�@������l��$������@y��
fc�� �u�-07�@�3v���+��9�x���=EY��%IkI��m��ѕ��Q�`/�^�R�`��.���0�9]��<�
ժ�#3:��(zi�8˵xJ�y�ؠ�_g��������UM� 3�5�98W�ǲ�!0�W��DU�<r��0�W���q���cjf��$*�/<��.V.`�z~�(Y��
�e"*�VݓI���)0%�	��(�/#�Ue�V�'�VU�o>��L\�:�B�:�(M5��(M]��.����>,M�Yn�!Q�Ϗ���EA-r����t�ir���2-���$+3�;3%��0����@в�Xx�R,n�*�~L�S�� �����
� ��u9��kHP'iꚕ?�@z��q�4�ihdm9>�oO��ff�Qt��;�`�;��� 0�������kD��R�Wƴ�E��ٶ����v҇	[��ۻ�������}�G(���	��-����m�2sii,aɱ�	���M�,w�W���Y���4˰c��ꍬD��B�)/Xق/�a�q����
[�d
XO3�@���Q��M�_��ui�&�yf�d�`����GE�BoR��Ǖ  Ƕ1�s1�R;a�ǘ5����U�(Bt��C�ц����a|�����]��G�G�~g����T�Ϡ(�3
k~3�l�Dߔ��I�H��
��t�D@�j�ǲ�Jh\�C�1��6ش�pO������3��9[78�P�7!=����(/銩Tf׬۝(N궦hD=��h�<Z1���� wR1�kD�TD���@�?-�|
��^N���i�0����A�6��;j��y�_����� H\1Ь��[ےg:�wciy�E]�����2�"��X�V/�&)����S�D�;�ѽ7g��{Cm��9�ի�'gH�J���vI��
���܅cg�c���d��a+I�!����6j��¸珬���I(d���"�P�(�,����O���8}ǥ�#���R{~�����~��� H`zv����z�)?��2 V�xa���wf�0C�<��{�%��	�*�]��a������"�HC]GW��zs�9i��P�<H�SQ�F�Kz{���خ���� F<Ґ����,�/�◈]��>L������|'��1��]�},v��O��DC�ƌ$�6�]6�됉�w �ד��qU�vTZ��Gt��Ĳ+� ��~��㱍�W%Є�i-����N�U�d�b��;�H���i&;T�^�J$�q��{.G|� ob��-���B�;W,��h�T��E�E�2���`<	]1P�Е$�;�Y`�ị�7��5m&s�8Wz���Anq;�#2[+Z�M���2�sK{�4V����`zC�Z�ky��]�Ь�I���[��Z8�Q�/#��ak��x����T�����߰�,�����_3I~��������j�mӪ$�S���;�P��-�J��|E7Pƌ��8�,�Դ��:�\������},I�0�����47�P�}i/����"НkE�~1����� d;]��>���ʇ�M{�~�VU��c�sS�?}u��K� ��>P�*&b��C�y�t�L��}_$�b��n����!Z �������P�ߧ��%���x	�����u�*����c]lWmO̝�vO<Q���B0`h�(�S�R�y��L<:$f$jG���$��^ ���-:�=�;	0�d[�a�b��6����I(�Z93���n}-�!|H��5l�#m������g��Å- �RG/~f��� l6p&Q )p�pVn7沟�"�a,&*�څ^�9c�r[xt��	[m���&�M��o�=..B�Lj>�8��I�?�5��=�6/�,K��H���p��_�н/���h]��k��Pf#����b}e�l��f�sF�N���m��R7��EC/�����fy�4#Bu��w{�D�r��THl紞{f>�К]���<d�&�a⚷�q���Nm��0+]Wۥ�'�:���tPs>M�9L�r*���7�4��J��T�;:=�e��8.���<\1��b|���C���b�.yk��r$��<#<z���J(�xGI idA=({�	�] ��Ug\a��[�*�����EI���@�#����]M�f�c�7�:Z�}�5��̲W��pƻ�'�4_AsS���	�kw@�}T@�%�-	�o�<�!LS�D���z��}um��J<|G���ǋҷv�yP���?�lP�8\-��'$��vSÉP��7޲gd∎GE-����n�C�[jP�j&e�L����3�ְ�߅�'I�Cm�}�����P���Ϩw��G����q��G�L�Q������ ����{�u�[���ƕ�;���_=�,ڛ��ό2�ba*�q���.���9��}$���A�+4�QF�j�������
}P�!�cIsa�Z�R��X-"*U\�*ō��B}���:�"�����N�_S��{�5��.k��X�����w\�8H���E��>h����52�D���ı���
Zޅ8�#g��Ļ���i1cy�Or ���]�<4=�)Fu�m�O�=�jN;�ٲ�Q���8���;:� ��K����vR�csi�<�,��#�$���T�>?-\�o��C��g�Er�K�5R�>�8����dYTG��a���{��B]��U[��w ?�Q|-�m�R�vŸf��x\�P�H�iY���G��mA�<x��?)ZH�a�N��)w]��+��Լwf�_��������W�v��O�$��:ˋ\��im�7�r�N��BR&k���&\��Vom�T͸h�[�Ey�|���b��v(�'�K��$E�gH��.�zI(�PM�\#8i��
7����j�� k���W��j
��~y<�lk�LK塛������m����zr�\��H�F�u�<� T�u�dl�!ސ�z�i��6�X�x��\��N}�		4˓?:���,��1�/F�PUOl��?��*��GIG$�t����e�yٛ�qf�7m�$-�=������$-J�wDR�UH��yCw��?��KW���Ck��m$�=Ƀ%R�}�y�)��y]h�r_�gN�e��>��[��	������ޗA���=��.�;�s0J�-�?bsDR�~:�g4��IqKJ���� ���S��F/a�/�,uF4���8�:~{������ �����a��8f*����N���b8���'OY�{}�R��\RQl+{���	�y�r��������ҷD� I:/�g�$]��� RM���r&�_�ѫ
�|�8�!�k\��\��0M�-�k�S�Z����y���mo��騿�<��=W0zT��ҕSaZz\��P��?����k��l�>�ϛ�4�Q���-!	f��?���I5��M۝�azuZI]��>	���rt��|�q�"�'�P�i�ȚB�S%'���Nn�O<?^�lOE��
��� �G@���f�F8��8BM��^m��7V��gܾ��D?���?]�bV�>:[�\ڊ�)	+�E,V��.���2�t�������ފߑ#���[�U���}���Y����S�B���1/P�)'���T´Nw�3�.���Lq?�al�Qs���ʅ�^����C����|v��;ݕ���*�� R%����5�+u����,�z|aw�	�K�Z�`��U�&���@�b2	�ݜ:2����x_U���`Q���Б�E�[���.哌�x��+ G��=G3��!���>��Сu�ذ���>�OT\g�+�wrD6.�]���k�� S�:Oo-��l��}�� �Ӆ��R�WOV%���0����i�*���D>��嗞r�����bw�������K#�k����o�.l���� p��~���*w6�լx@�ńs\��Ji�Q�N8n��h �6�Y��S�z-&����	�\�;
���i��o
��7�p��4|�,���[NYfy�z�|��[0�&�ʠkd-<��w]�o��\�rK���(O2�S���|[Q����_טM���'0��=�FkX=Z�or�	<�-���_B�\����3�ʩ�ibC=�*���I5&>:\c��S&ߠ���1%dlk���\����0��j@B�
h��=��r�'�:���l�X4��¶������VD��Z'v�N_M�5�}��=�n�3�@C6�*�����}�0��9����#��q.R$�u%
�sv��-~l�w�5#@N���Z"l՝�@�(��+�9SI`ݛOa��9]����HT$Q�hP�D��7cf^׼��/�����H@����ks�@��<�KZ����M���!�����CJ��x�Z�� ��?�`SƩ�k
c�w�yw	�[i9G�dc#�H+�J���nx꬐�u`]O6���v���"�x�p1��\�N��:�~w�B���Kx,x�b(���"���JN���@9�u:���"��`nϞx���^���1ۂ�F����J� �.�~�����E�>���LY?�4V���,�ր�Cg���:�V<]�N��%oW� 9V���쟆��'��wЊ�F���O�y�4d�Y%��n�R<��5��qԖey,�@���4uO� �����<H\��'K��~��Τ����	Ϛa�\ 1r������Ş4����v��*E��\l:��#��< �/�U&�t�+����LC�(]�����E���[�M��<�FBΦY�@�������A�Y�rw���з��,O*��������"�`��f��!�X���E��"��w!k�@�v���E~J����	�lٯ�TdZ���3K�K��1g6E/	5����6���n�K�cs�������J@�R�A4�|�$�f*��X켍�fQH&>+�'�@�����l�VN��!+UϾ7��N��H�;�:�n?���Zy`����eݼ��tB���ָ�ELV���K��g�z~����ƫ��T������G\x�a�z�?�D��.q�Wܴ�!�. �	*�H�7Н��J@.��,��<lT!�[��[E�6�g҄Vu����Mۋ)6O3��1�J�:�
r��la�d�5�̄���=G����~���֊�R�7d�Z���Zr)QrC�k����]��$�f��C�dX��涤���h;��Ch8�6�_� �}�!��NC���Wf����� �P�u�k��"�`&Y��g����?�[� ��I��5��� ���^w2d(�Gm4�)(o�����M�=�B߷I�|sC����/�@{�6��J�=�Eɳ�D�4��g�_*��Sǣ�!N��!l_�XO�m��~�k��v'�
�����Hx��}�@��<c'���2m��b3m]����sJE��-��à��X�E<�E�R2ҵO^�Z;ԷKʛ��+�킚�d�>DВ���1g�rвs�/y�
v��7���ˀ�*�̰�%��j�I��^aj�;���әv��D�h}�Ԑ��T=�����V��4+�>���[Q-��^�]4d�W�O�ې������b��Q3(�c�ƒ��$�v��F��Pwe�i����X�P��)��|��tt��\?5����g�>W�P��0���I�#z�г�Mb.$�w��Ρ*��wV�Kf~�4�깹7��˪�9�9��+�<c�˨\Y�ܪ��mgl;{T3���Gh�z42��A����M���s痬�4i�紊$���=CBt̨���6߭� �ೳ�Q�r4����l�D������i�{I�/<D�p�"�0-7��@T{�s0��z��x?�.�د���[H�K�aQ�}҇@ø갴$�6:������x42n��Y�ǫ׷��w��,P�C\VÚL����Ln����F���;�v�`S�f[���4Q2K����n*?�G`�#�����.׫��*��4fS(p�ߚP��#7x�x�f�.�/#6��I�Z_9��R�{Hu��-��W��%墪Y�[Rzy���P[6�ɰ6��2���ւadz��o݇�P7gK��X���π2EK��Z���g�Y��5
�Pi�	T���&ǹvI��m6�����Ty��y%�T��^�j�C.O��s�t���y�z介z�~wF�RZ�Ö-���	ɇS�̼�����f24���T��`�f�h��9R�V����JA;h"�x�!��ԛVÚ��h,�Z`��M���s�4Unr�x-�vK���ɴ,;�6�d6 �Z��{����:K�l�6p!
�+#]K�	V����������˱7�Y�m�v���t� ,u�����6{>�V��aL�`���=,ʌ8�k������qT�܍$C���Dq��..�$_�Z��7�i���\.�D��G9[����7W��׈��%%wQ���"?���/�T���3{Q������(�v�kvQ�*Y��>�?��>�+� �<mӣ��m�i���Ė#��v�♔�wk�GEq�꩜���\�G�鴎0jgb���Ӽ�B�2�LR>��e��]7k�9C���۹E���1!�<�kY��J��/�,kU�A0�{�7�{� "l��'+0�6+�l����>Z&߆�}C9�Eu唧f> Y��58~K|gt'N+��9�g�i=��܋�tg���86/�xrX�
և�V�d8� ƘL�V�ߋ���j�(�ɼ\E���KC���\�qê�/3,�To㲈z(�o�Ƅi���C�h��E�"`(���T�7��-��k8G\O[-=TP{+�!1�ρ���r��H
A"yB��.o�nU��=JS�m:=�$97��k^W�멵<i|kh�6��v��L�}�
�¦�oܵK!Io��1C�K����(�����lŝ�b|��^ސF~���:l5�$Ȇ�:��0]ɴh$�TQ���(e��s9�6Ȉt�anRn��"C�^�U�H�Ζɭu��C;��Ē�^ݝ�C|X��1	���C�?�%�.ח�95KR��F�[ow_&���2�$o_ ŗP�J�����o��`�2O��t�h�G�ll���5Lw��4���Kn���K�,Vg�@\W�/Z�4(���_�x��%T�>������ <D*f�WqOҙ!���<�d�3�u	P���+�w����yD��	׃�y�����ص7�R��"��a�����#�AN�@3���!�v��J0f
���S���*moiA�s;3QN�ѫ~��k5����:J�.�o�!�#@Į�,ͥ4)aE���!].ep��t��npkF�8)�ε���fT��m#A���L��L!��O�x�S�,44�	o� ,����M�|��X����k�M��tt�`�hɆ�z��JE�|\q�>h������M�V6��N�`q��=�@�q�d�
m�Ā6�mőx��q��cV�hp�����C�j����U[�݋�,؀<��[xg���Z�Q���!���<Kj�.�<�ȕ��ɡ�ˤB-%�FoʛHy�	�ۢӢ2.t�p��� ��[@�P�Z���? N�	b��a��$���>�ӒE����k �)�9`�-u�G]���Y�P�����<6ŤP}S�1?��3�ɇ=�X�������2���7D�HD+22 ��a[�-��U�9�uƌ����}Q��x�9Y�	܆�P��!�Ry���PE�QK�b�� I��i,%_L�?ތ!5�\�՞f�եrw��&��!W/bR�p�d��<�+J������g�2���R0E�.?ʬ���!�v8�n�_j�`��1�3��1&N͙���1JF�pZ
C�N	��/sRA@+c��y�^�-Dau(�>3W��e�P-�7d������4�!�3LK��t�,(��@<u�ը)w:�F6� �CÑ��K<`��*�x|8�ҵ�]��fVV��A�JB�}�Wyo�D��P�IOC㐓���8�h�;ż�g�t�8�����dJ�W�Ck]��j�	эDҾ�-R��N��ϸ�V[�����K�̟�¡�U�G�Tu���o�Q�����.�\��=����9�".�����b��Hy�s(�ૐ*�)�8�%�o���*�����Vq#gQЅ>�R!.<��}?U��'������2+�׻�����O~;�m- �~m��i\�J�����Kt-���(�[iEf���:IQ�~��b �q�F�E�U�^c����/Z���}��V�&�I%�����XE��-4z~
�$�uQ��]/"A�=iʾV��_"�*�Rڙ�����<X�uv��a>��=R���"X���6E�l�]�Ĵ����3`Qв5���(ᗝY�����7�������؊���Yv*?P��?E�eW�CX�b��Eo	�j��p7���n�r��<f�vP�WlƠv�������K!d?)��O�F;~� ��~XVC:�Ϲ�
������$k���>D )���Ɲ֏��J�I��]4�"	�7)ŵ?�k4��	�w��7�l>k�X���}'�T����o��6��.�$����+�A %��jB���&Z�d}Eq�֋zCZE�X��4��9YyjPU��G�����d�%î~]�h2�T�WbU�/��D�G�^B�����ԉ{����Ә@eX�q9�2�g�vYLz�PL���DZh#
o�d��C�D�F���)zgˊ�|.hF�x!�o������@�2�+3E`�Z��dwi(+�:�c�i�46^3c�aw1rN�!�ނ1�g�,X�,�D�%�S�/�b?��m��3�he/S,^l`,[��(����Q���/ ��D����sBh�X9y��j�1�#ύ'�T�'v�nKNS�I���{$����Wx�s�a�#���;ҹTX�SlhJ/���8���� ���R8�,'�X�SK��In���Eor�x��q��˻�m�}�Jhc����QP�hE_c��mֽ�L��ld�� ��~�}6ZY�ߠ�s�:�p�ߒT9���xȜ�2�H��|N�}��ʌ�?0o���h��R�WG�{{�8�	��L��(�����rw���h^Q 5Ü��l����f�a��֡��J��g�����Ty��gS|T���7.5��N��`�2��s����E�K|-a����	��3(8�}c&��x��>�B��
����
�8v�K��XvN;�GM��%�����`չ�)�z����ςv$)�z��`+�6�0e���t6	Ь�p�x*It%�ѯ�`th�h�]X�	+���K�{D%�����u�Rk6�	O� �~&��<�rv� @��eej�i�`'Rn_@�s)e����$���@��l-�\�C�� �����S�CڮA�2��
����8��sfv��1b���1H��?�X�z�{���{.\ǫG����g��v��Mx#��y��~,�I"�\8�c�ԋ���[���g`$�c�����ʼ�t�Bji��w�t�z��u�-!Y�׶��EyU%]?Rɴ1W掣:a�͝P���}!���S��P�7�U�o��<5:c���#�{�T�v��.��~w�H��X���ٔ�V'��n/�|�U�3��+���HyZ�� �	ޜm>���Rӥci����)��������JƋoA��Z6��M�A;�6G��0nq%� ��0���)f�VZr�H��9|+=�M'��+�^]��Msê�,��V��Ɏ���q���c�/K�i���-�g݈'�T�jI�ֿ���1���㾑��&$�=0���^^�L��;xЬ�W�>��q�����JsA����xUu)c�.6�<�QT��
�X��'�/^ '$Y�����K���]o��e_��}f��5c����z�����c��ֳ�A�p$o*�P&�2��qv�VB�	msLDQC���U�,�1J���B�M�!h��&c����3��''�	 ����>7'Rz�=�g!e5��xQ�C�/\��#P�O~s7�ل����K�`�#<G�X���i�4��&̡F���ʶ��|\k(�����Ub.L�e�K�@�I �lc��KK3�b*�-虳��O�J^w����x%�+�,	��D��[�Rdz�~g0�1�� �2�l�HF e�3��l�����O�����3������F���t�	��3*�7,e�NH`�����u��}�I������qS�7�=�J@��n;��u��@֙�TG�o�v��f���5��9���������5:�F�4;I=}Am�c��-ײ<�H�5�h{fK�4P�fç��E{|k����t9���;�4�Kw�㮐�L��fЙ.�9��6n�7���h����{���%h/
����z���Y`����$��N�9,��J}TB2��:���?�|h�Wj���*�tx�ďL���f�:���B�H����@��Q���F$�a���Bd��k�:�b��;@��D�F���R���,�� �> n�����k�{:SW
C0��DeN�V�B�����H8��6��DP�>�&`'�l��&Z�9�,�<%5�:��l8' �;�?�m!�N(bV��{��!��B��b�5�����j}���<9��\����|�u��kӛК�}�,�E�w�PZP}A�H� X���D����k�{�f�'s;!|I_/d����8Ǘ��VU��_�[�Z�bPRxZ�ˋF��"n�ܾ�y�h��CϏL.�D��`u[܏X{)9�z(n���IQ��ꈅ�"�#������8��'�%�E'>�-V\�4D�;`��V�B���NN���MR]
o#�C
�[�v�C��p�����2RT�my(a����C�����g�d�0�΋ ��a�T1��n�? Ʊ�v>Cؿ��bF�]F�"7>R�^��Õ��73��&�T+"H�V�(D�����]��Ǜ;Zt2P^c�$B�7��R������GP�L�|�v��ٺ�q�`�H�sO�K�i���;�����8�_eq1Z�E�e�vg�%�A��s�� �'q-��͝�x/g�� �܇��+�h��g����&�N���`/UI�*ǫ6�LТ���c�-5�:c���p�9~>�Қ���C8���?����[\�U��
�E�/J(P4t5۬�@�����}�w{��X����+��V��uc��k��f�&ʍ�"g����o�)�r_��Q�6{({LO1z�r�
���TX�YO}N�9$�V��O�d}\�8������]�������\NkIWrn���1ұY�tUb�03�vG��RCZ��"P�;C ������)#gc�VU3NqmWeON��_�Fظ:��9����hVzh��进�V�9�xd��;�ϋ��H:J$�d���J�+Ff�?>u���]5�E����h Ə�T�q��H��i���x}��ء�t*�ĳF٬IS<���?�N��TD�U�٧�Z�y��H"\[�����h6
��� LJ�!M`��<^:Q�TJ��%��䵣�t���3ε��W:Y�pCЫ�)v�"�vh�|p'5�@�-�3j���@�ܩ�D��%�/Z���[��n˺P=�9��s����u����ؽ�[ʅ��6�m����j�Р\Y~}��V��Ù�~O�G޲�J���t'�x`LO��22�C�Z�	HZ�$�����{l*�C!Ry1meJ���Í��űӆ�����BDnL����N�����=U/�̘���S�С���D|g�y�$�� gLi�ۘ9������Ô�Z�
�P�L�oc�inT�; �2�3щ,j�g=��(ǵ��ӹ���RB����n��K�����Y��N>��/�����:�w>]6��+� ��$�F�Zk���Y��{�^6���S�-E�0���zg)¢�SW#X�48�!l]8L��{�Ԍ�U��y�WsZ�d�uc���,��(�a�;�gH�XvQ*�Ü����4�}�,�|��:�fP�a�[�B#-�M�r
��]�e��E6(h�B�,;�E`�1��SM���,���q[CEvs�[�����g�RW
*��͜��-/����iX'-�s���-:�m�����J��EVj�.T
�2s�s��/%ѽzȏL(O����r(���0M"v�J���<=R=�X�2�h�����0�"������"]�^���fN.�q^�E�Jl5�-�c	��6�]Q���$��!;>�n�	,=`�*�6G��$�0q���*�eN\$�������mPc\�#��e�74T�jB�Of�@W�ţƀz�����.fj�
`�÷"��W�f�����i��;�����+f�ݫ�����x:~Nl�1@`��0��e԰������	L����0��8庋����%��!7w��uE��Z���r6�۱�c�ȾD>ڇ��}�Yڣ��?�,w0�D�\��t���A�=GJ���ܔ��Q�F�#��X�|�b"2W�1J2�8u��6��������~\����J���� <4�-C�*izh-���=L{��'���R������2���ޭ2@(����5�6\�h8�[�^��
dI�x���`��$'�J���E�{��ޘ�'mMW9ҨE%�e�攦$��C�, X��D��m��掟�����������"�	�����RQ��l��쎩�;HZ��#���Dk:b0��B�J�;U����/��^ 4)�irT�a��0�V�.�EZh�vG]��EV4�}�Ԧ�&-��"��7�Y`͂曩�|�M�~�qW����ΆXUH���%Au��/]�/\���̉�Z�U X�{~!;p5��E��>�x�����k�%���m�,����c&���p+v(�l���I�E;{�7�
�J[ݐ�$��ki���ֺ��X�Y�@��.�7�U�*��-����U9@G,�]����4�����c8���h_:�V&�3�}��S[�Bʹ��4К��5p���e?k늕��k�kCH�r̬�#4����
Zg�&�eh�b2�]�8&t�bc�:�Hd>�R!���0w����+�k�"��b�?[��y.�\�Z
��)�'��|��'bHǪ�6Eh5A{�k�Z�P�����JN�L
I���8��$ʦ����ǈ�!?g�{@�h�0z y��@����^c>p����v��̞o@�]�#��z�HJ���%x���:xs&���d�Ʈe���h�
���q��'�ɰ�sc������z����K��H�KE�{Y�O$~K�g�p�$t<.�s�c���s�]��mZH�D&�%�����K��&�SG�f��K��w{�#|�Q,�6�1�^��.�k�&Ț�T�!ׂ�����m��/Kk�H��EBo�:��f�	D0�'����3��jCl�^�q ���ۺ�gy>�c��c�1E*����S |����>gÐ$�4]@G�F�u��`h� �m�2�b��/�~�+�Vx�N�}!y��Ŭb�����ڏ��*�
dq	�C]��#�w�� �}����"Wlr������;źB��ф{z̷����jH%V�bB�M�%}X;��K!�x���:�IrV��-_o�ϒE����+!�,��A)�Ɂ�>�7���j,�m��2Vn8����l���ʑ�� CZٮ
�Z��G(�}��%7�	�M��&���"d�A��?�+1�K��#I9��(g���2�inc �ȥ�)Ï�=�����,|j;��A�������c�d�cr ��a�:������&�w�Vvg�unw�!�OuV�4�v%)3g�`��m����H����6`MML�Mq9��.ȒXmu������{93!�U�2J�����v�A��M�JT�;y�}�6�*�YK�{] ����,�Y�m��� Ip��X`�������gB���`9��G��"���W�����־�"���|�E�/�mK���lû��z�po��W�8��ד���0��5�>wɄ��X+�Cp������jwlT��S([�5���DB�$�S�e�7������·���	E�8h�)�a}���+pM09�	�+�������xł�2����Ȓ6p� ��M�ψ�+����� Sbp���ܸl�ޞ����"YY�c���Rf��4q©����Y�hʘ�B[w�����yY5�h`G��J.>���Yڂ ��{���%S3���K�ReQ:�-/�+x���-� c^ei�F
�u��|��������=1UՖ��쭟�u�Α�eE����͟��l'��k��N�,�F��]L
a��@�~\�Ck�����ۈ�L
3t��8�Tu0��J���^L~b�3�8�ϻ��+��������*��k;ص�@�Q�Y��8��a���%���dEE��4����>�oE��Iw]"�	HA\:�s#OD���[�,�	�>�9�݄P���Â;�T?�{/ٜ��P��1�	 恋�QX��f����Aŋ��D!������ӡ����T���ꪏ�p�Њ/3����A�l؄}�d\|&�)��4M�������M�� Z����y�
�Zî�:\ef$��ѡ�<�g��`�2дl	���q����j?Ņ��I�W"���/.&�ԸM<�������e�� n�)8���4��xm�UM��{y/bU
�&�X�⽏�	��J���2��|���,e��+2O �X<��^QI�6�+��"t��khJ��o����|�R��hf�F'� X��}T���������̨c�;�O�K�~�pA�����y������|�$��@��s,��H�GM9��3`)��K�чV`|��x&.�����Ж� �*�k�K���e�G0�r8E&?Oios�u�7�:�u$SM:*i��U��<1�6���d�q�"gG��m��L�2��h��&��1��JpTT��SċߋT���y���X���lpգ^�#���p�{�9��t�;~Hp8�	.d�Უ��}<9�B��]:eB�����'�HqC~�dJ�
���B8�.��;��쿾t�2�qMBBW@��EE��y���R$Y���"��wB/K�E�T�oSXa��]y�#u)��Sd(m�ϕ(�j�����q�7��:�E�L|h��A:4��s�u_�������^GI�>�4Sv��a�Yu���:1���j�';J�.�2����j��z��9������B,�~ڹq��N� �C�x!���i��\�\�l:!\�7MZBt�+?x)]o��%���o�(*���ȳl� �ۀ@�ca�45��$R�6��F$����x1pb�#�����;T�����:%fO��$�����,��*$�x�H��[<�8u��6��-��%��5���Ş	;!n�e�o]pO�T��fC���7��Ձ�1��n�iI��+DXY_�Glm���;NGT(/���9�[x+2������P��?���s]I����L���^~ͩ��#,R+�tD�Z����2#�+`����Cݜ�Y���E�w��_���{l7���Y|T#���'W��	;%�F˧ʓ^;#�E�����i*�ꔲ:d���O��l�m��2=U�U�\�K7��Zx�煃/@��g�0�a�]+)e$ ���1J8��IuǄZ��]Fg��{��^l��f��B!�_�3+��z��g�48�N�W����!I6ȉg�u.�3��bL�� O�-�
��	Lۍ�=�����߷��V����01����;]*|
')��X%��
YL�n6Z�W�
�HZ9�U8΋��kr�PM5ҙ-Vm��IDBX��.�=�/�0/�WE�N�K�|6�vS4�z�����@��?֭�	�E\� or`�����K�3���-���� �N�7WS\�N�;kn:A��$� |ך@��_�%׸ ���?7�Ĩ^�e�*`�=v|�S�'��ք�/��OS�^�sA��J�#΀�?�5+MsA��6�	�'�2�g�<h�g1sN�(�s(y%�ېhD�t�.�E��3Ϭy������^m�؁��q� e�n��S`�3�P�o�0p+�2]�%F����wM��;����5="�.��������S��W�]l�o�
�|^[�,9@~�9��ká>|g�vʘ��n�Q��j�u�Z��;qN�2��8?H�4�3�A�%�+��2���;����:"er�2��/�ƊMԢ���1�����I�_2ܟ��EP���� *uf��iǠN2���PR����m�YV3zl��ZY��GG��N�T��9`�3;��<<~-+�Ҷ�q^lH�kD-���M�'�u�2��x�ڻ�Q���~z��ho��M�h<�Eq�!��[�5*T�<��˽F���dǥ���N�������R
�ֱi Q��2;���=7vc7*��]��N���܁�2i��$[*5����aX�M�scP/6�K�����Rb���4�����r�j�sxuC^f�#�_G��M=�goW��R�)������<Q6�ծJ���ig!�*r7?;�Ǻ�KB�!�}��-�k�F%� �l{v����u,��������Ӄ��\�����������@H,�'5y{op�3�J-"����ψ�B�g���gOh<��b���9d_A���ޯ��fvn�x}N6�v�a�u��c/jN�G�M�v��9�i�+�����MD���SiU��5o��SA�pl|1�fƮY+�`;;��Q�l���]����ՉiH�]ðu�������_�Y�# )ƭ(V������*?���1����� Z�Q.���yw�P�<��C�/��GF�"�4}�.d�Q��r��p��*�3d�nˌ~�i/7�L��=q[���Є�\&۹����?��:�{[��$��T�)F
�u�����LYn�,�39@pޑ�!_@����ua��$,�71���!o���4��
��[J��B��}��&Q�0��}k��ؾ}�`L��y��$Q�~��P�湜�CC��W��8�/�_Z�+H,�%qǻ�)���-.n��û�e���7�_h9�x�0��XT;x��?K�\������G��`*I���`�I��<�����[��y�ئ�:��Q �
�@Z�'�J��}�4�^V�vΟ��� ��1󑌒��:IH�.�qB�����~��0�oY]P6���w�,{8��ɔn�\'%�)�I��ų,�RQ]��dZ�r��_����B=�ʘc|�?|�O��l'�(����p�u�����lh���]���0�M��z�I�^TW�U[C5�l���[,�n-q�H�W�=�<�!�tP�2m�k���\���sG���p��0��Rq�fk7\~ݓ�PW�B<a���R>��<�楀��f5�g�nbd �����)R�AL���f!0k�q�����L��F�I���N�8��wZ�e�p���+��Z��>��h첗=��!���N���-q���tξb`d�-�4�'>�W���(�mE)���h(z�yԋ�?0����>f�gO2~�b!�	6�.�|�ֽ����|�o{/Jʳ�9%�h�F�fG������]F��,��.�p�c>+6���<r�.��_��'���+��z�;G��  7�s�.o�P��������2%�����w*��� ���ߔ!��n� ��6�,n�����*㆚��+Q��.NL��U��p�_5���(n1� ΖͿ��$���\�����O��KPN��)ݏ�5ŰҬ&�*ve���7e#�`���t�ڪ�g�M����{��ʺ�F�6	_p�be]�XO����!��80 D>2�n;Yd����>?�^|!�j	`rZZYO{	+�Fj1k:6G��wJF�-k6�1%����e�t�Be����@F֮Ym�3\��"���Nˁ�rԛ��������V�U�9�ݤ�D7��"'QGKxi[n�mɑ6�ɉ�99j��;���x|�FA`G��o]f�dǐ���x*F�{�޾L�o���#ǿ�}��Bhoߣ�kE����e���,XV�>�<��dIu�b�ƞ�3،
~��I�)��h��7_d��W_h����Ȇ]�ǳ�ӆ�/�o51꾻�_	f<?�����PI�n��)��J��7Kup�ao)�F����#"�
X��1r>�˙�>n/���c�'��mxά�!�hz��M�3�3n�Z�� ɏ��f���ߣ�G~D�;�?$��}�� �����ճ�V�u�z���.\*祯��� r�ޡ��K���]B�o< U�mXh���.��g�x��ߓ��,�r0pQ^VI�1�	��2|/�0��^��?�տ]8�?<e�O��j׉O����<��dm�^��O4�n��*�ט��6t:��� P4��89(�`����r�eHh*Dҟ�J��p�ɗrE�_0ъɛ��o8ms%�D�0t���k��p�?6[���ď�{���|&��A����/��o�����l���T>NΤ@5�)4f�&�n�}�ǁ&`�|4KQ)>l+X�ڡ_���ج�O�jX�[���VX�sY����8���5q�^>��#�����;��5�&X�6�������!/"���+��J=|[�E\ �ي� �ob2�վ+8�m���\|�z��	WB�*o�8��ʁ8�uV"�+=�T����h&�j�^xU���*�C~����?J�"���$�'�ֳ�-����--�R&���?��kc!�(��a�87P��Y�ObA�r�a5���!�L܋7� �TAMmK�Be �/WGP�:X�tp��8��
K�`D�y �{����gA�����s�������s��)�*=mY���p�ȼ�0|C��b�`Pǘ�s]l�F��ߨ�6g�_���v�ƶ*A��f@�6���3�J��p<�X��~Q/X��U~�9?ѳ�fſ�=�Ϩ�߲����ܴ������ܓy����0圛�S�>]�E�t�]���^X�[��9�m��H��Y�f�����V"�>�*�V��x��9�CV��]��`��$�OY9Z�oC�>�u�l��u���W�/!�N�/ӳ�?f>�eO�1c��lh�h�Pz���ˈ��B�Ȓ2��&=op����=������H�I��3�{���=Q���m��t��Ϳ���
����IPsru�G�����~]~��x��`�Aa�C��ދ��玓�
�rz��)?��H�}��|\U1s��b�_2j��a�tS!��nK���������Sg`�լ��i��%����� v�kOO��{3� �h�F��D�e�Q�?D�r�X�sv�n����dG0�YN�/��Wl=�wEz�R��U�����[�I!_�r�{�����^�@�?�5vA�c&�r���8��'"u�o-^�f���D�D�t����+nHL����,�&a;���i����.��Mh�)�#z/�J��s�;�Կ�Ќ�����ĭ|�:�Y�N���-r�_s.О�I,�C�,n;~ECy[-&^Ӿ F*>ⳓS��(I26��d%$m�\��b�)�H�bΜ��,~ͻՁ!����o���$�ac)!5scb2�|=��z Vc�9䐏|�2����=GA�6N^���t2�zh��2������݆�����}�\���(׶��;�8�+:�"����X�u���Z3x��`cu#�j8��O��]:��%��5mJv3�:�������u�Rj��
g��j�^ �����N@��u9�*�q�NT�O4�C2c7���3:B�Ǒ;�1p���0��.��8q0Rٝ��uq��b�2���G��M�_/<�b��[���~!��E�ģ��IM����4���,�(��!�^'
?�H�Qm+4�>���]�g�L�>T@�eY0�}��m�	yD�Wd�K9��iP�Ý���q܍����V�P��
�u����)P|���z��`��{�G	dۄ���j��|a@Q�GsZӠ�A0��5�&*����N�t�x������ء3m�o��E'{��X�����oYÐb����.���Zͦ�\)=�T,�H@n��[������Q��d�J���I�u�|��H�*���� A�9h>	��ƍV�i�sD��7��������I�:l��]�2�P���[|��u��z�%��<� ����#����ҖP�e�׽i
�㘖'��C�1\X�)��E�!N���.�b���-��o��O:��tW C5�X6�/��b�B�G�[6n%F^�#��G#��"�k�U�����Y�����f�79g妨&��OK����A��yw6¸[	���@"P�m��vR���b��=�L�C��RN������C9F7d�H{L��S��H��+Z�R+`0�8���Z�۶Ǡ�Ndv��LvX<ͷ�K�K��k���m�̆��!�Sz� �p~�0)�5%~�8A�t����ܧ�L-B������Qd8Ҫo�����.ط�K����{^k�hSM�ƫ�1\��p�&��*X
p��aRk�(�I�kZ2�4��_p�{�e��~H"|~;�)1uX�Vf��0uy�|��@t����Z?Aw�Ar24Ybx�ۿ��4N��Џ����Ü`�����6S��b�Im6[��;���!"l˝C�U���\Å����j�dN��@ �ދ`��G�����r������ҡi֒	��j۟�]hq�x���3�I>#2#Db�V�G�<P�6�
�بʰ�h��E	�[�L��5�d�\��~�1���uO:蟨�z<0�k|��#HP!���Y�,|��eFH���C $�%���t��0���~$�hڔ<%��$�e�ޔh����(�r`��y�=P_�A&���­��,��?�P��^H��R[�rI0v�����y+������X��(,.Z>p��:
PCf�I��H|������e[�ڭV�Ϳ������,�Cx
!3��yH�*�x���'<�������81���n�af� wt�@ej�Z0��[*l�u�=ߎy��h9N�'�2�j
r�gv��)�(�<�K[���I�
�4�	�e�D>V|��L|�o�\7�E�SV�U�4Q�E7��%�:0@�*J���Gb;����P�f@��I�$�Ǚ���k2��k��[�|k^];���9U���r��>�A���������J�=��P�m� �[�Fj�r�����(��pqdFݐN�{�Q~%9�"n�*kbG��ܺ�ιt��ŕ+Gr�����)���$A�a�S�Vý�bPNǈ�N�	x��B �2��~� �����=�'Q��g	��$#qOH����W�8hVRH?nպ�� �*gX{t��a�c�8,f)�����<nZ�<�r]���7��,�@��Ԛݪ*�5�-vP�������I��mt(����Z���J�|w����}� �i�ތ������N��9=]i,�L�J���?y�s��0���֟�"�X��}�h9�=�/���1N��Û��xb^��E[D*+�Dy���Պ���u6��6B�rU�E/w�~�b)�W�d�KH��r����B��Z����9}�o�u!;�op���DP�	s�G'..h_���"�		�M!���X��|L)��fT��W���O�6aE���:7^�7��b��K=��A'����]��w�R�~N��\ӎA���ic�VF�jȽ�U����9N�I���������qw�i[�x�W���Z�;���V	ʺ�����YY��m�W:~��$�W��U�)U(-���ժr�k����I�#�I'gq��|�]*K��T�^��1p��BP�l�9��;7
r8�B ����������u9K�Oֈd�q��{��y���g)�&�㍠'q�1��q�+�[���x��M��Ͳ�8Th>E'��*0��T���U�u�Ķ�>/1��)6w*�ە����jZ�^�?ODz�R�B�!�~uG\��y� ��_DZ��!�k��c��8��(VM|@u&n���ŕ!�1:<� 8�;�7�.켦l�1+��y�(�r8T?�q�p��8����|��jH}u��{��+�@��- ��߿h�ֱ�-Ѓ���&v+9���~r䄽�Vz�&]���ۖ� B�=�p�������]�C��
�qwlɡ��"�b6r�6�FO}ߩ���z�BB+�0G�,��`�Dr˭\>F�͈�:�+Y���#Vf�}+��,�؄�����w�k�S���>�G�b0Y�H�@b��AA��f~� W�񨴺�7uN�T^�β��h���SR�j���>Z0���y�I�4�-߯ɀTI�4 %�~&�VZ��k��w�.{N��'2׷��ֈ5 3�O��DI��X���/Ku.'�F��7%,��ݮ��N/�����[�&=�y23�<#�U�,���:��5Ư�4��G����/{��,1<rf��W&k$&�F�;���Lb�����H�D�ROx����~��F�Df���=O�u��on��t��y�'�&r=�
��g�m�&r�s|Ԝl�_�⼾".&ǘ3Erw�y���|7�s�`X�����t|���Φ���
z7ε�\��q�/�O��2$v�&ab�O���7O)t�++��������[6xJ�;"n'�b�y@T�qf�;�	�*_�u����?��z~��������q�τ00u��$�~?e\��i�Qe�����y����	B�S�\�{2����F� U�qB��V)���[��[� 1>��3���NƮ�R�fo!��/wG�_"<l-CBwQG��"c<*{�9��γ���'�!�sYd˶ij�K�:�(i��oQ�Uj8
ș�8޴q��Ƣc�	�7�U�NI��9�w+Y�M�QF��ԁ=V���?ʑԅ�`ڝc�GT��wTK��,QHը���9�-��ù3�����fH�9�ykB��� 1�ƫ�7�@�#�4��o4Ty�ٽΞ>�MyM3ݷ�g��gj/Rg��d=��+�[���3��E�)އ���6E'��85&���[*y�H���o��;�w��% e�Ǥ�����g�j��X���7���)/2M!;+FC	�X
�Ѱ��9��G��!�4O3V�B~iX_���<ͰV�y=��$3�?�����\�P�Ţ,ĲFlLj��M��~S�w
�3����K�I���X�vg�mD�P�uݨr��oI(��|*�)%oKOO�_�����)�*���4�{.}pw�Z \2��p�K:hG��Fwd`2����7��YR����~c��C�$�!��a>Kgz���)�.q�O�s�B�J;s��*W�Q�� ��Gώ�|,��5\�~����Y;a,���_e6��nF���2A���_�l��g��.h5�S���R�Κ@�C��+�<�F;*��<$)���~��H�_ۍ'�W	a�%K�y�	+�
:(������ؠzM���� �ި�۾V0�o���yb��E{R#��Nڦʟ�v�JM�����cs��D��p��n�����A�Ձ�Y5uh˅�g�t_iA%S�c��[�XPs�
�@BH�$VFi�$�O�e/�H���K�"�AVU������y���ʄ�6�D��^���'��c]\�nÔڣ7l4IX����2��c��e��X�YK�S[
�{؜Ǳ�j�̺��X�bI>��85�FH��T�e�:��՛Tw���6�|9�/��4�������D�Vd!���bqW����W۱�P"$I{rL���A7qudGrb��Z`f,����I���P|���"��|~RG��A���md��O�@*�2�^F��.c���#8�f���`�C$'IJ����c6��;��Jv���q�� ������R��2��`�m��.��^{��Q� �lU\��

�rj1�X��Y��Rt����qU1��<�CR۵;�c�e:&ʁB& f�6��s�3J��YՆC��ch�`���C�	��y��Vh��mKj:�zh�TT�����K>��X�ZD+�^�%�Z�eo�z�c���}ѳŬ���b���Բ�|�͈/�����B����}�>�Rp[L"�����9����O��CoRN6�!n�b�4����E	�������ڒF�*��oX~�*%��,���:_�}��>G���r� �S�_˂ۿ��m�����9yT�^s��/��F\페ݝ1�F$W5���'�Y�w5�(�O�d�x{Ƃ��·�����%Q���ҋ�z�4����m��"�H5�6�\U8�k��AV/
��ޑޡ~roj9K��]���/C�^6���#��g|���zl��ۑ�W�6�b���f�mb6�\}]o
���(��v%���jph�
���;��F�
rZ9@`������'�#�W�5{�!��e0��*	V�.�4��:+��Ws�~H=�}e���t �j�+'����Aą�+F��\����7�N���Aς����Ϗ�T����4�KF���0��������m��܎z��In=��Gk�+Ss�X�����qA]"��$]S�Z*���7X��+�t�{�-~?`��7�v���1]y���Cϣ�6�����M�Ќf@�������S5�@[���O�G�^�ͬb�k�%�F��#YfM}�(L8��h(E�	Smݧ�xT�k��2]�K�17+��ы���'��+u���Й�I��2\��ۀT��B`�ͮ�%�G��s:"ǀ�����yk�L�<��ٹ��8�G3�c���!�C�J�:�X��˞���ŀ��Pv����V/1�-���ڏW�ū�P�m����Λ.H �>�V
�X�ݡɜ�P��E%�)����rc�4,n=Jhwv+ܬ3; �mc`����Y=�dd�\����������<���WNt��t�-�1W�����ɐ�Q^�/"�Wx5���a������|�c���x� 9Z�yx`b$a(�X.PA�y�����iù����A�Ny!O��a�Vc7Y�jg�x������;O�C��fA�&L���TY��g/����3QIl4�Q^�I���U�ƌ����Ӭ�;�@�#��r��t���+3�v��Df�q\}�;�v��t���>o+B.l��fD�X�`J5�S8ۂQ͟یy%!�t��J�H"o˴�I�˾�D~�
r�b��a��G��B�i����I��4v��Ϋ�Ɔ��/F���@����	�ց`��g8F����6���@������Kw���QE�ъ�b�Վy��x7h�i��!��qJqB!l��X���	�	;�Nu�7�G	��#n������0f^P����T��x��R���D
��4R��\I��(�2b+�7���
2ek��rHd ��^���o�A��$<����>�( �iL��㲊E���G��FL`���i�
��,�)14<�e��4��3�� � �f���4d�5�N����OCb�8���!b��X���ƥP��%�sj����m�e$�:O�Q��LCo�=�!17:iBH?�v��}]L>�#M�X�pƅ9V���Z���#��U��)D��8�%�3�'�5�؛̄� ]�Tw�O��E�*Jx�x�ކ� 8�|$NDr06�iN�[�� q[M��-�w�L�R�(�5�b�E}�ء���wx`��s����_�9b�K�Y��_�@L`Ip�_��j�P��},�O/��� <mzt'�bp���W���t�A#����Ǡ�'�LY����U�h k�qpWb9e0��o_�\�#*���&��@(��/��(RU�y�N�����:���qao+^
���h*R�+�|mu��L�}���%�W���P첯�1!vp��٤iN�'�9�q��s��t��$�K:��?�7�V��Ht�]��a3$|�taѼ��t��/'`�j����N}���Ǡue{�Z,&_�6m�C�r�E<9�ڢ������O$8"k��b4U	��0�ozNv�����ӌ,y����E��KV���̯,��#<$���_Iv�7M
���^��Y%4Z�F�H�WN:��;�"LRurۘ*�������*E��/-��@x��2O�	�����<u	��ț�M�&X��������O�94��<jo�����R�*!�<�s�"%��o�4�(Y�ӫ���@�y��B�2�t)�u��P�y}a��(EC�x�<Q͆X����K��3 ��5��4�ϭ��o�\�-���5�A�n��Fɀ�'0 8�eT���]q;�!˞f��5�!](�z�����4:R�� ���1I�6Ўj���B�2�&{U������;�C��ݷd�V�*�X��4/z�!ㆴ�N�ԝ��Y�}^��Շݞݦ��s�3�����c=�f(e7�;���:Wa�툓�*�dSD�̎y�?mq�����CH+nD�q-q@�^��|[��������*g*P����G��L	��əD��}��Ց��tY��>+O�ݔ���:��d'������ѐK�����ʥ.��l�,�a*��q�V&�t���[��$:�CpO��=x��֪w��`ߦ+݂�g�'�!ꬋ��PR���*�r!9+^Э��Ҧ���$bz=��P�QY����y��+1<�熉�lҚf��*jb�ڼ�r�X<s�p��F��*0�m�i���kzR	�M�'���!y�t��T �`Q?ε,��s�k!�JZm7�y���LI��A����������|Z�8m(f�ӕC{�p�}ԙA c�	�H�pN9���!PF�Ce����M����	ԧ]�R�0T�(^'�1��ܵ�awD`Q��x9m�E��A_��4�b�u\X������/������p.���g�
��))�5P9Ċ�L��,���{l��aK�Ir�����[ �)����Mq�x���H�O!�ȟ�&E˩���\a�6�`Ħb��HX��Lf��+�ʃ,�C�U��ۚi�?U��-���K��y:�sgK���:ۊ!�٩a5b���a(�J6B�#q���4k�X��&To�j]zj�W�zb5�~q�?����r>%F�t	2���7$���+Ɠ]*�w!�p���:}l~uخqm��/.�c��؄Xՠ�j��Ř���� 엵���X��M}�v���jD8�(+U|>a/����uM���b��� �G�-��>]sU��>ܛ�:���I�4)��w��к��^T��`��¤X3d�L�b-Y��2u��u�qk'=�8�坄��J<�M�c��5��q���Z�4 %9_�C���A���\�0@&(=����Ʒ��¹I�9Ǩ	
�\>e<b�����u�۔����owsb(]i&�����c��E�k��TNR��Jx�~�#&`r�f�4S�L_�ql��;1�qۦ8��"x&[
9�`ٳ�+�z����c`X��q��,z��N~c����mR"EYͩ�*���^� ���~9\� �G2!O��N:�lh~=PlE<Ս���a�޴��E�������"j���<ŮP���B�/]�ADL�^���lw��H�N��&�E":��(hS�)�n��� E'1ÿ��p�"���*���5A_Q,��{��/�Hz� �֥;�u�T���}�� Im"�]�<mE����ߘ�;��|^\��oaC����WSnS�S��!*���r��i�Gz�Z|Px�.׍Z4i$U�ۦ8��2���h̕V�X[�c�E��͉:��ΜS������q���I'n��T�� ��(`[e޺(�ޝ�+�0k��⼝l�T"K�d��e�(��w��E�����8i��Ő|*2�H�(]�0�huH؟�ޭ5�ma����[�_'�����L���~�@uW�}\�S�G����/�K�s�}טud�4����&l���kXŜ��f��ÁT�6G-zh$���*:�d����:�5�N��f�F��2vulY�6�$��#EY�ᲂ�ʙڑ��6�JiG/�(漲m3��%$ƙ����w�˲���Ap'�'�U���-<`s?�	�ƨ�9n�T$ϟ2Y�c��8�՛�m���}=Џ�P>5:�p��#�L���9ʬ���;��@]�� oe�>�(|op&��I��.��u�8
��E��vb���J;5a7�8�o���~^[Ƃ�$2�f�J��f�(�j�R����;q/j������yA�o��2{P)��:�R.-d ޫ&���&�,�%��O��p���<��w��XC-^�\_[����݉wi�4h.F
H�٥	+Ą�\��g+�5����W���H/,��b���
�c\;�i�{�dHL�ZŸ�B���?�{�m����78ҩ�b=~��&d���t�~�����^$ ��\)y$�ʩ��MYL٦*��K����������_.Нx��y����w`�X��ۓP��o��q5A]S�:<�S�moڸhD�k��&1�y��8��3��������ި�J1\��]�V����v}p
��ač����v8I�% �ۗ��:�C�?��1�Rou�eQ�i�~V��S�X(�|�s�x��@	DcM��,|��7&���p�k\t��o<'Xt��"n����N]j\�c+�,���#G]��0�_���ܻX��`��2��4;sI���tD�L�H	L" pB��"�q�t�޾8��
����5(_D�`A�!��H���'�k$xl���]����>�)��85���f��?���ݛU�,bO)?I������R��R�YΛv��"������g��GxA#�M���6�X�uw�e�1�g@	�)2I�LF��,��ن3Q3n�D@�<6����\�wfPKK���>���Mn��C'�mη�)��[F˅U&D���|)09d�l���1q��~��$_��B���ݸE�|c��:OÊ�7�g�BW���c,��	�����Mc,N$�~�$��eF�O!Y%:���]؇v� ORUi��.�xs��y�~�uNLMD���^�2u��ɂڛ�#N�\�@)�7t�%���/H��XU��GKe}��V���$�}�}�����(Hݤ��β ��|������d��U&G�AN_iM�SPn���&�6r�e^���}�nf�׋З6Dۤ�~.��u����Z8�{[,1zy_��&]���2�uylVz���A])�ۉb��h��U�������n���(�v{���o��X�J�c�#<5|�Ű.������J��t��_�s,�%�6���L;OO%q��㻓�r_�rG�&�&�u�6�ɽ����w:��J��:�j�Z �/W�fc����'��k_O8��2*w���p;Y%^(��@� 6��8+�)�冣��J|�(*�jT{�,S�dHm��yyI�Ar�F������/�ի>��TD�:��;��F�V%��m'��{zq�98zU�򧐢�W��,,9SJ��Ek 1/�
&�\�}S�-L��Wc��6���|1�j��p��ȑKImW��.	gt7�)2�Vۆ4� ���4��� Qe=��覭!*��j���}xC[>A|q���P^�}�����U7A;��l���o���Q\��awC"���6��@c�]���,s��S��HM�Z�Nj���p�C�#�B��`��xlp�M>�<@./��9���sm*�óJ��e������n�?.���T��'%�
\p �h�ާ�t1��� [�pyZg`�ɦNb��WF�n���	�Y<��"G��}��?�Oj������|Lu�j'��I�<�}���Q����_�$1Yiljj��р�� >���HW��i�$dǬ��U��J�~�{�	1���Ŗ���0V�m�+�ܺb�Χ�4&��h�e����+��n��5O��N�s;=��0�r>�F¾�ݒ�'��t�n�+h�6Z|��;H8d�h�|ƌ�Z�R���#'VZ�ʏ&&J�EH!�QF��n{.��S��dN�X8�:K�gzBc,�fb۸��������հ��.u�H:�SN6#��|�[Q�
G�#���|����	
�'���� Lt�o�M"��P��NK�#����w��h��q�_;7F`1]l�5�`�V���Kљr��q%kE%A���i��2�F�����#ɂŚ�K����'������H1|���"0�_!��r�ڲ��Y�K�zV|�2f��F-�'�J�C�5�cK�+8�m"	��B�'��O���<���<�E��#�fN/��!-Gƶ�.R��!�"ZFΫ��l9�HK��ɭ���M��2�b��rЀ'��}܆�v{���5~�]�Vo�Fݥp�-��S����N�2�;z
/�x����!�bس�צu���_��e��*M��4�(ŝ��%9��'��O���=��p���4N�\��[�����	I���C�+��LL�*���H�{\pW�k$~�O㲥L|�b���<���3^Z�k�5����,���]�|��&�C�cR��D�"c�+8�a���50�
ig��(�%�VU]�lM>��g`�GU�s���K��1[b�h�TZP(]���6M@W��)�U���'�������W{u������9U:@��mz�B�+�t��$��ۊK�������sV�PƲ�}���e��$�^f��B(���m��e��}��a���Z�QZ��~%��HFA�Ǖ�R�h9PY�"H/���W�b~�Gx���q���	FD)n� ��P�ȹ�H����`rӕ�P��o�����RWO��Zcf?@��"�UaJt���O�$�LH&��Sʺf�]�+�>:s&d�Zػ�`�t<�i;=b��l�m����m~����^�@O���1��L"D�+�uNVedV ��/O	UQ#=�����<C�r�|���Q�D�}�p_��zq���"ߚ���2��F���`iN�֨s��I����:m����u}��,�4���L��l|@q�a-GH�s�{mW�}Z�h[�r��o���ļ#�/%���Zh����g�t�BRFϏ|�D�6�P�l���+��CL�9��<���� �?ﴹ$��tiN��I�7"T�są�y8�E��?薋G�9�ݡ���	�K�Q}m
}���"����)UJ���^�5(����X��a�g	B���r�{2��ָh�c�>*6��FbihB��)� �f|M��2���!*�Q����<[k����-Vހm�6�9|)�i����J������G��˥M��L���r��jw����b	]1i��5�7��`�f4��r�g��>�䉫��,�MLsE�ixxlVx,�D�-����х2��#^����;�9�Vz��"O�:��h�;23u��N���a�}�HǥPb$�?�өZG��1z�:̧���K���}�9OZXƔ��f�����ڑ+G�[��D[t�� o��68gm̟��+��HH'�-%�T�#-���*�j&�������pe����p��,Wm�@|�g�P�O|?H+ٍ��à9�<Ш�UĤú�.�P(�M�m����S��d[rMs�0�����y���n)�ꖋִ0v�Ú/dI�d�^?����"�r*������D�;�޴#R��Q��:{3B�D�d����3�T���^B�`�h��rCb@1�<�5���;���䖾뤷������=�_?K@�_�x�����0�����Ľ`d�Oy�'��K�(��I����ª� ��x�cAN��z�hW�aK)����*G���B�߽��-�����=&��R9H�M�Zq��:P�K����!�Τ�cz�>`U&���=�y<�oP�8�B�Wj,�Wz6s=�)qb�Ps_����թ�L��0��}�!� ��^7����o�Q�����T��gY�Γ/���Ѐ�e��(����������ϫ�/enh=Fw����@�0���� �����>j���w����=�o	��5�Sl��Ÿ] '=��@�!p��|���sf�1ZT�'��n���x�ȓ[(�6X�7L	�yN�TV"wRJ�Ш�[s9�5�ۨ��Kl��եjJ����[S��X�܇Sp�?��t����rӷf������m�a��@��A��n��<��)H������J���ȓi�P����"v�J��A+��0�#46g����v8: ��`�&s�#����P&RI��B�oJ 0��С@H���BG.��H䔷iUĥ��{;-fKV��NS|}f��0,k��^�o6��b�/
�!�O�@���/�g�d�`���e��I��-)��S������$i�V���Z�z!Q� ��6T%c-��n�R�}�ҵ��e�ެ���b{��%������LV�}F1r��W�4����'��]Yr0��{���M�W�q$sr��$��~�5dI��]���vv�C��C���R��θ�,`
���!�PP�E}9c��5�i�w͡Xw �o1���|�jj���8/���L�M��%zK{�Bx'�Wvl�w]�.�2��a:�F'�l�/��!�x6�zZ~D}ݫU#�I�T�]n�\`	��Ǽ�Jc=�N��)�G�� ���^h)��c?{X��t�6]b�獽�US��y~�B��rc�/�>��^���B����)}�6$���~	f�>�rcɎ��W>����(��)vFݥ�BH�U�T�7����}�X��j(C��2���y���,)��#K%��FYӄ����.
����U����)R����*&��eh�ٙ���6D���S����Fx��2� �\,@c0ن
� �yJN@^i�c���J��9�J�Y��iY#ib*���ζ�}�����~��q��AjDUX����Cn��9�F���2�/�e�:��H���*c0MapgсF��\d�kq�X��Ys9�I���]�����_/f �Jr�=����0��@�H��KJ��:	\����H!�W����v2�x�x�i�;���#3*#�F��/� �ҋd��%�f��,��Q��Y�T���	�4[�@��%~w���g�~E������0�yM�.(cn#��n�Rv��Rl�YE�%��/�r�V��,>���b
7N�66�"��)�<YN�m	Cmt�� j��\�ɓ�vXQ��&+���:Qx�r0E�Y� ��G7�����ُ���(�X"3�$�0l��Hyj�_�����]c"����m1�[��TAn�j�&��wFw����ʒ�W%���Mᱬ�V_�e}�o���=�X|6b̄�6chR!��@ �+����t�l/�!�cgPVd��p$��1<9M��Q EK�Y#���d���Z��/�3��pZª�z~g�,�T��S��_�M��΢��cx��E��m���c@S~sJK?��_W�>[�U-�ngށ�Lڒئ�p�EE���A��Ѵ��ͪ�hD )�3�9J+Ӑ�kC��֎2j�!p�?/��WţA��>}}e7�������Z�����o�0Z�f���hMmK������W� 2����\i4�y���v��@Mp	G]����v���|^k`^��)ת� H|�I
$_&{�W'O��u�?�w΋\���$g)騙�vJ�w_��M�W���.�M��=�c` ŉ)	����<)n��J��x ~��T=����0��Q���1d#�gL��Tݘ�6࿴vm��@�*�('7���b!-��.�a�R�}ອB��76���篧�a8��lr��w���v���
׌v�3B<�.V�����8�g&�����]KWn�,	��dX�1܉+��`�Q}��[�*����,�i�K֓��B�8J*����Wy��ą���a{�DaDߘ������.��p�䭦��WA��՗i�T'����!02�d�w��[� �	��t}YJl�������[�B���S�^.	;D�ƫ���ko���E����pc�ǀ��M����<qL��a�I�6my�.���5
�bI5<���J��Q�0�~5�ivr��}��,��)�*w���jx�Q�M�[��
G�k��-���~rB���܁a���:��u��D�5w)�[@��N?��ο�HdZ� ��zҳ �f�"z�m=a�}���q�(�c�thV���&��&(H���wt�5��-Aq��yG�����W�#P��"���[��Q�7�b򓿮[7捨��X�
ʼc��~~y�9�hy��^U�S��5�\KP��`<"L�K�SzF�"G׷�?���<Cͻ��+!�`��6��ڞ���@�m��b.:V��զ`������מ����|�+5����_��	���NG�b�Qzh��l<g@��W.�q���:+��3j���Q�2�����^��+���	R:H1e�A���t�`�y`�H%D��6hǄ��)wG����{A�Yy�`O��/��%�5:�|[0Y��������<��y?q,]��m-DۃF�����G/	��64��gh�[]����c��ەaL�:v�L(��)�������0V�f�H�:Z�FH��G��!R�Tf�LC4eQCr�xh[�@q�婑����8�������s�k
���KdO/��q���*.T>	w^G���+�0M�����V�1�5��Q\S����{���m+�R�����]eL�_a*&�-CD�G�f�!�*�3��a�g���#�cX�2�? _-�B��;���S�;)fƒ[Hj��O|���u�u��{����2c��%��W�7t�ϔ1�p@#�����k"++F�_�Q��ma�ޓ������nK*�DoK57�+OF�� �a(9��dW4��@�5,�+�x��J�v!u�$���1x�JH��7s�J[;7��!*NV·��H(d�"�5z{coi��4Sj8�u�'V���u_���un�u3{!9���I$n�OZ���d?U�.�A��ψ��]Zw�z���땇�C>�u-�I*�)�N!%�m�Q���֏�{�I�	�E�~��_+�nr�E~�r����HRCbX�/gK�'ֆ�?�E���kuS��aܶ��\��beU,�3QD��r�8SJj�}�Jٍ$�O�ZV�H�L/./���qc%�F���Y��q���@�;ᄋ��w���|�")b���i�ߒQ��,Ld�k��_�Xb?��M��X�,�+7���';L�iN�eCl�L�Ry{�q]���[�?�=eMT)������¤^���Q\¹�ً�~����g�\d�~0������X�NH�R�n��v���t8��zh$X���=�o�&r�������>���ּ*�^���%��"�Ӯ�{�f6��Q�V�YM���
+ˈ�k\��I�s�J�x�Q��0�]�$G;,�%[<�'�Q��mc�y���gR/�E3����)b�&���p�F�
�p��U�yF6lo�ϩec�	����3,�[��i���(�}N�ij@%:�1�)�.^��)է��E��ΪI�(�a45Xly19���K����f.!ų�T<�!�W��2�P���ab8�-������MJ(8�;Ο��w�$Fɲpxx���Eh�����IR�2�������"`���l�j�N��Qp��5�Pj::��J��\u V�,�'�x��7@**%hT�
�|����L��R4�s�#���a]�3�_q'�0ck���}ub�1�L &�V�(6O3H�:L��&�>Ŕ��P8����9:��9UB���l�T����FK-Lx$6<4m��ٷ���--��<	ZWv �, h�в;�0+����]���O�n!��IH����	���e��%^�+o·�kH
��
59o,��Qrv����hW�ߦ�u����N�b���6�Y�DT�mqx�ᘄi	���-��^b"pr3�#�>�tnG�̵'�r�	(Jm�Q�;�{U��^�5M"	wl�7b��vm�a�S��Y��υ笁}%\��饾�v*k���.��@EP�ĩ�ڻd7P��q~�KCPg���Ĳ$���7j�,��=i[�|���=9G�@ʚ�6�y���ٰE��U�ٮ�c�	�*�I��>}6KWM�#��:���^�{���p�G����x�%0��CC&�iZ|���$t�-e D�b��X�yѳT���|v��W0;�{�W��܄�*s�M �:��UzA��߼��WIv,���#��"ڄl�e


b��1�_+��W$yc���äY���y[/��)Ds?Y!q�v�h���$��K��y]:9�' �U��rFh��ZO�����5y�8Ζ�oMoW�nf��￦���nօ�����lz�^f��1ð�Q��<R�"U���î��&��z�����NC�A�!��|���A���L� ���E�!:@��d	Q�kWs_g�/�X�E�ZH|��Wzoܰ��J����Wɞ~����U���>�K��yN�E��c��*��h�b���[M7p�T�MW	I��B�y�Q�
�����#4�L��<�L-�9�A�`n�]�3r��T�(�gmb �9�k��{�Et�D���l׌�ˡ���%�|t}��$QQ�xAGo>-��eߘ#no�b����-��o��q�XQ��t�5uC~��৤?3��%L�Ȯɾ�E�ErD�T������V�~>��'9�$�L=F�	RB�6�N���&4�� x BI8�y/��*�o��^�$����?��
 b���P�{�'��:O�#�6p��.��Z�dwv�G���ޅc ����ԓPy�N=����Q��q'W�*R<1��@L�^�
�}F{gy�Ö�D��f�������V�pq]/��VKZ\#������e�K�y��h��	3!P���m���\�21SL�8�׋�y�����րdޒ4��k��[���Om�-?�e�C����#�"��I�������Q#�@���'TU��6��v��֗5q��������+CC�PK7�o3O�����t2�pț�vjp���=���/(ӻ�����g�U,���Vc�G*�����v�Yt�H� eyZ�2m��.�Q�E�E��r�6ě�wI��ϴc��A�|+��P�8���>׳B�w�	zz�s��eq��5p�,�u���c��jfQ"^*����c�y��ĵ��K��쑲dp���eɧ�� � ^;�v}��mϙ���dG�|����O.kmsMI_��@���Ҥu{3#�/�`F��j��Mh�����E�6�~�,����L�]��a=Jw +@��_LS�D��±n^;z4�m��C�5��ۆ+�^
n��e@s���E::'��	�7�>o�b1��������W;����ڒ���h��H ���X7/���R�"}�r&�m�@��*�q���sZ�����~u^]��&��D?�+����ȼf��Ø��I[w�N�"Q��$y��*k>X歖��/A&���N>�	�IU	��x�Vw�j��e^�t8*�H&�- $r�<r(w��ڶ~��c����mRφ����(����o�E���x�`�n@�ɉ:�3ȹs;� ��IyN�/����z�[�50�_=X�fA/���U���a�9,W���pٗ��Q��.�%Ub���K� ���ϧ�U+�l9n��"��e����v�X�1.q��;�>h�A�"U3Q�[�JFƿ��^:W�� wI`�����/�`��Dhp,8�	眬�A�95ʯ��q5=����Ѷ}2X%�W^ì�����ʄGo7������OQ�yZ��u�y���A��R��]Q>R_����#�����8���
A�q�"'no�"��U�9Wĉ�!�M����g���DY�r��W���X��H���iC	w�ӡ�W�d����n)5ifN_R7S��B���0ͽ�� &��}Pٿt�cƀ�q,]>�:������*鍩���q�(MΥ3�#�_��Ϣ#�%�?5@��+],7�x�BR���h�ǻ��i����
���N��-��X�A'�HƸ�ۖ`����ڄ]��4Q��j]7V����e4��H�Л6v\ڪ}�G�`�0�v�4�5�y�f���5ݚ:��;|7�m]���;��9<I0�BA�Xs[?��=�h�V"w�΁�#ڥƂ�0M������P�lVX
h=���-������7��a��є�?��L�I��&��r���_�pu�R��lKum����Y��o�Ա 4���]������T�#��nM$��~���U��Hڏ��D���h75~^�L�%N�csa�!���C>�uK8�e��^�Bɢ8%k>��_���U�@�,C�S�L k���Ά	��f/8�n����2�Q*�l'�I�k8'?|�j���t>��BC,Wy��ٌ��CD��c�.�*y�����/
�R,��pJ �����L���Bj!����,Ov�P� [v���J8^)��`�����@$H��ӽ���)[,�]W�8��Wu-��"@N��n��x��қpq���Q�1���p�ԏ�dT!&��9n^�gs$����l�P�lh�!�V�!BI)�R0�tmu�r�P ��K�-/�y���	�k�l��?N�q࿴���
���3q4�pm�ڀuu���@��h�Q~�Q��71��7 wM�\�8tĸ�����>��I_��d�͟O!f��W^+�R�?�Y@ȁ�.]�o��wPWJ%�UM���:.UϞ��9�TZ�F��7N���7�EN�;��-�Ǭ�� 1o����}�����|��4�(�~�]ܥ
���V�׳9pEI��5� �e>�kM���1%,��O���ٛ��s	I�K�rj��ME7����B�X���I�M��C�!��-���{fn[�q�f7!4��NJD ���&Q����p|QZ�䘔��C�M|�ihG���D�a�������SK�ɉU�o�\�S$��1P�Ed�Pl
	�麡"I�v����>��teh
Y�հ!�
l�UCPv��{n^_��l���o���U�@G���G��˾�}ŷ��e�<�c��T�[m�Jk"/��v7W�	�niS�9�{Ϸ�S�˱i�i�[����f?o� ����N�B.�v�:���/ry��p���A��*��;�TLAyR�M��o0��97p�T����|���.b�#�X	y�x+�Cl�i�g�M��ƌJ8���y4ݖcy@{��+.�X��Bz6�Ϣ��s�FR�:041zhq#YWnٹ�1}1����9뷟'���O�~@K�+�(a��T��Ve�����ڠ�0�*�&v���Q����u��,��b�M�wtC�T�]=���ڀ��z����WVY�^��&�Rҁh��=]�w��+D�n �W��1��U�]+=�z����7A��ʖ催����
ēv2�ߛ��o)�?)p���(KT�+K�v2޸D�8�+!^��B�
��0�k�v�Iw-l2BI>�o�R-��^)zvwv���4XC.v�������̔���r�Tu�T��p{z��N��mZ�`ԗ����h�"u����a�A����ݭ�D�XfQ�B�d��º�5쪳]!e��Բ���-���V�mM|�ӧ�u��k\}��B��|jh��i+�����r����&��`
rZ)��HN\8z��E�4���n�M���6$ߺ�㳞��ܤ
ZZ����kdW�C���XG�_�+�B�Eͭ�E��ڹ�����QAjR�/���PP�i�~5��f�taE�`-����U�i�`��
�@��+��y=0�T�'���N1����i�'Ôdpo-q�hPN�>J�8s�mAke�0 �l�S�j�AC:��=e�
��G�ķ,�a��E�+H���Q�ں�oQ�{�.Q�h��J?qU��&���!�6��y��s�}��2`XQE�괁Lb�|+u�W�������P����g����Z�V�ҫ���z�;\x��qz�����_�X��OAgBJ�_��r�'ITb��D<�"�ޱ��1�G(��1߇��]�V�S���a�	n�د�B�ZX���3_�����4�o�Y;�Ē�֗���q��vB�:�x�-��~��VR��Ws�7d��N�<���{�*�ܼ|r������;pwZ�e�D���*WN����z:ܒ�m��9DEm�`'�_
?�!���b���F�Q۬�5؄u�~�(ƾ�����V���1<�_�ƄE�;�����h�9^n��P,)+=�ڄ�y�	hN)�as��?�#�n�k�B����r%�N%V����]	��Ť�����W�B��,{�����1���&e�7���_r=R<{-.�{��B�Z�р�#^�dC��Gl�9K	=	�\ڏ�+fż&z� n10�ۡ��Il��sؖ {�j<y���7��Q��m���S��f�����hm�!%�h�@�w�%�T2YOk���ɹQbǖ�]"]��665������O�Gp��j�0ޛz���p�c�| � �ye	��ύ^�?݆�8�H]Y�-�H���*4vO�)��U�__����F�[�8$����(�$ۄм�ũb`�a}g��b���2�g�$n9Fs@ƜóR������S��y�@������֏f�x�/���nW�є�0,5Pf�_-�;J�;)��+�i5�,��N�X�]ԏ�-\��L�aHd��ƿ����P�e��L��.�P-�\V���1�~��v�/��h��L�K���l��+�y\%�N\!p�;3����c�*܊�= r�ARz���E�1�͐FJ��<�^��<�����g�������!y�Ξ�a��H/��oP�� �<�;�ݝ�� 7�w�{y�'�ؚ୰�X��lÕ_~���JIոI��E��#ķNAR��]#�6M�i-��S���9q�������.*�Pp�8���Ϳjf�ޣ����(��Ip
֎f���:�@�ù�h���<s�E�/�;~����Sr,g�y�8��s&3t���6�@�J=e��1��Yf�7.��!	��|BrP�{�C@���3�հP+@5w�'�A�](&>q����A�xg�����6�������t��H�M��Dk��Z��!��b���8=�gނ�#�k�%M�S��j����^�W߾��2�	p�N�-_KWm��a1����,�kZܳ��G��f[h/�6�"�5�v~�����Ç���ͮj� ���Ul�oѯؓ �=����"Q�����F�`Q
L�\����-���LP�{#a����ҔH�^�753���ս�׈
7�Yrj�`����k��I���g~:��
� W�^�*�@�T�2ut߷G���v�7/�#`+�p��QX�j�� �6'��ʇ�9?��Di�DmT�	�j(�_���v��
���� 6�^c^��� /ZY3���TG�y9�~6�&1'N�qT̟�%�=��Q�;���Nr���#�j��4��ů!�Ԉ���f6��%��Y�N����>zV�x�N_�􄛣~�_��4Ν �,]�2��V�+
���!�T2�)yR,)��|�l���"����V�I��d�K/��&����x<���nnk�Zpe�g�H@xt�1aX���K ۠�|��\�%Y5D��=�J�]�Ŗ�ȹ��LiV6�#������wF�Jf��ߵ�dH�<L�vpmt�^nJ��T�D�"%��-��G��LM��Ifu��g?�<@���I�iW8��+���A���_W?Y%���;��}�[�d���5�Q�L\#Emv�ԏN�B�"x����+���9=�X��!�#��~/V-��j���9�܉���f��@�>�����6fu��0 \�z��eu#KU��[�/v[�����"���7���Ę/�6����*IS)���೻	Y����5�B�n��c��V	��j��]�$f�5�������?��"	��m+W���jK��|�ozX��Y�+]�����Dx��5x��4��\��#�H�#�/T䀆�HOaih�dB5�ݥ#tEvl��	��ɨ�d��?1�$x�;�R��57�� >1�u[f�3�l��bs�.�NX b:`�]�c��=k���Z�O����Fr?R�$r�3����@G'ݣ{ɚ	ީ�B�)x�o�u"r�A�.�f(�[�/\�L28�� a���6Rq+��֙Fj�����L��I(#��lH�.T�����q/�j�<������ᮚ��Zy6�tt���\��Ey�M�}�wF�o��)��\�6=�H��˩��.ǹ�ǲ�/��s\4���lO~Bs�/o���]�q;��|�[���>�`Xn���"ԛi,�@�8�%�Y�e
��\�=���������U��}��"��<��_�<�E�r���|�-6����`�@��`��� �$�m�ί�v��e�<?W���ѹ��ià�r�f�դ���=#�u�ۿ_;>�ѥ�����iC��?T�x���{In�p����d�� M�Ir��(���]j�riBz�f�b��L;K`0����{~=qyL�G�*:�G�&��V1mK��U�X�߬��ה���jp�
���rV����|:��
��L&
c�/��؜���k5���u�
}�vIA��5X0h�UOR�g��Yx!2��K1I;!��z����z��n��h-�0|y~�����p�ۤ$����
|�|��@��W4��^�.ޮ�����2m}H�_�$��V:A�p��]Z �`"w��.z�xe���JL|���&t�Td$�����7%ƸkK���r��!�8�BH��0-��,�/eP���%���e܆��� ��%r�B1�]���K����j���T�67C��~<M��3n��v�4�sїP�,`�s��@�瘵���*��ZL�L�r'�Zf]�5�,p"iw���Y�0��3yY���9����(��D�!Va�jJu��kA�� m%������嫏V���o4�PS�ھ����'=���'����a �I�_n�_ZJ=�����ʅ>����X���*y���,U��w�!�LK�n"�-B5�G娀�]���J $݂��6�3o������i�'�@�_�v�Ǫ̚q���~B��-���>ؤ󭂉���м��zU��� #���q$��~R̆]���@���Ѻ:ti��n�k�C��*~�*�&�B�ֳ�5�B���(��u�o㹙7�ߝ�&�É�~���ݯ�\�$�Y����u�8C�&w�^���U�Q���K@��2!�RAP�d�={�z�T��S:7��,@�iѦ�&��F槁Ub���K�ѻ�K�\�t����` p��Ǜ�����'���M���E��s��� �:��̈́�#}��ȸ����>���p3Z)��؏���Ȫm�RV2'�C$�[�&Z{��ޗ�� vF�j��:���U@g��D1
F��X`\v���i~np�����kH��BXi�.�'H�l�ZU|�r�D>EL���J�r��� �:�r]���GT�r�P}�s����c��Qɣ�5���K���,V�N>iB�Ȁ�IKy�G&9},W�ݷ�צة)�5�R!>P��Μ��U��l��B��S"�3�QY����M4���G��S�S�q�,����s>K�f³�4�������6����#8c�l���XlS���L����%,�tJ�CF���jQJҹZ(_�X���Z;�K�湫,J�Oh�2C�-Y�K�;7o���p<͹8ZWq�a���uؤ5u�A�ۨ���ii�4��۰>�U1�u�_�:?�
���~���.�1�Qݪ�t!KU'�ss> ��U-M���N��~��X�l��]]�&���u�&9:XP���1'c�\j��/f����6�j����Iz��N�m?|���rpQ8I�ul ����'x��fo!��=��3�����s��2�m���ő
�t>{�5�r�Hr*�h�g��k1>?��	���S�L&ٖ����?�J��-�Y���IƧ���"�i���|��[)�DP��(P���
i?�zQ�`G	�Ʒ�J����e`�`T�ڨ���>
eK�ˈWZ�	l�R�>5	Ϋ�z�:K:�O��W�y�[�Q֪U�Я�L�����@����>	k0��ה�Qj��h<n�$�����cX,
�=�,��[i��4�>[lǬ��x6^_��]I�2*�OY%mc�iS�T�egTu�$�Roq9�5�N���~6ͽYD�D#ïΦ�1�g���}�lZ��z�ƙ�XtL�vw4y�B��pp��I�F���5��eA��!�q\�`g>���V L�V�����~,a]JȚ_�7G�@e>� )V�����Zي�a�C,�V�E��?�� 9(o�Mx}݆��R����`���M�c��쇿N�!�_i�96��aD9m[/#sN4���nu�����(�%'R�k� ��-�?���N�H�jC�b�����V��K�-U\)-�CdTg����F%U�����;c���#)�?0��ZygC�Pm/�i+>�a_]���fm�?g�����'H���8(̛Z A�R��9*Q����e�t�P��>� �FdDJC_D��:d�/�vU;?!g�f�Z$H�ʫ��$j�{_��G�
�w�P�^Aώe�U�ݴ8B�̵�f���I�2�$淇����3�ܒl�/����L$%�efD�o�|��|�~B#��3j/֝�o���X-��j� HX'�T��J����⚇U�CC�H�0�?&�LӥnH��Ǩ65PM�x�	a�Gg&�+c��5Un)�)��4��U���َ���Z�!C�+^3;[_,��M��t��s Ǥ���h~�Iux������m΂r�b��o8�:ތ�lKv���(~��J�b|����5{U�[4^޿�G�<8)ځ�M���XGH7+U����/*��Q��K�5\�!k��Y�e~�&�7�Ӡ�؜K����S��O���O�K����0��y[ͪQ{����?����jו�;5l��{�q,6:��(L� e�!6��:�"L8*��ב����(b�x�&)@�Cx��'�-p�
y�=cE兀H"1E\�V8(� "�h偰���]�a{�h����|����
�οT����v$��۝�p��w��"�*e�,#P�j�F*Fav�/{�$*�-�|�z'�)��1zW49��1'φ�q��^�s������Y�)�%<��2#���;���-�MH�_U����4�z>X�K`�8���ocBe��G�q��~�h�x!�t���k��>�(�v�w�����=����r[_��uE���
�������
Qv���,�)+�r���g�lf�T��;J\��r�z���<�y3[�w�^+�K�Lf�;�ei����'�t�Q�в����®6 WTaDlFN��[öݖ�-]���=���K��dȈL�û��߶�.��B2��lRʗ&�N=�i<�"fj׳+l7'���a;�%v4�Z�~	�	�m���~�pa�f٩�i{ܿ[��T�^#��BKEk��]@���&IR��o���U�W���s|����̵��|D����o�	�U>9�İ�Yx��{�\^�u4�WW��"��?>��Kp����%�,Y��;�O��K�VU��D=_��s�nEm* ]g2��qg�s�V/g��"���M��ǫ���|��L�g4�����Dݲ����5��$�?\	1}S�W���i�Lr�*�)β"�X�Y�� ����O8#o\��$K���B���ُ�~�i�9����n�#]�[�!:��:��ܳzT��0ӻ��H�1��u�4]���h����3i܀JN��
@�?���Bb�l!a�Ri'�^us��cq���W��Ă{��P&�&�?qNY`y{iI�/�99���
�*=�����S��dx��թ0��E���<��z�35(W�f�?y+1w���<H�G"�;�u	�[� |�$�%���`����gt�8��'q�şJ�Fg䗿��$�kƦ(���)ܑH2O'C�rr/�f.��WFT���`�/Y�PZp%$�c�ugHV�П��%'��s�)8)�rokcv9'�MQm�����g�N�>P�F����3r���������Gd�����_��@�����E a�s�3����5f���o0h�.�/^6Jy-�vP����w=?A<�Z�.܃d��@ιX��E`z�v����Ү�q��z�I|��Ph/����Y����<����.!�ŧ�i<�����-��]����=�{�v@�q�5�ȰYs�N�|�5�2wIӽ��9a6'����!ԳU�"H?��O����	L*�x�lv���ҎXH$߅[�|���A"�Y���6��'q���Տ>����t.�c:�W�i���n���R�>�"R�EB�2�����UN�_�bςG�֦�ج�b���Zo T��SD�Ճ�u�ڬ�J��mݙ�&>������柙ԐZl��;Š%l
��cYA��5�<��B:���#������Y4U{��JÒZ�Nd�)A��5��s?3��S��#|�[{�*�Wf�߁��{n'Aޏ���- ]4J�G����������^�(����+;׹�73怏E����&���O�#p��J��p��4�� ��P|�����n��Ա���4��B4d��;SvU���qV��[�oN�}�R���NNEܥ�{�b�U.Ἡ�m��-q� #��9���6$��n��/s���_b�x��c��n�(�����9���v(g^l%x,�خ����'�S�vs�v�n:��������	g������/�M�马_�o�:�U���1Nh����]������n?���%Y�X�!el\�S��:��H�ko*��������	��S�%�b>]��ja�9�[����[صc�z�A��ce4n���N�[����� �g�;��ǧ���*��^d��<�b�(��%�3�	��zJ�<SIG�x�������YM=+m�����H�3��ud��wE���R��ǉ�d�C��a�H�y������{xb���@���&d�>Z�{��88��#� EQr�d
�SSy�d𕍞�>1C������L%m�s۹5�1x��6���VFk�`)n;15���M�&o��h�/�6�MGE��ˌOp}%�.(X�SX�Z,ؿ�E���n}.f;W�̞�%��� ��Ԕdؐ�M� "���0H�t�������Hj�٠�� !p�C�0G��.d�-�]��a>٘BP�{Y a���`��)�ݚ�=o�HP���jôm�=�K�B��y�=<q̔��I�q�k��>�s��/�䗴�ќRh��bҡ#È�y�#l�.�����%�4��+S�W�2#�q�/$#�<Ħ��iA?!��g�ke�1�|��g,hK�>R�RM����$��+�U���%���p����w�/��J��{9FI�X�2��x�0���Z�H!��fB9&�F��_(Ϧ ϖ>w:�*��CY���白�x�N�]B�3��曩�e[���;u���萉��y�����ݣ�,����>x�]�ce(�qh�8�~�h��SZ�h�]�hp���ؗ��C��y�&�/�7��\<Ic��-~������Xy�BӺ���g�0���joA#A���ܲ���e�x*��u՞�|f�|�J��e����aS\���MЈ�?!��M(�%^Fk����Q9Ҧ��5�������v�P�E��b?�p!�X��2�t-�k�bv�� [My��1G��ڝ� I����S�An�<��̀W��H�J��� �]e���n� )׮�b=�ϳ`~�9���ã��:���h�b�\�M~1^W����R��^�qm@o�5"����r�7�|KW�3}�K�R��=�A0��@�����a9��ZK�ɫF�K����d*�G�J�	�~��u�9!ӎG�衍�!AB����Lԋq�!�h�D��2�jB?N13/��,�����+cK#��g��(A���6�����+��ukZ݃j�h��@fX'�q`��N�K����
���GYN��D�Z�3!��O.�|��֌q��_�Y���������=�H)H�]Yu�w��>���`�^�R]�����|ѿ�	� �܆�'��z~��@&R��!Z�A���	��5� �Usfm~�T��|�y���S�����8��ʚ� ��� �ɱܽ��2�@(:��h~=eI@�e�9.(d;����ɿ�$P�\�����ic�`�b�Β!<��A�q����8+���8<�n>� Dr{�)d�r�ޛW�A&%ú���t%W����zU�ۼ�ik��0��[]-��?G,�U��/A��P��V3ƥ�NW{a�]���un3# ���gӱ��2���\U���u�
3R�ş����ME{����w�񦺪6�P�J^G{*��ǅE���q��|5YFY�X_����┗6�$Ο��d~�I�A�+ �uV
��/ob���:PП�fd��\BN�
@ZF8���P�+�-P��Z2��1��O@J^��^���56)c- t��ڌP1ɻ���7�R�Q������g)F;w0�O��R�AO�(��鏯���׬rO���������v�D>$J�X��u�C�A1�~��)��-[�)#5̓�=��M����5���U�Z5F�!>
6sn�A�:{� ��#�m�*��V��I�b�(ꨖ�w��� ���*E��z�X�vW�l�/"�j����t��BA�F�R��p���"�WR���%M���G>�1�%�h��&�*bU @T�6P����zf��-��܈�1�G��o&L�Y�=����nH@6��8!�ɉ 2r�
G}��T>�r0ڏN���-�w�zu�
V��,�	���&F�ԕy���BO���Z�M����ř���S'atb]
�T�����+�����q�ز��(5n��J;ҥ� 0 ]�D>�)d1����#���Q�>���F`�>\v2��3_ ���}@�;�K�4�Ԩ�b�D���5�g��..��жbEf�J�S4O�,���eg�#5���k�#�}-r#|�[�?Y{صb>}xb�GspqD��5�k@�b�d4bj�V'�x�~�"��j�l�u�.��Δ{�;>�z�iQ��!u�Ld���W�݆ka�Ñ��W��v'VJw'2��d�\����_�΅ޕF'�fܩ�P�M"0���� �yٰ�B��t	iş��3���~R��-�Y-��j���iع��-��c�1zΪ�F��*[�����s�E'7�[���1��Bѣ�GH�d�2��:�����f�uk�q��)�c?�u��x���&y� �EB��UV�z_�~~f�Y�����>H�s�v�ZRS���h>K3�b��ё�FC����< -��V���b0�B�ée����%���nE�i"�Á����l`�ݮ�]�h��f�*;	8_�9�[9�'���9O���@�N?��zݼ&Fa��F/2�܊Mƴ��9v�}���W�>�-wv�T��X�_эbD�L�1;��1���v`Nj	�I�xa����Y�H��Q�+V3�;�	K:�[�B���O���ӎ���ィ[��
ވ�2ئ�r�S�(ʝ�U��m5t2z�]�cu7�z֒x-�?���y^$�GC�yi�������k_���^�<m�Q@�	�#@�<���BT#/���ࢸ�So3w���yBp3'�i���!˘/��a�M����C"�Y��lE`q�̟!8�u�m�%dJ��>~y�w�#O�٥�vd�������sL[�����\J0��X	A+�Ho����I���)����'n?��[6��M7�;�k�ICI[@��-���P9�~F���@�Wy��:aO͘
��h�sA��g��D>��x5��"bU��)	��ʷ���T�x��u��4H�`����y�[u�Nu�6��|��Z�U�(B'��2�k\;H�$�w҅P�mt���2Y�X_a�}5�:=�uF���^ܯm�E�#?��
��ɳ�^F-����/�U�#�!�}<�[�v�[_֧�"������gB�d�U��y-$K�F�ݧ�#*|k2Qԃ�
��D32g2@��T�P��9��c}�C��:.�|��y y��F��4�6��?�g�֥F��H&��Y�]~r��0�����WY�����~Չ +�,��8�����+W�ϡ��Md��B���/�Jʹn�)�������-f�a)�g��^����i�Ú�O=TYoz"8�! �L�~�i��� h����{j��n	1������t�P�.��l]��HiJ���X^C�Z�㕞��L��:�K�Zn��Ꮠ����Z������N�dt�fO�F7+ǯ��rI��2N��=�i����������dDM ��aC��!�cs�4pe�c���D�>/$1�|����Q\1�)�s��럺��5F�
$���ڲ�5�p8�l;��q�>:�&9JuEq;�i� ")���Z��#�=�Y�����7��ad�]@Ā���X��y��ā�Ȱ�!J�һ�0u`s��*Hz�iUK�H�P�>�㿽#��҈�����ymqM?��^�E���(^���ർ�|�EϟOY�yi��0h��o���
� �E��(��*
Ai7hz�"9M�/qE�3U�mdFմ7�I�z�K�z�k�gD�kQ�w��FVD����v!*5�cA���H
�u]���3�+��Dm�n�j��n��q�x�m�܇�B�a!��� ��Y�iy��fg��`�3��J�J�N���{T�#}�o�}:��lH~�v�4�Bʤf�Lxы ��6ŵ������yB4���N�=!���ݥ��޶KS��ů��U	�An��n�H�D�M�G,K�{�U�$�m�?q߷{�-i�EUnѩ�xb 6LI�=�6|Z��Q nh<��iF�X6�_�c
��[=}PXt˖7 �5eX"= �.g�
y*��I ��x��������3��ִF�HE��������a%�c[;�c0�2*���>�}�[{) @�s��sX!G�׭�RW�Ű�϶s�Z��[��TɲӠR���nO��I/�1�)��h�E� 3YP����7�1L�b����iS�DT#I*�j��܌�l�-���v?%U9Z���Q�+�MN�%�h
#�2��kI�6�[���t�.]F)��4a�����ۯt)�����[N����c�$S��Ѿ�}�-���v��Gѐ��P$�����J�����U�����uI-��a���#�ݦR�����e���C��^I���utcgH�l�"��܂L/�䲣���!wf��U�tWԅ�S8��	�-�M����GnC
�qi�5������-�x�P�w��a�{�Ȟ��OKm��� ��0_5��ųKX&�]	����> ń�w�kqi=KMBx�A6b0��K�<E�p��v�ɥ"��{.�zT�h�jsޱS�o��G\��`�M���:FY�1Xv{,�A�|����&ZFH�6>�޵z�<����w����W��<E��ǭ�D����Yp�0H���T��8݉�:���D�{���_�\Y������0=��
��ؔ��ϥ�����<sjm
�-X\�j��v�Ke�0���T����0����j�*�"k}�����m߻	E?U0wd�� �i�aIk�pQ�n4��3A	I�F��1��&������r�k�M�:�_���X�N��;C}��$ixy>&�~�)2�hHM*��ə��@K�m�y�^H5<�BqVɯtH�]m氶�&K�K�솄�bo��'<H�0�0E��j�������v����H�5qQ���.����p�b;@�~0��#���u�舠�"��́w	�"���V�4?G�nO��|r�U%���OQ��ED�E�J�+�dÙ~W���2QMv��B�l+D^dc$٪�LKŮ�L����*=źd}W幅��$Fo�dRvap:{G�-[/���ʏ�Ұ���h�=vv���8}�tG�#����2�0����{���;���Ү+�?����h��u4�#�j3�'2x���	%�(��=��'�D=�?>hwf�D!}�DTKRF6=ϔ��]b,QmE,�e��ٙ��j�VB�5��`;G�	�)V^L�a����E��&���e�
RJ�%�[���1 Q��d���)\gvz!Jރ,���q3vT"�.��m(\���W�p\�G�,f
{�}/������+���u[B}��l�`�C���G��P��(dy�r�i����Ȳew�pR�����������,������Ey>�F(d��o�Fa��B�_�:����@(uO�>���O�hW[�n���=bo7�0�"X�`���*�hn���+)���zv��moe$��-�,��V�Swt�r��h�F��(�A�U�%��'ڥ"f���S���lJL�8���[\	-W�V�@!���ök��?��N��O��1��U�O�
�̖.���g�^R­��ƚ�MmMP�g�{!����t��_I�_��K�n�_B��L�.1�0!��_��}݉as��}�w��N���w[�5<����<�#mÕ�_��z卌�]N��T�G�ꬖ�`W�:���@�S4C_�q���k��O)lӲ����lU����)�#�'n�'1�bȪ�_�u���=GV�}]�����%��y��Gr����ݴ��yG�:���L�s�����Eۆr���qʓ��X�{�}�7yF���Gi�	D����_�U�x�Ƣt7���-���9h�6N�3RK���zӚ��Z��=E�r��d0L#�aO1�ٸ��6�T�Y�]+1T�̥�d0�i�y�>h��J��n�uܗV~�4����1�=�"C��a�ͭ،��	���T�N�?�3S+�a�JD�X�zx��AԒ}>�/f���Y �tV���=.�����L���B]j�OYH=��8rR�u��V��U`���D�	�@e��D/���h%w�1�$�%��r�8�l�}���,k#�L�SY��pQ��"gL"������.����|�2_���E��c]N�5�{H�)�Ik��m��*[���\f��ja�Ǵ��e�/�U��3?H!�]�S��~��5J���c/��S�y�F���=Tap�x�T;}Ɏ��+�}W��N`���у$�.���Y�
���T�n0�s�)BZON�B~�#����rԥ�&�au��>Sy@4��I��͕�"�_@1�\
�B2/��P���{X�,�i��9ô`�2��G3�q]@)$�T&�hP6`3��`��ӹ㏉p���/�&UQ y~�)[%[Pr�ԉ�F�b�j�ƵH�>���x�7�%.�j�����+q����h��C�rde��9;ɽZfS�p��*�S���s��r�����!�@��b�.(�Cw�j���j6�4��%�{�Nr�I��'9�*�r)������K_�� ^5�U_�da��yۄC��VfA�(��<��4S��46�+���G1OYB\��Vc�c�w�}��~��Hy�>7]f���Z�4 0𱢉�`/蜫��C���f��#��E���Z�4/����92tS8',f��Fn�M�ܫ��W��Z��+[�m��2Yu�%�5ɮm�x�Y���?px�g�B5�}݉ ݦQm�����J���º!�]���E3���DH���:���$�KK���BT��ʠcQv��螉:���n��>1EC���5�m������Z6�M?��t�6��h�dbc����o=?y�٪��c�-�`45������d�&���6
�o	��5�<n$�$*�Ke��~���������m"<�sg�"W��_v�J�	1�� �S�9��u/�u@j�i�L�����6Fh�_h\3��_�����Q+
E�~l�+��Q�B��� �K��]Jfڷ�h [�y<H؁��A{ E�U<Ӎ|;��#�c'[��q�91�x1����'�}ڌ_�Y��A��.!�&����K��g��U%���^x��&0.�V��[�'	�Fe^�,�hgǽW]�����Æ��6�"��|F�}$�Zʙ,j6��O`AkY`� Hk���Z�"Kݳ������,.[�h�������ߋ���EO��X�X�r�3�*�ww����q�}�Jpź���S�#�����%�����\i����\��EJ����`�U�
�l��R��}�8�.�����q�^�]�Dt��$��M ��L�4�r�e��Z1��y�[;�𽌸[�N��1�P�'��$�(��a�(��o�E�+h46U�t+*�`��~`�V�V+dHA�Y ��z��o�JȨ��,� ��3FQ*\M�#����j�&Ȭ<�$ONP��:��� ���(�7�^t�T�ޞ_� �R�mM���z|�S��,�mJԸG��BK>�\B�%��9�d4���{z�=�	8� #qf*b7rXf��u���6l�N}jE.�0���r�	0f��仏oʘ�������l��)�X#�d=�4���<��Tܴt/\�!�'dv�'��o�^�����]��e� g;�"0{���s���r�*��T�M%�'d���@݋~No�/��"�ot'槢��W�wՍ�`�t��]�|h���^w��i��mH���m�}�y��v/c/-�:3sҙ,�� >;�|Iअ�e�\�?~��:��O@5~MZS�Q_�C���[��%]����no�Q�=9K�F�1��՚�uw�_����6?�)��ﶩ2LW3~ �"űN���EK� 9��gu�=��s�^ɯ|�EX�o�G��_�Lj�]||���%��zVj[�k��z�A�����N�+�u%h��ɘ�+}�LM{Ch��Ԅ� �A�jՍqr�###�N�e4���d�O�����
Wx��K��N���/�=���[G| ����|��B(=`����5��� V�X�|�-�4jP�g�9��R�Z9f�VjY[�P].�7��:1]1=����l8f����CETED�%��
�^��S����6jCcB���H�@<�.�Іj� � B���|��YS���R]i���_|�Q��!�t��D���%$Q�-�E�F' �"~A۟�Z����%�$�C��^�#�Q4r�C�yP�;��P\�1��r�_�����y�+�
���%�Uy�g<�x�$LS��6���;g�U�aM���t䗬�ͤ�(hpp������]����9Y�7\f�g���&A�Q��LhSϟ��܏w��ve�U�e�
�禞�G���.괥u2`���i�P��Z��e�;P6��'�~_�q�5/�Ȕ���68�D�>\�U������}�
M �Ja�^��o:����u��-_%� ��*������?����CK������&���ٗqk�|Z�̦(%�!�\1=Y��o���K�e��Li�jFC}�:P�Y���3��Y���V�8n6v?�l���	�sCʸ��_vFo�{��^gӥ13Ï�DB:��9��"& ���CPJ/2��zC�@Kݢ/�Y�(y8�'WN��%~����o^_���M�R6�D��3��vLM�-���c��o���d1�&���9�o��J�j�����"���EӢ/�D`�\_=^Q"I*g�T��>�[��)w���.aK�!��"1QvB�UC"�AL��h�_���NH���:��J�q���Ѝ���	(�(��э!Q��l>��lJi��A�Gm��[�r�OX��)�8G��۹�P-A&N�+�u�=��%�P(�x�7���V2�]��o�=�Qr@L�7�U���a�Ƣf�^r�m�W�p�~�v�*����k-��c�`���ȣ��Q5��?IA�/�֊k��ף1�;�8�h;DL^:�X�:+@7�`a#�;�cޤq=	��9���9!J#{���+�d�@�ф<�!�����	�:�:�gr;3�����d�O}���[���Kjf��g>���5� �蜶���O�Bo^<���0K�f�I6�kds�$���	1#��|f=��� d^Z�D����*➙��)\>�{Yo�a�Ө-��+������M��f�1�ީ*;7�!�D��9���1�����~7JGƃ�ڹ�j��#�y;��4���D�I��nP �u0n�؛t�RZ�ϑ�� %�b��Ou�Xn	��;��&��2J�/��}���uܭ�ᯌ���/7^�����L��ܹ�-ϻg��\&�����!����!%oX^�����)ns}�ȸ\Z���+UD���VM+d��J�����yq�k���@[M�o�OX|#vg�B��dQI硃F#<0JL�l�`�mVܮߦ�b>����.�sT�U&��^ZU���*��F��\Uܐ���Q�M�� k�ڋL��aB	HC�	mM@�s��N�	�s�#�h�S#��Ġ3Ò��	O���O�i���LPX���+-n&�p�.  ^��~3��F-o-�8�m􆲵j�%�6����a�y��]�V�\�M�{:�	�\'m��bО�����GDd:�!��y(��7h�4G�(�����[u�����1���j{�B�Ν�Rzɝ[#���Uյ��-oਬVF�u��w��d_�	�����|D�� ��!b2ь��ko0�&2!4�\	�1a�42��=��JU�U�|�&28h7�V)�����1>���C���r�α��ީNB����}�	��y��Yf�G��ꌴ�)�ں$���,yˌEBFG����-���	��J ��.��u�$�����Qdk�x�z�G����ܢ��?��)����yv2��!ku8�p)+Y!���A9�4iT3I'hs*�<�k�X>-�l?���N|y��*����ę�F��"�_)L_���ctNB���F��&��m��n�� �U�j�$+��]]`mSI_�_��[������љ3��EhY��Lt]{��Lg}��Ǯ,��ϣ�%��$�AfaQ�V�c�e�7���U�a�������;G����p��;k��MO�c5��3���w}3���X������t�U)�
!1q@��N���v2g��{ʖA2V�"�� ,��(zeH�|μs@�����}�U��4����/	�~X��~��6}.�L~sbgR�����n0DY����6M�̌��Ģ3M���	������� �9�;��c���<������TC������e����$���~s}ݝfw���:�x�D�A%2̒f���݁-��� �7CF�x�'R��q�B	�4�+yf��Zg/"�{"0����&��˫� ��h����C�I�od����N�0��w���{�+����=�Ьv�|b��@�Q��j���F7!�}b�x�Nˡeq�2U?^�M}��]��m��KL	�ƔK�IL��r�PX�Ɨ�	��7(���Q~��.օ�B��-����ـ�?!̈ε�5�2dv�<o�>Gu�Fy2����Z��
<��3�%!��.u#�`��Z�p�1r�G�rL��	��{4 t�N��R^�Y6�k1����R4bh�(�𐁉�{e��`�� ��.��I�%�F_�o��6pQ��K4W[V�)���;G��k������J8p�+�8��p�R�c@���r����HB�ӞB�gx����7�LV��n ��Km�Eo.|��+k�/��,�e^F���|�^P�X��Q�(��{nv�-A:1݄���n?v	���Spd�W�j.8�ovT��>/M�!�I��yzV�4��Ath�E�`$Ah���T�P;�%F���g	%�O=]Lj�d�ך��P���1�Q��xԵZƼ�G�
d� ,:�r�^D������� 5u���n�A'����B0�*#� V��<�[5�UpI���W�"rLQU�l�ƍ�Dyғ/3 ��' .����}d��I/�z�~�r(wN�y�Z�ed6�2��B͸E}��a��;N�#9��9�ebw��ߨn��+Jf��%D����}��1����k�IE'��e�nGз�1�`�ͽ:'�F���9ߗ$&�yO<l��d���7�����V�9,����{J�
V���_��_6�):��)(◒D�ۃ����z�����ƥ������{1mCŵ 2�r���H۷���HT��=�*�;������ށ�Z��+�#5����7I+��c��+�)E2����6��j�ܟ�Эԅf����2V�C)>ShK���c.|C;�Ye��S�FaT�t���D����8㒏�8yJ�]���y\�2�f�����,&p�Hj�|�Gh��R֊q�rWl큷��xef2�����9���lD���oEI��k���sn�C&ZS�c�����{�<-ނ����|Fn�����K>�&� ���4A?y�0I���~6T�f���ȴѻ���gt���L��?�~��{ٔ�~m
��J�k�(��[7_���`O����4�P]MYԀ�Q����޽/���M*���`�v�-M����=a�{�ӟ�x?���hdl��CA�"���ǋW�ĺX�`�%��gYJ�O`qB���7p��k����ˎ,�����k�sƴ*X��+ ��Zm=K�ǆK�]ǉ7��Л���a�� ��w�zM������ �$?�L�>����]�L�"����~��e�T?���Q#w�cj�) o] �l�%�Bb�Ni���"�j�Ǯ#���#F?����fm�s��%)�y���>fw���e	�v̿����*��ü���޽p�о	����3\�܅��TX�F'�@!\�u��E�lp��E�0�c��N¹�߭& ��Y�Ûx�V�,��#>a���'��V��|@��ۑ�f��F���8q8��8�4�T�V�m�D�$���4n����W靠���Q��MN_MVm� �O:��z���s(6�v~)�-���Y׬�^1��&'=�y؞x|�TKS�TA�U��۱a��0��n����)�=�]n�Jm���K[v�����౥������s�zyr���X�mwOr�����)̵%H���Y�d�5��t8ۉ"A(��UQ<��ؓ�u�`�	鶺>�l�d���ڷr����*% �!v����=y�h��7_̮�3腏BX�C���P�z\;�)�[��ɗƭԣ�"FH�����s��֮<���,�����?�/�:�_�0B��B�pM�d\�*�\������[Sl�pV�@�ؕ���Jz�)�����t��%$P������� ���Z���p�'�ї�a�gU'M����c5s��Q��ڼ���3��9@���j鷥W	���Iu��������7j�9�B6*J̠P0��(��9L�V'H4���F���u�ޓbo�=��e��MtR���+��V���O��v�N$���R���}�����ym��ҫi��IŇ�ܚȱ�ߢ�K���J��ë�X,0�Q��tLXFe�nL�����9@���dIڜ3��ã�U	{�y	�Y7�OO99�_g�)��h������E��c,����Z)�G�CQJ��1M;���eX���T*�Tr��K	�R:a�Y,�s�S����\�b��[oE��y�|'�4��B8vf�V��W�. yF�91QR繦�m�zy^��BU�mWML�q��ǌ���^d�n��^"�(S6��w�}�f��br��0R�Y�qM,��B�g��6������V�_�^��H9|�����s�}ջ�����E���5���/0�����h�̄,���<Q6nd}AQ	�����9�>S|�7����X=?�3��l�"q^Y���g�TEz�R�uW�+| 87�ڶ~ǝ��i�
���4��&�P�1�����2�y,��6���rF���|K	7��4�����U����t�(@koC�ā��@���ΒT�������4�$���r��Ǚ�H书:=�$S�>2�{����*��f�g?BpF��Qݐy	�~��>R��kIj:xq�g�|�f�a�Tu����6���Ki	�Zx)���D�<w|K��x��x&&+7x(��j>h��sџ�;d��:a�wܐiy���"�xq,ၜ񴜆[��F"H��Vm�>:[m��M�PZg�þ��2�n3Q���ל&#��bKr� 
��t��ƙ|������|��Œw��+�.,0Va�Vŏ��j�����u����Gb�]��U�嘂/R�)�� �+�rƕ��$������=ֆ�pFLD�}l�ݣb~
�L�.��|�k3��;$�m#C�q(��*V����_,:~���+3Tx9����:��n ��ޣ"1Ô���2+P:j�śŏι��Ŝ�r �O���>0��7��#�gwe$��4�l��ꭣ����˟|����­I�)��z���W{,#�M��u�MD��(�[<��,`�;�C/|�#����P�|q������Ţ�dG��NEfwS�9�!*b
���M�&�u�K'f�9�H�����+K.����N!��<�|�c���5�t���Gԅ>Ӵ�Q\_�u*!�,��5z��.�hs(_�#�E��>W�"�׫o�c��EN��Fɳl� Vp��Z2�7�~9G��41��F���^�Ft"pk���hq�n��DAJWȃ�Cx�ρ���m��ǿw8�����v<"����eW�m�T�D�bLy����ާ�#�#�A��<F�b���燸c�_jk24�N�cB%r�A����I:r.ד̲�&�k�D�4�(����+�lVy�M���9�fC�0 J��;�J�q=���)$�JD�����^��?<�?�אX�&�g�A����O��2�Dc��M�.l���^gjg���.��.�_�1G��U�b��j,�����eT�QK�U�i29ޘc�?�C(�DGtǛ�B���
Q�Z&��^O�A�!! o)|{�E�j��h�� *͢as�< o&T�T�A3�D��1���A�G�M�*+-�ڳE�b=�.��.��x^o�ՋA�fB�x�
��EX��,+�z��1�X���{�rg�2?C���g��O��s�l�4�}C)!�)q�&����@��N5W��Xs��	�R���y�8���6����\�k!W�D�_�_���~&�Yk�^�,r��#���?�,g{zb�G��L�$i�~�l�00Y�v�aa� {��fj���)�F&%��@��	�^���^"�"ػ������r�:��b
hA�]�$Mu�bN����	��t�}c���3�����aR�i�#jR+Aǫ��W
�U���Q��]���+R�9ޗ��(U��0E��s�,6��h�Կ�	
%����m��F#�U�2Vb�12���c�N�l��Z�}��z_b���N觬Gr0h#I�bx�!=ޭ�/i�e��㏦*��iF}�5o|�������[@bLE>�צ�
xl$�&�~C�R�6�6~i)�]��T�kz�����������hH�i7B�����c�bH��d�����=g��_�� V�9rX��hn��K��ͫ�
Q�B<(����я��XjZ������y�+(����	�ا*/ө��X����_nE�=��QD)Xz\��Q̇��i�A-S_�0K�8�&f���5<�����'�ZM�#�� ��Wo�rPz��z4��t<��c^�ק�=a���"nFQub1;d͑�!k=�2 ��X,�g�(PB\���]@�?��x�H����H�x��kF���9��-_�&s���<N�W�����u�n�$�E��m�d�"�� �·>f��h���y9�����g�*"�'
@x�(�/�
���E}�	�+��Ώ�U	e=�\��k}Nh�(�0P���KJ5�Ue4O�qj8Y��HZk'�b����ɓY7ղbde�^i������	�ʅi%�jI�4��s�PtPi]QC�]�;T�x����z�!jU����H��(z�=9��-5����n��ϡq�����ml�pE�}����/Lo
ʻ�[��g�3 �3Qu��|VR��:S"s�-���ԹQ������O�fː)���Al`����C*�3�vЇ�0���2^�hrZmd�,�[H�%�Vϻ��1+L����ZQ����qä�噕�H�ѷDniQA��oJtj5_�ӧ
��.k��[�wT�C��Y��.y�e������dl�9���������#
A%V%u�|�˩@V�b3��H|0?�e�<p�� ��o��0|��1�A�v$�eh��D�����{{Q;;�%G�z��}�R��L�t�Ѭ�E���"]��ƫ�X ��>�����П����.f�36k���'�(<�� ���ڋ�����E�:��>_e{���Ka���!�~#��8����ޕ�'L�KD�]��b8��瞼���b6_�p����﹗|�W���&%Hd�G���`��%G��Us�u����#�����1�&�3l���'���לІ��>�(q���ʬ=3+�҅*�J��#���ێ�<:G�6�x3>���B���ե(-j,/
������a	��3v����m���F��s�d��5��w[�RK�~o��NP��=��2Dx�s�p���.�$j"L#4kh9��=M���c�o�~Q���yI�����'��I�R*EW;�&���@΁�'��e{ێ��=X��qɊ���UHY#��"v�+;�*K��S�}2{X�?�3���ߚ�.gD/���9�B�.K*!Cdi�'���	_8�Wۼ�����4�q�I+��W�M�7�Y����)s�� �r���˚��)2�d!���)pbW|p0!�1��Dk쁧5m1;,���L�(���e�p����'��#�s���-�~��C��7�l��~�w�G�T͡�"KE��W
[V9��
��nD�q9 ��("�0U��1�E�}��Ho��œ>�E
�=�/)����\��~}�8a����nė�N ��'� �.T�NȨ�Nb����ɭ*y�`�5{-he?�m���a]V�>h�@2-i�{�-k�[�
�s�r��Ұo�w�\�Qs������FHq�����n)T�w���G�?ڭ�ې��2e$��jc�� ZiZ����%L3�X{�=΂|��i)��d�{M��P��F�ߠ�g� <�+��o�a�>;oϪ��1�d}YzP��l�����}\JD��Ѥ�\�DSE0O���?q,��Ȭ��X�r����mA �����t��&���I�o�e�������X�m�}Jϼ��\����7-t1�Ȕ�l�Yp{N��R����W[U߅������=iޅt�լ�&Y�(ߊ	f%]���e�J�1�+3bo������5KK������Ol�C�:�����~��6���v��@@���u��������I�^V.�x,�'"R�=a����9����0�F����Q���~�e�9��r;e$=�t���ڲ�/���q��7��@Gt̕�����n�e�$�^���+��9*�Ss���@$�'�Z��PƐ�'P}�����&>�ks���O��ֶ����[�	�0�����������z�8���� u+����Ȇ�jpm�~^�^��!a[�i�_�H]A.d�N��+�L���ҡ�Y�dE�x��r�6{j�l&DD��_�U/�)!��,�����
�M���?C�������D�|��a��8CE��
���Nv+O�����V}Bw����~�-⟱�ӏ$��)	���e�꼛1n ȉɾ���I ���թ>��D�Fs��d��D�K�:�_ "�L�ξ�x�~���P�e]:7�Z���Su��x@*�{������sm�%ɲ�J���i%乆�턐��pٰ�ث�[��������6�2[�E8����縖5Q��TN��j�tFQ��Ӭ) �i �b<�2Xc���/�c�J#�5��E��$�a`�������w(�+�ƊK~Y����gL6&~���(�lL�웽I2$4dI��gDM��q1fB�ԏ@�тL]4�S}�,p\����I�gTT\�囷��Y�g� �/u�r
�ۭ��.ҏȺG7�=`�&�H.{��i]���f�����O�-]��-�Xx�:�T̡�/e����<��ʔ7����`�����P��:qϷi[�ָL)�Uv�=�Lq��+�����3��1�	��0����tcT�|���K^��-�V[]��g G�-V��V�����Z�۱r�����g�|gBr¼G�6\�a���U�ٸL���ʪV��u9M�U)Y���O�K�����vB2� �m>HF�R�ɵN�Σ>iy�"1$ī��B��TP����	������k�[SwK�u����v�.Yԟ$���]k@���i�>�X�n��/����"A��&���z�Vs����4L���ĩ��%R26�*��+��3w��y��`X/��ͭGXLT�A������4���%�;�0RH��Z�4�H����s����2���qy�J�̛g|����!�L���1�]D�$�Ԣ���@�ʊ.��'ِ��/С�F�[�ǁ���R��ft�?1 e{���J�����{�7�^�A^�	�,��)�ҝa����ֶ�X's�i�����@���p��W/�K�v$Ud@�-�e�Y 8�0�.ʌ�6�PRK<5;:�(��j=`��'�l�����o��F�[�e0nHK��^�)]��`=�a�g�6��5�3eر����K�T� ߍ�����xm��D���C	�9�x���d�
��j���Y=���8� �J+(\��&]�7fx���g��.���b1�YeW�h��m�����s�kB�f��V�B.�B�������A3IJI�Ipf%��s+I	[(�YH���T����Q�$%A�y`�����E*��q�K��Pu��@c�Qs	j5�@�K��FBK������y>+gܰO�=�|/����\l�;0^�;ְ��Y�������g7�l��~�V4�E���q���咭@��Q�W��FMX~߀Z����3Y���h�Jv��b�XF��P3_<q�-�ϩ���`?1���hfd:�s�bc�KCu!�r2*� (��E
:��
��dR��^�
ʅ;cr��!	�����$����%��1-i\��tj��Q�^��9]֪Q�zC���7��
m��>'��5.�%��?g���v-T��6��^�(^2�ou�
�G���7e��/	֭�Y�y�oXL�
S�v;�*oW<�Թ}�(3�߷�n��p�i�O�_����r2�x��ҁ����1�1=��q[;=��?����d[�ªl߶�Sa��W
���ǃ��c(B�>5ϖ$���D�b`UR@?J�k�9F%�ԬT�0:�-j�$kG	���w�EJii�=#n��~�w�iI}.��]LIU�V}�Tg*s�r�_o[�FW׼�3���-�{C�I�^�}#������]�:h_#S�@���e�.VηO����nk���FJ�Z�U|��>\b���8F�
���� ���
�"�㗼J�5��V��h�����N!��\�ࣱ(�
u/oBT����5R�pr�܂�f�f> 	�O�5��&I��-6i���[R����a0K aG�8�E�*��$�{E�Y��p��K�}��y�̟꣨(�w��H�Z2C���ۨ���6b�~�+�G.<��+���m�nK��&G��9����iΌ�๊8r�i�	��T\O�f��	��wpMQ�^#͐���6%�z�'�E�ǀ,	���E�)�L�Hd$P9Ƀ5�S�b�Nm�'vYJ'2�ۣz썥�z��oQ[9��{�,8f��@u�����WxI����-yCF��ʠU=����Zr���!ӽ�7v�x,� �rŇ�u"D�`
W���g@�Ta����TX@��`��1S�I���>�tN̩��)bY�w��2���h�)�`��Z#�{ �y�`
>J�v,�=2�n�}���^�D-�a-ݰ=��	�0DuL&~#���k&�$kl-n�#��?P��D�/A��\]M�^���y�$�C!`��(��S�ќ��e�$mV1{
���IcOԷ��cw�0S�)v��vd����wB<�\��<6��އd���nʽh6[p��rWt0�O݊�5��Zம�;�i����0M;�-��o�<990]��D�-�&���[!�3���>mƯ��z��.�"$�/b��~��r0t��!��_>�8���M�nU�5������Ht:�����S}��|���iX��nӯLx�O>�tN�/�p����	����ͥIJ���/ځ������+<���2���>nQ.ܼZ�ut�{ָ%as���- 0|�H&Ea�툠[q���r\�z�Qά��K�0r� �uLS�R�]��2�<k�@�XD����9��4���6�8Ġ�(��6�(KӅk��Z�:�Vu���E�>,�}u�V;������qsL�ǻ>�sgn�Ök��P��Y���]l ���Gc�mX�`��G��>8�j�UQ�PaL#w��}Ky�	�l-Ǧ�Y<t���ѥ� pg��I�b���܋�3���q��D���#L��P���H���Ɠ����_"���[���}�cO��}�(���F�.���2m8TH�3��PŐo�V,�*�9j�d��sX�r���G�uu��'ѡn9��^6������*�=��� g�M�@��s�0X���m�"a���Hn��v4]��r���"R���{�ϲ{�v�v��2���f�����k����N��m�} K���e�������9IM�K�(��rA)�����j�߉�[y��M��u��y���b��sД|G�E����G]�I�I�9
���v_�nT3�$�Y���%\͞��L�����.5��[igSrS3 ��Բbby[�|c��{U�<? �'6cz:q�w�I��i�h�?��[9CH;bm�>x肃e{7��S�y��+����ݖU�fy&J�B�I=~��
t���-�3�`�v$��Yq۲x��oT����d}7�b�Hb��ss��ڟv�]�ۙR��DG��@�{ ��ΘY�f[�����>ɖhTm(U�Od8\E�7���7�]x�$n�)��#<���{�&/{4���@���z|�֑,��j����_W0��sm����?H�9�nR����55����R)!j��"����J��cЌ���R%�'��?A�6�����X0F96ʧ��H0�T�k��4|tMԚ�ߋ�5��bZ8�J�I+�|[,3���}G22ӄT��?H�V+�Hg]C|�U�Ș0�n�s�����G@��\B~�a�㳖��uC=	ө����L.��@��&}y��&bB�K�UT�G*�SBޑ <��t�u�t����$�V�k�!вГ5a� +���@�}9�J
ϖ��'>A!�4H	�w�){��7V�15c�?���C�W��
����ۤ��+˧��C��U�����:gePd��0KGM�?�/�:��������(|�$�!�����䅲��
7֥4��B���=�ohs�́dω��9�,��/�}x��K);��o�[ᐤ��˷��P�ATFc8��=�t�}��¾�f�um�1��&�OJ�6���kQj�|\�,�]y���K���ȅm(2i%K�QE���b%���W*��w�a�`��|2��9��ĚzI/� 铻���s�}�^�P	Sv�,��9EHG�>��������x�g�u+`8��c���N&�+����^� j�	m�Î
��\:�ǉC�z^ZH}��������z	��'��� u�6d.2M�!�ϫ�?��~{B"=D�ͦ-Ǧ�i�
��ث �t�P�&h;
S��a�ZgREʺ\�n�b4����Tq ��u���w����'o,KM�BAS�(�5��l��|�A�o��J�� �I�<~3�h�O��S�J��|�?��/�L�E*ar��Jpc1�OORo������S�Z0��K�߮c�%u�*!�Bԫ��j�u��fP����`H��|������2�\�Gז3�va��h2��n����ȆF2z;�gq�o|�N�6~��0�]`�6Y�b�6
�e,�V��U����=��;p�j:��\��b\}6�D��/�b4H� �IeR�jO�J?"݊��.âĪ#���B���L��5�*Y�_�
��K1��Tx�>?0���~���6�*$�c`xk_�%G-N^����u��֦�1�V�l'������q�H����h�^z��G���H���?S��Ia�g���J�u$�ݥy�d+/�����E����k�y�Q^���6�e�� C�����=����=�;)��!X��,�K��KV).ݱ��.��V�~E�$�1��dN� ���[,�,lx薟�7���}�X#i�5���ƎQ��eG�xl�"@��;��˄���JQ�"v1Ӗ��q��8öjțk�q�R���� .^�+�)�R��i�$�� �l7Ϫ~l��҃J��~�y�qj9�Fy�tSZtW�'���E�Z�z/t�%' ��>�}��u�����*�𘑷dIё��I��4)bv/7�.1��n�9F,d�&Y��W8 Op���{ےܤ��빹F�Ә�J3,���3��m�R��Sb}�:��L�Ɂ
����nQ�^���NrY�J*�;�*^�9y��3O{o �"��:5<�OK7�و����'ֻ���yZ�þ���$���	�K��H�V��0xLs"w��e�(�ڷ�]Ƙ�t��Lg�B�T�G�)�͊#���[el�H��N��"@c�@8*�r��]6[�,�K/W4!�?�ӆ�	�m3�4�Đ��\�W8�Q�<+�F�R�*�a��dRvP��~����Z��gp�NL	TѹQ�.�7+D����uܻ磊Iw`�� ǉ%�ǈ0�{���/�Z�ُ�o������^�ts����x/`�(#j&�zmGPe��d���&� m(f��@�P��%K� ����4l,j��8���O�r֊-��}�-G.��
�re�/�r"=��il�*�}��:8b���u��	7��7DT_ѧ���⫋?���	��g��/�"�O�{�&�<j}��n��Ѡ�Ҙ��`\|A�д>�G��E��L�4M� YOS�4�0�q�=�g�d��ꇀu�T�+[������1���hx�/�����kA]��wړ`�@�u�e�1��-mO:�T�;s�����6[b�
�|�`jn��&0�6�o������� q���tʖ\�2�{'q(�m��(٭�wS�R��3v;�`Gh7){��d!���*�uHY��8���� ������4:���w#;��L��u�$��3�0ѐ3ԃ��)-�bC���`G��T��J���Ί��M��a����)�@��P��ږx�j��zf !x�[�$�x���7c@�K�����M��_W�� 7u�Sʎc�?J���i�\[,,���GF�%�G���I4��1,Ѹ�	�c��t�+I�Xn�1��8���.�xqicS��`{z=����h�gd
���\�j���Ú�o�� �n�Hl�c�l0�yr���,�6��(�	�s�0�����M�h�^G������T@�Q�}U��<2��i�Ё�=s�����"���J�d�(��R�$])T�'G�ӎ�+ē�L~��n	"iZ�v6�^�}D:A� ��G�5�տD�񪉢��Ƥ�ܚ�����r��3��?����rDM�,̧x2�?�%g�_ ��Y|ؘ�
���~���E�<����lF΍ -�5 R��h���G�т�C_�v7MK�Y�Qn�wx|[�i)�ٰ��~+�C�fC�6ĵ�"����a4g:�{�k�B#��S"�]0ƕ,h�[�'�{�?1:.�π��w���Лu��c�����	�	����?SS6wt�kÄ��SG��v����� AdW�䮱�W�Vv�EeD6��C�V�^��Zn$0�*sc��Q��%Cԝ��;��h?��ܚCρT����ZmAh�@�nYQed�"2���N�����c���g��:�c�ǈY^�	��N\m�\�^�3B��<����lx�V�������\�[ -����ԇ�=�6C3;4S.O�u]^���-THc���1�rٰ�W�%1&��!6�?R��� ��t�t?qW��ܘ[���q/�idb�E����i�#ޒ&+{#�U�􎘶ƀ0�»ل�Lٌ}���0���$l~z�9eTuv�9v�c[�5��M����(���"����*w�
F�(�sdqnЇ�:}V��<��nJc�����@6$� �rxV�-lȳ6��`^��W�Q.����q�P���Y�UM3+��1�b�Il2���b�-���c��jR�`��K�4Ya���N��x���saM��4�w���5�R�l!ݱ���3�c��l�r�E]=
#�K�su>!Ġ�����ϴsx	��\���)Eg����"�J��q�AF�{/���5_M�;d#Z)c���p��g�~������`�oէ���;�$Ż^4K�������� �W#"�E6r��� |�S
�!tzm6�Jh��K��6��,0�2C�[`�q.Yq���:�+g�Qc��t3�J����𙌸�����B���x�]������ڹ��MB��Һ�l�TE9��D��j2 ��G��޶R�2{S�
`��ׄ()l7�r�=���z팷(�j ��� fW�`^�6��&�!�%�[��R���!��9��_F����k���J+0� %�PV� ��J1W�N%H��=d�nirޙW|�2�mk��3F/1�յ:d��	�650��sڎ�/����o�˸.���~`�l��}VZ��8c��%?Z�h �N�Җ��t\����ށ:rG*��#+ϓ����O59�LO�h�2w�Mv-�^�z��^s����1� +Ԗ@�̈``Q��c�C�Pi��	xF�B:�r�=Q�;W8��wK��jDͯ7)�I}�.UEM�ľh���~w�.��!A[@nI$#M_��dE<N�e�٬l���x��r X�L��q����b�s��LU����R�rS���9ׯdʫK�����
5q�N���4�q�c�J*ѭ�
�a˭�F�:߷���F{���Bp�9�܁E�y�qg��wN['�tz8˃קd�8�![��r���Ƴ-l�n9�c���#gM���⨯�"(���^���'�'����v�鸆3��ы r�C��)�M��6j90�&V٨�vf�1�4���-��H��r�gtcj{�a���{v�}�OaQ5�����Qm,��/z7I<�!6�T"�Ҧ�c�/;��N��P�|�P�K��Y���ZR���O6��*�%��>�} Qf>ղ?�Ő���fH��q9�j��k��Aی�J����]�HX�R>䯓���w��z���'�H?�N��f
�6�g�W�D�޳T�%4@�u���]a���C>;�S�����ʔ0�+TR;��"b$�O�|AP���$��^�`��_�q�6�	�!.�?��U��ao�ݛ>�D�d�0�B�lȜ!Ł��4�e濏W�_�ٳ�jO2�3V�Ikʁ�0�A	��Y�V�!y��F��Q����C��ӓ���H�{T�-�c�Eހ�����R(�^�a]���-�|0���"�u�\�.�W�����l�*N�� �gC���}�߰�T��q�\XK�X�9�K�6ϗ�l��_ ���⌉��-_j�'k(ҏtv6������{ҭu;��8�~2���oڼkƿYv�Y�x�KQf�/�Fʜ����Բ��I�7� �=��"?�]_uǘ�5����~�!.���F�/�)�0��#rG�K.��% Bc�>){���2�Y�S����=�}-��]�t
�gLO�rrQ[� !�=����5^zc�o���H��}�(�4��qMt�e��c裵�(\�D�s����/W^6�&s�} ��>�9#��(Ph�w��S� <�|)��A\a�RL>�Wg�-Djg�؅v��3a���NA|<�4�)��+��pS<&H*����P7�^A���,~��4E�Ai��[�[�l�bf�W�"Oc�麘�g�pJ[����3�hɟ�>��pq�P��A\C[������n���7�U٪,5�B�`�7���\�E�e�ݑ��_�{n��Oeg�{��&/�dI,R����LQ>��T�`� ���pk>^�?������:ɗ�	Z�c�8ݚ(���s����2�)F�^+��CN�uE�첚�+z5޽Q�
R0	�'`^�W�X����/�XZ>ݍ�Gi(NvZ�!&*�ؔ�������E��Q���L��U*V��2M��wyu�ݽ,�_ R�<��o��ad�0�x��;���B!1]���UQ�a�]�W���㲕Oc��m u�$�� ,�E�K�x�Vf�%hP`�.��ުݪ�S����ű,�l���i�Z4',����8��1(y�}S�A�Me�I,���~��������[�@�^����1���]�5=��r��	�ܳ6Sgi���4����>�;��FN��	�S�M��������<����&,�3��ӌ�+H�	T�{RLֺ����@1Muj��q����oxux̐C�j��\��hk���7����/7*gA��t���YV�@)���S���"0��b>��=�����Hz�}��)�p̏�?Q�f�(����6��Yg7�dz`��'0[|	%��`_���&JP�)����y�T����m�Bhۏ��1�SIY�x��n(��=K��1�*�����J�Bz���.���C�ΰ��p�� ��-��$Eu)�5�l����UE�I�n�4�~��6�px�Q�y�c��de�-H�֍�eC�k[2t�8R�""q�"1���̈́6'�}+u�߽�6\8s���4�g"(�z�>����G���0N��U^N�u���̌e���-ͷ�p��@h����1��#��&���Z�6�[#�Mm��+q��/':?�_�e%�.O}T�=��v"���3'��9_B�/"��\���Xt喜��:�#����_��=��o��~��A��{T��}�&��Ս�X�c����so\�|ϡ�.W���-sW���b@eݹu��Ҙ*��d+�&B�	���p�����DQ#����dZm�[�_��z$9K�Q��ëX�9'� Y��^p�D^,���e��m>\�t ך&�H@M�w���x9����E�J��a��Ei����=ɴ����hi�9���:���h�'$iB"�"���!�D���k���t��;��'��?lQ�����
,�:!+2��O8�rPE��mǸɯ�W�Ba���l�Y���g��)mg��Ƥl����dFZ��
�� ,��D ��BiL����� ��<�޺Q�:���މ&�C;�k�H�I��o���^��@�k��r��e��;�B�8�Fg\+a0�)�zO)�� J���y� z�?��'���*��Գ�>�3/ə:���'�u�Q��j@)�(�h�!� $�Oc����mNL������_�Q��HI�����[ Qo,���]��4���kr(�H�N����'����,������FЎ���%d
6�����Р��������b�׈1�y6N���;�T�b�F}N�.į8����w^&g�	=��M���s˦?�e����b�Jf�B�p�����f������/=�w��7���'K.K`�R��3�B��斫jMw�Btg�*����O���Š� 0�O�2/�H_d�+{��u�
,.���h��ݩ�{�W��+����r��bk��((��9�:6�r��:��u��H�GB�t���$�sYP�V�8�|���K'.�ƴXU]Z�l��	�EM(���KGj��pG�Y���ٟ.����W5�6Gw�`��j{�</�5�Y�YH�C�R��7�q&ݔQ��}R|�k�a2n�����\q�&K�aDb�]���Ql��U��磥�N�W`B	\2s@�ш�s����l�M�x�� ���J�sH��J�X�FωG��h�*\�#��|���/��[�
�S$�mt�R@��8ޛ�� �����c8��fʷ;hg�8]!�Pyņ �ĘI�ι�k�<��E	���jd�A�P0tJ�`����$}�̮�fH��π��t9-i�|������Ֆf���R+�؊i��qa��St�! y�g"�� �hCB��l=�� ��E�L�xUK�Ϟ��­�ѿ��~逶zGǏ8>�A��m�0EC�YQ?*$������]�E�S?�~��X��X+	��a��p3;�m�.AU�E��5�)���(hrW[�~��c7���3f��$��r�?��F������tF(sRXr덶���s�Hq@2��J�Z�B5��z�R���7����u +�E��F���	�(��)O�/�a#���0��[E��B}�t�,�"E)�Gά��ޤ�#!J��&��mU]�ph4��z`"b�nNW�[5|\PV��$>����ŏ\^2͡�1�˭��c�ȴ�VX��j��׳�CA�x��r�l2#N��l�L�S��.~�"{1�̉VR$ϏW�`��lT���ÓO�x$Q���F���
�B���$C�\ؾX���5A��y�sGv� ��:��t5�>�A�|����.^�4���/�\.�wˬTe��Rn��v7��Q�[�PL���yD�g�@����Z�i	y��3��/�GT˶4L#���yXr�X�CG��"�i^d%�|�����K� 	�l�'�=�'�l��e�����w��M4EǙ�@f���Ƹ�mY���@>&���YG���W����|��)�
7�U�%E�@6G� vme�Pm�(5��+i��g�q�p�źn5dz'ԬyiJv�#�
c�dv�E�c�G�Qp�\����c���T������n�K�w���lێw����5������X�E/�'3�P�=7��NPm��J�����ՋB�7o�j?8ڎ������tV��#,��i���>��b�1��2�j���$~���E0���5��:�
*��i�8���*@��!�R�ⲓ��s�#}�ك���+aD�6���8|��R� �B�W�����^G��% x�}/W��_=}*�	m�b�6h�v �7RUQl�8���y)��m�ܑZj�o�G����`{-\gZ �K���B�T�N�a���xS~N��C����?��|���l�2&�6TBK��� 6����MvkT�Y�I��Z Vu�ꤾ�%���Yfgu�Uѻ{.Eu�Bû8�h�p���cg@uv�g����:�8�f�_W���R ����K�I\\�_���8~u�y�#ɼ��q7.��x'A�����V-�:K��UE�H�ɕ�Q�D��b6�ՠT��N��^�Á]���XD�6!t�x�!	���[���kK����-F[�h��}r¤����'�BP��2�(���_��Y8(�v�:=����ʠ=�����l���0��[�V
�0\��� �8i�WE~�^$�թB_�d��tx"����7V*�u�|�Nkar��ĳc@O�5oQ���{ڸ�>�b>uyEvE�=9	O3�u��e_���7�6���3u%�.1k�ef�{�+�
��[8
SB�,��+XJ�����F����Z��p��{o��bn�~{3l�8hud��tZd�1x��eϢۄ�j�>+H�|*�#Ґ�
ԏ�o�(��U��3��_|C��5���S%U��O]v (D6�i��p��α����ºz�u����}T���u��;Flt�^��ԛno��%�d��@>U% �HT�[�	P���KD Z�t,�xw|��A0��X��ROl���R6X+M�����'y(�HJ p'��4�bP=\t�5 �J[�Jdgڍ���fn�ʸ�2"qk�>����0A��=M��[�m!ĵ�L!��Q1a� ��bz��=��I�Huʜp�����GrkW�-.(�$�y�,��7Õ�<�1lGz���Q�$���q_~Ʋ͠qK�+�c����T[���lj�c��=̫�~��-��!{LbF��v�W8�}n���I���-ES����<P�{_�=G\��J!�n`Q��1�Eu��
�}K"�8��'��3ڐ��uc�΍\�S�[cU�	�����R�WW����p*sp��IX�ܤ}�X�C�6�����_�b�_�'�L��-f7�A~>@���Dӯh5e�/Vߌ�zp�Ҭ��S�YH�F7�=Z]��`�5��_"���O�������~`}�����AKk��2z��y7������3����(�E`�L�]��`	��1<(E���N3v$uK�,���8���>�7�Q��Ǻ��t��g��=<���Z��fI̊Z� R�>�|J#GQ����� ����v��!v��7'ͳ�T3���fه�ًo��^���>��e�lp�Á4������@,}"o�ͩ5���W�u��B���"Zc�D�t�ܻ����-�mv�e`D��)�ڂ{���U%v�=�?�練�	?*V�v���?ې4��b�n*�Ϛn>�NTtx�R
"�g�	*Y�{�4����z�JJˇ�,q�R���T�c�5��DR��%>�ͺ.�ݖ��5(��%E6A���Q� ���Q�X���-t��Gʔ��o45~�����D���_�*jޤjP�U'gr>
����܏.4: a�k�ޞ��<�iߛ"ܢ㲭�֬Z�g��L�:���^aX��S�hu�2�����kG��*���qL�F���~��О���;�VIr��M�"�X�hݢlڏ
�X���Z
��Y��Q\1�X���M�o�j-���`|6z����;���h_�S��3:���`�ޅ9��㼲��ǽ7|�p��s=x�Y�	p	��J�;�'Ǳ�Ԡݩ&~ۿ��M���x=׵fz����-q��x��#�\�J$����9���ԷY�[L�'(;WO�'e��dXsU��Kg����o*�W�� �E׳b?��e�:�;p��Z&�͓��Z�g�b�H(���Z�!(����L{���fK܋�`��4ƈ�f@�1`F���"\`<K��8�b/i~Wd�g�R�'�w"��/�6Sm���V��t�7�+`nL�7��8�m[��F�������}~]�< ��Eg?rB����x�$n8�Q������YA�i-T�{֠��Z���4%��Ayg
�l����qd]��`�?E�+�Hw�#��7>	�x��a�g�ݮ�z���'n�΍�rq��F1���ΡC|����!��P��7s�lT��
x���py�M�ad'�f��5�(��i�?�,G�S���K��[���>�i.�w�l
����]�=���-:��q��`�6�k��j��E�<'ۅM<,��yMb��F-iAL�`����R��f�Ƥ��J�2�@��)�������u,�U�P�au�[w�����m4�Lplj_���H}Ҏ��w�b��Y��e���Q��yJ�V���o�пɌ�$H���nZ�'��=�x�q��J� ��ux��o4�p6�L��+�<�}����Xټ�m�ϛ"J�R���8�Jm!t��-�}�6]��$�t�r��/Ż�r�Cۥ��j���ilgM�w1<�ns?5=��me,T�#E$������S�ł�I���APf�j7����h ��"�@�����
���|��H�Hj�L���_��lNM�b=��"�X��8sNy�����y�=���#�������Q6���7����LG�hc߲Oi�(��>�އll��sJ��T!YӉ]�E�<d�d�+�˂�ҐE���tDA��`@/�l�w�r�ĉ��1%גM�oI&l��g��(gQ�^�����H}����s"�� @�Av+�{@ʗa*[��
�=d�8���8�N43@�Xj����������^�3��o��%=Zwʥ��a��E�Zrh3��R^���\__ ��_��gR�k�d�}���T���i����I2�Z�
pF0��`m�Y_�'�TH�[��"���"F��F����|��qܹ���<����M�`�����|�Cʼr*�~�+J�-c�w���Uk6b2���]7�����T'�����;����OkmQ�D�:�s�� �i[������]x����6=��A��C�jr�N� ]ҽ��6���3vfj�`���;�y'�8��<�X�6�{;R�E44�晄��0gM�����,'�H պj� ]pA?�
*�ti>������X���P�Q�=E��"�H��w)h6�	���?���I; [BN�='�kYVh�ׯa�j�2�P�Ȏ��?K+��8��.s5��M�GǑJgc���U&F:V��Qj#b���W�́"+���W���>�����M�r��/ � M��B!J�]!e���D�*Rن��C�IB��["��3�vGW��s�t0(��b�5�\��7�4�B�0�ܤr�u��G�(i!ۺ�gT<W�w�-m��J'BZqO��nAJ�{�"�܎K�vP>C�d��������MdOEj�'�>����,����aEY�W��1��yd(�0��u��;^A�U�y�$�d��] ��jvY��T��i���B=ڦ&O 6��VeZ�f$t}�V�Y��.5g1����1oN#���i�(���������W����Ѹ��uH�2����3g翐=����+q��k��?��3�<zw��7=�/�.ʫ����<:AEnwn�nXnl=Dn��ˮ�<p�z��灱�@�GE���ns������Է��m���_����},�V�?�����g�0��M���`:�~U��' 7�o��d?)��� �K@6��z��$�.�W���z�j�U������@�%�	����(