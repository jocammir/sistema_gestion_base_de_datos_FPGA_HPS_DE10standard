��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0���C	�i��E��$��Ȯ�_�� o�	��,�}o_l�/5ո���-��Ff�16��6z��ԫ�{�C�"Q���h���2�H���������8����� GƯ�CSo� y�X����o�)�|�)������<.>3 ��(�v�wnM#3B[��>��^6V�۞�B��>�p�D(�����y�|���x����m�F���m�%c�d�o"�˫�@][_���~z#�N\g��!'������0x*hk��,	��{�x�/��*0�t�ߐ"A֜.>?n�_T����bC�U��|r��V`��0M�ޤ����������ռ3^q�RE�z#����#<˟��Kpn��b�8i�	�Y�sA�2�*č���D����,�9S�yN0^�T�Y���{�roT��tǋ�Δ_/��xkM�c���W�8k
L#[��l�|�T��p���g��u�R��Y�j�`�,�m�f]��-˗⍖n�^���z�lD����1�V��c��Ԇc I|k`�Ub�Ǯ�]zƱ�c6���Ё��N�6��?�y�����B���};��|�s�s�}PCQ"i��Wi�D�^����Pe/�0'or��S�Al�-�����>�K,��^��GP�`h8��T���*�?܍>�Ozϐ	�e�=8�<�W{�@n#� D��7���ö�媧�u�J��'z7����-1}�����v#��5�wS�S9��&�w���l�C,��b����с���@<�o�}�$	N�N��>����Ĩ:X�;�]9�54$��GK�(��b�a)=�$��˷�ڲ�n�0�K.���a"d�d> A�E��E]{�ֶ4g������|b�X��#F9JA��O6��FY���  1�{�j��G�W��q~*G�� �ٛ�n9&�ְS���l�����尴y����n�jh�o'ȪL�/� ��3����9&��JfB�#��o	���-��x���|Z+yI�Z�hE�|��HqH1)?ĽSþA�X�7f���y�n�s����� ����R�R={�Ϡ�
�݈d(cbJEM~J�Y�
m�zq���g�������X����.UJ~��>���˯�,�{�9��wЬAy6�K�1+��\��2�7˂!S���ȯ��kz�EngnGI��8�Ts�Y��r�_�������>|Ip̸D��k2?���?�"L@Om�xq/�Vgn�K�G%un�Q�n�7h&W�,4V�۰$���ʣ�:.�{ ��@�l(�������>�#Xm�2�\ �N�
���f�qɱS��.j���f���d����*��d˽:�:�^a��Í��V�M_��v��:(wd
0u��^�\A@���M�w)0��qIZ��NȂ� -
<�@*e�Ƀ�0��Ża��#l����̒�����A��*7�#c�AWU]Y��������7�J���V  L}��V�b�7�A�W�oR�/��#�m�h�kxH�0f]��\\|�L�(��_4�)n5=�a.�x%fyVab9�V�/�l�������a�Ǘ���Ϸ$��9ځH�-��w���&@�E$5��u1x�`k����Ҽ��
��QƩ��Nw�ғ-�0�@J,��C�����.����+)�����9����4�@��;Ïp�o��Y�(���kLv�`#�7;��&���/�U!��Gw�z�W��Y#cؓ�_k��&��UTR�%3ۀ����(.^�X�
�:���͋�@���.�5����_��Kc���M�ܵ� l�C�pƁÕ2� ε�����;X����uM}��T��I�T'�*β,j'�h����;L�w�e؜M2�R�.�Ju>�%��մ/��k�����kY<�r"����왫��G�mU�bh������rp�hJ���G��%݇�{��qV|�%8}�P��w�i&�Ac|D'�l�(W�Y�����%9������4w���u)��+�	�+����6O�2B�Bw��=��?�B���UNH3ZKna���r���q�m)�q_��x&_��$�6[�
#3�2+��;
��4�jnj:�-�1��*� ��V�ƻ�^��B����d�y�E����7#H�E�/�+���q3%�_ͽ��Qx��OL�*la����|q	�u�힛
�`^���v��»�����X��䨷��J���d:ƶ���4N %ĥ��A�xz��T_�a��'�*bm���^��(���&�g� U8�k��/E�/X@~X`����3J�Vy����Z���
��t��o��X�{�P��g_�Fj6�[$�{����5	qV5��\4�QM����z^��:3XV�9/�U�O~�)W��rf�T��&�m���K�/>!
kg}b�WN�� ^���)�,�(���Eg�P)�c��x�b��R
�׭�ώ�.'�E���%�^0:-7<���*{��P2���N� �9qe4ղ��h5e
m�����??a(��)0 R��ީ�)Q�:�hx�m3
f(���5�|&�Db�yE������-�>�0Tp���jb�O�D�ꝁE�ξe�K�vB����M�T��y��j�3�!���4��Q������=%b'"�F�3 c�h����@r)DWZ�A��p eBOE<�x*�$�5׬^J��T���o�;7��'�M�"k��Y�̛��t�D,%N �9�2Ԫ�'��#��!�f+�&ϼ�"KekDHJ� (Cw�̋��<M��Ҟ�Sv$˻�)>\^.�Py�l����Z}Z5�b�x>��r4�/Dˉʔ�ty���_:ϭYѸ�]fQb�l���v#��f��Ta<�+-&�Z�d|e�\�=fc�Ú���Cse��5��(�s.�{\s���,1��=�{�L�@�۵NɅC�D9a�9��d0.�9���Y���O4���8y�~Ҏ�0�+CIK�� ��).�w�3�䈊�8}��V��"��u$f����oږ=yL�2�=�w�h�n��hV(7 ]9r�d�z�i�?�{]N��i}E/�t�C4�E��g��J�}ٶ��I�cY3r�t)[�_�U6 4Hby�2�w�\�ł:��df�8帻o��e�3�<[sjr��8u�e��P]@�l��Mm+��0��ȿ�ƭ��5;Oq��r���I+�]����r'Js�zI�Qɐ/�H�$S���]F�-P�Y�5�eT����ﴷ�2�����먥B�6Eq'm�t3`{o�f)����#�YH�������EO�Y�T���Oj*b5-ן>������Һ�3}�S�����&�%]��u�k�����=Iݘ�F;�v	��i<�y��V���!��>DN5�cݚ[�b��٠	�o��1;��[#�Z�L.����=ἤ�*��b*uL��T5�bkԟ���ԇ���.�Z�gj�~��tG��2Ĕ#�y��S��.�s�K6���ޓP���F �D�hf�F�̑�vÛS��� }�=������|!��0��H.u�T���Rf�K$��zF���9Y�n$���:����)�G��0g�z'#ZgGg�qv�	���ߓ�tT�D�. �3Y���z�ᥰ����
 ��n����T����=	/�-h{k=�q��h�~���_ىy\e|�1�enL0�9o��OQ����xezJJ�8_��}���P_\�W7�f�ȧi�B��G�A� ���ݒK3��=�g��f�5��v)'���T�I�
�K?!�4����Gt�͔D����<�7T��}l3$�s�	����:���ݥ�_�{JT �f����f���(��V����5�u�S�c@����U��/54<4f���a�㭥c� �z��}tKQB�Zx<^�>oٺ5mk��/P%-�9u�J���$��'�Fgܕn���1siUճvS#t|.^���¢�X*�u�
�9Kh��_K� h��D�ǃ~�MKU����D����w<�vr+�k�3$oxû��G'���p��q�s�Z��i]��d���랇P:���G�b7�\�O��܉
�i/p�6;��v���r��Ì9O;�ǔ}���p��\m��<�:,�+}�Z,�N �xd.�p#<�����T۵���*�B3�Lݶ�0�~��J&N��P�+ƹ%#L���>�!�x~E�Jǎ n��d��y�$��Qi:v��*;�S�1�%�m�8!��Ń�{�G�af�2���w�����&"�l��H�4�e�ơM\��.Nq��h[w��-�X��ڴsc_�^��sdsE�i��`�T���]J���6k��N8�`���jY��	T	P��՟j_4���T6�x&:sIzQ-$ҧ�=�i���B̎���]�F�ddgj�Om�[G��l�ut�q,p�PMVG�G��eD�Uzq(R�L��m#��'o1S�h,���g� GKUM�07�c�c9nf����`�Ï;d��������9�����I�7�V�䰀x�V�efB�j�c�RWۃ�lk	�8�'/��]]��K��D[��_�Fx���1�n���p�௠��������R����u��W{�� �)��;S��fI����[�l�5r��C��uK8j/�m��;�O��]��%Ѥ�Α��8�� ��s�VLƢ$V�1{�#xOL
�O�����3 ���*J��%���lo�<�}MZ@th��|�����5�P��g3�"��u�Z��lΛ�����yQ����76�1�h[J���髢����:-��.��M5�w��G�<��C#BԿ�۽��4�l�6�"�ڻ&����Pn�n�T�0��.���M�o�
U��+e� �oC��mlu�IF34�L|']��X-d;E_����Ǜ�����	��=�+%��+)�_������o�W�Fk+��A���$�)����Y�4�b�Op���q3x�a.ꀺijp�j�RX���b����[��s�1���>c]zŽ�aMh�q�|��Z�_�cY2����_̻�����bj�����=`~m!󓔜��l�)�<*�����w�N��2+�$�[l�G����U�c�"�it�N�%�&(ö|L*A�P�iǢ~�#��C��q��P��a4<)7O̽z?�gP����O�!N5n�&b���r�z����-@��}�x���#�cʵef�5�����7㽩�#�"|����W��*lR�=��M�1[g�vu�d�O[PK���KuS�P'��" ��&/&�s�G�2�Q�G�����w(µ�<#{3ze B~��?��66Q[�V�>FT�0��_ձ�b��=%�ҵ�B���gMI2ɨ0f�%{3w�JֳKT�»㩅��k�|Ж)�mE��C��[��m�Ɗ@+��Ρ�w���ω��G�c�K&h2���w*=ÑC�Q'�B��b�?X+o����^�5��5b�yɬ�=��sEY P�~�5=rO׽3�}���3�xYڸ<�t�E�&���2TO�m<ц~���*�f[w�f�50�D� ��Uu�IMz?m8f��S�8�Q*�-h�+"K�"u\`�H�$�,Һ1	7�By����T��ߎ��9a�U�<��&�J�n��F�N,�WVUđ3o�_aA�y���&�<Az��n���%;+5�i��x��r����ڼt��-bD� N�L��c���
�tAoƝ�����#)����LW�@~��>]8����6~f�6���ĩ]���[?���"�P��X�]#Ҥ"&8�P�y�?�#�2?j@�줸����ʭ�S�"�����^��E^�`�� �#b�L��w>B�HU;�]�D�6>_�$��_�O�m����!R�۫5!f9(S�`�C���7�A�wVI�j�ɩ@�V���t����Ѩ�zU�2�F
��	��+]q�h� �&U�N�+v���sc��掭J�˗�o����1�v�� 	<ׅ�������S���#و����n��W��C,w�⑴,J����8w=
Y���to2��|ς���0Q�`�r�D_��'R�ң�������2 &�<}��ү�Cp���ls!�X�ݛKF M��f���/�(Z����\+�,��7o]V�ۼ�?u�敖�e<���F#��d��V������38{�rV��X�cE�w���nO"��5��W,�S�]�n�K2WS�oj�D�9��Z��z����f�$Y7O&�-󊪆��JP, ߥWz�=X��SF����u�u��rB���-yy�Ci�g���Aد��G|.
u깿V^|�q4���D�J�� �°$�ڝb#T�87��Bw�7:�A��[V�}k~�7�.ʀ)��J����͘Me� � -�ޢ�빤��|�Jm�S>9#/	���w���}?�� ��J�2s7Isx�#��L�Lu>�J��g�τv�xx��sv��1��D:�_��5��(��@�t|5�@��w�2�}L�|�i�U4"� ��v"lXO�*L$;�rd��,s����0��4}zɐ�z8�|���U'��9���/m��Pa3�,�R�ʯ�g���o"��i��H9�L
mjq�pВ6]}|U-���0���O�]Q3æ� ��bȻ/����g�� c ���aIݸ �_��l�}��,�9xPx��Оdj!�K�l.�.���Z6#Ҷ��G���n#�3k���!v�	��[��8�W�v�{Yߵ�C�Z�e��~j:z�R�i
ߗ(�����5�Ĝ� ��tf�U��J��!0�E���O��N�K�J�{�����]�v���j�"=뫂�P��:P�'���fw���UuN HX���Q�oX�҂���gI�'ܶ�L��D�n!��h�D��
���e1��]1����yʪ�0����g�_�%d�=�~�����߂���U�F7bk��Hk>s��n����O;:Ќ��Jr�'t'n��i��'����7y�)*�lN��ˉ���d ���� ����!Ъq��2���NB�;&���r`��βY8�=v��v����=���=����?�g_ �n�I���Ni||�rװ9(m��{��Z>O�;dH�t}����I��
y��X�݂e��
��G�ι00H�E׊N�L-��Ń`��X2l���0�b,���R��AH�#����:����D0�P��Pu7��J�P��ז���hCW���(Z��42�dӂ{�g-���>#y���W؆�� �J\��U9򖗺#�~�B@�����C|��De�8�I�����p�����_'d�C�tI4aU���:o�N�)@��z����9���??�y,�	����~d*�"e9��9(AbLK�5��<�:�a�/��*��j�vXGU��/�1m-A���������>�+N� æE��~,�-�6��鱷5⾌D�[Ϡ2���~b,Y�N4c������-ٚ���ȭ�2l��	��4�U�asۺ�u�C����Q��E��ˀ���;�_&�ɂ/T݇urG��ِ�\#�oT��qY�ԑ��t<����	tG������v�|��=���&���	dk�<�jՑ�d�׆"���Ժsl?OZ����B&�M!#s��0�3#�"�k�mیY��_M�-y!�Gq�{-���	��
[��u(t�
ntw�����VGn�d��+���ذ�_�.�f��ǻ�)p���h���q�6���>��+��P?2PPm��h"�E�J5�٨˲4B�a�0�3bT9 ��S��6�P(���pa[uOr.���q��a�@�j��q1�<PgȪ�'�����!5����D��-c��AxY�㜛V�xlf���q{�a����m���;�Y�W0�Iyw2���r{zd�Q뀏	�^���+�s�o	����w����e\$��%��M��������	ï�6AN�NyQ��^����šA��B8uI�Zej�.��kU �3�+�'3p��~s.% :V�B��������M>�����������(l����;�-�B)����O�c~3���R(�g��3Wh��ۥJl!e�s���7��ǣ���Tl��Ja�aFˠ5���9&��<�21P�*p�a~"4ŀ��~N"EH��Y�y�.�!�r�.@dY��{���Gq�Fg�d�+#�z�7I���f9f=q[�_Ձ~��,$��%�#�5�<����b��j��ÇYE��!�{��;��rw��1�Q�S��ͧ�PȮn�<x�����MUE����C���̜`�;f���gqEy�u����@^��z��)��_v�l��VY�v��\.l1x�3׃A��2�����y]v6���cAN�Fl[d#�r2Ш ���8�9���UH��� �Z`�RN����Ա��:���p_�����w
�>Xm�2��[�
\ �P���|�����"�ˢ����7���1���,{ ����E��'�9cc�=�t�N<b�	�����z'[K�dW-|�^z�c���Ny.��4OCh{���B�v�Dh�聺�V�����FZ��Ũ:�_�Q�H@�zOV�p�^.@S%D����P5w��+-�¥���Cc���-��^�B:���n��$��x:���� ��ۨ�Gj[����3�n�j�c��G���{�:�lcP��b[��eyl1�[��,,����/��͂��s�N����Xg0�%�tҩ�r��m���'�|��jYRd�ĩ`O�0������C�.��W��*w���i��Hwr䍵����G��K���'�7��[eR]zֺCݫ�\�p[�Pe�stL/�{EpU���ṩ���P;��K�7��zW��ԒwNh���m,:�c���a�8/L��M�y����c�e�b?ww�Q�m^�O<����m[z�I�Щ�>wa��22Pm�C�x�{�^�.x���5�� ��(�~��47�G1X�z�m�0�U��r9���"��c��s�M��F,�X�!�5m����ɥHHwE)ؾ��*�8�{KV��*+��v�S8u�} �˭G���m�?���N�"!|М�2�¬�;�d�q6Y�Ǻ��P��ޭ��[F=�.�N ˢ7#�"�k��/�l��6}Z���������dH����	"!���1��8�܇=�$B����r=���ǐ>*AQ#�-��e��"+ҳ��+�NnU�V&��$7Ot`L�q�6�n��3���v�bΔ��=��\�!T��PU?_�?�M�qh�:�c:� o�юիa��J��C��5�SB��w�hVW��?���_
�Ҟ�p�|�Cs��Lc������>la��$��:���J��?0fY���I��k\�=���O�CݻbkQ�=-�D�~�t� ��s�bp�1�m��zH��Ў�
`�'��E�{E6ňy�K}��ڃ_�@B�ie̞�Bnv��,F�F��<>i`��s�̹�O�N0��Y?ۡ�;���6�*YK��z�U�$�1+����̻@6݀��\������8��HB�= O6�Y�k���O;d�k�Ӆ��Q�r�]��*Xkfp�"κ��	�g#w��-t7��Y���g0K�[����p�mx�� �s���\��_3���q�=��6	2�D��M�ј Y �K��Кx���j�}y�_7��^5���B��Y�2f�WM��蟲�X��(��ѨO�#��J~��f���@�?�Q��b��e�wR'{ZQC��/��n��bt"�]�qœ��
6���j�*B��eZM35jA�?z�
�9(������nCO:�F�*F�C��*W����ߴ
�8})��xR�����,3��Oo���"�
�4�B�
~.�)nE/֋:Yj7�:Dm�VB��q�5:����ᛄ�򱑯��^��˯u�~�({}:�w#�_��3�a����܌����F/�:`s�$(�B�36�(H���;��Ih���N�[�2M�)����?��3FQy-�#nN�b��hB�|���z�ULP&t��l�	u�	�Y|T�w9:�.~{ٲ��jw����,y����$����<~��2?���pNp��
_Z�j)OV:�*�ue{���:��[Q8�a.�Y���2 �)�(�������#�='+1���R��)K�3�	{)�2'�˔�H^5��j�q��,�F��#i��e�e�j����g���E��	�0T�M�E��)�����	рS��Q�6p!5cm>(Q���N��n4@���.T���+�{�"]*��|l���l��.[}��f�����2[J�V�3��{|M�U�H������I�;��ZN�8�6kH�]��i�u	
���{�k��j�k$�i{�Ue��]1@�?���pS�н׋�}�drt��\V(w�P�%o�~���b��[A
�veE��N�wPZ�����`4-��
'1����#핯�*��H2T��J?�9���%��mxҊ��ܻ��)�x7$��TX,2x�x\&��A���|�ۭ�T�gG軹w� ;gE�MK�T��'UFvi�+$-KC'���6���� ��U�������G��O$�r ��z�~F���6�����Y:����K ����@��ej���ר>]>���� S���mG�{!�3�@Iܤ
��Y`��ar/_7e��o��n��C��q�J�P����9�Iޒ�x���:<̹F�9����N�����A�|~����!A��#��׈������P���@��@'������ri�b{6z��ʵL�ݸ��in« V3�v���e�&��1�̞�\�$+���j;�&Sd68��Zs��p��`����x��fO�E�t��	��K��;�o��H��o`iN&[�D �� �w�S�)����1�^� Jx&�3��Ş�t8y8S��ō����F�ܺ���
�hH���U�hU	������je��ў; K��)�wqa��^�m�8�T���H�wg� �Qɪ�
J�r U��\�ή�`��2Խ��F~��2�6�q�#N�����Sֹ����永4���?&t$ۅx��es�'@��KoC'��\����H�^��a�PNSix�dmh�Ӹ�*3"���R�P�.,đ��P�O�]5ۛ��Qar������8p��v��@��m�系wY����w�<\j��l��_�sǗZ8�9�A�B��vb��%z$��c�*�B|����*��o|I{N��7CC��ӆ/�i=iը�'��l���5�m����͊G���΅/�2�iڮ����D�;�|���W��ː��
��cƣ����<��*�I���G0��:C �c���;t�����r�yR��sR��m��?9�q���-�E���
"�ӂKALpROs���٠K�z'N~�r��|�)^Z�SKd���:zI�v�D?�"�s��rZ��o���6��o ���V�vn�v"~�����l}�ĆgF�:��K�8��mLRJh�ܓj+W!�b<Оe��M �oe�T���`�aRS4@�5����z]��j)5�B������> &��6�7�b#Mecx�h�0�h
ߴ�Ӏ 4��s>{�������RC�g;>�rK�>s،����Ά�·��6���z�/f9��"A�y�Y�j����ݳ��1ߎ�c��NN�K��L��)d�����8�TXÍ�Z͒�7��0k<qQ����Q�EC����f:N��*ܶj��f�V��JM#�%fK��ry�`B���2W�ɤ����D�Iy��(��yp �E�e�����l�v!ل�����1̓��X��
�ŢLD��z�D0��#u��B��H�mS�*�q�0N	���x��ۉ�B�jh���L����T���]�98�#8T>�f$��p
�s/#m���/�=T���E[Ѭ�]��zo�%9��2���A��V�q�zކg�-2����W�M�tE��Q���o������9��Z��f�O��� �E�U��iJ�8�~m6�z��|E�N��5� %D���~���sP�K�K%��U�y�f�๰Ya��G��yR����03:{�ߏ��6�Ŕ9����5yR�nW �b���b`HOe��X�U�Ѱ�ق�ٹ��F�4�,�{*?	�]����C�§R�?��ا�,R�R�e2��ȠhK���9jM��V�9��j�>(��a8�~X��Sݶ��嫀��;[*CUa�8Sxͼ�2#Q��Q!(��ëo��#�t�r�k��q=�ll�x�'�
�z�����C|�U�Q��Ǜ�>��܊H�z���NK.����J�w�Z{<��`a����uuo�h�����+�����Z��t��7/�bp����?5����uc%��Zg~S&�]bz��CF� ݖO�Y"����H��D��q��U7�Y9�+\z��]C1g1�B,�.!}�����\��P��d!�)�z�����2s4+����1δ����`4��Q�ư���p�w?U���d�;�!t�a��Ɏdɭl�N�PrG�%0$�G���w89��?�l��$Q1~F��o�"�D�!�O���:�zR��r/yJDe��������
��z��t����CP�����N��bU-��f����5е����{���eG���?���ػ=��4[/����~�U��X��e�E3yjM"�5<-N����i1�/y%<?NRS-�@Fn�����!S�Q�2�ҧ ��$L)z7�{gr�x�;pˡ8�ų����)����Z�C��l@�E�Lf�
�}���ؗ5k�����u��F�i����ؼL-�>:�
���+���zd�!a����AǀN>���/�J�gvѶY���x��y%(]�w�k�i����!@��o����;aMS�ܜM�����|�F�L�����g�����f�NdW!A-t��H|�	�S�9^�>��Y��n�{���8�s�2ɛ6�p�b�'m?��IY��=?5���\���gc�v,ȹ���̵��F�W�a�M����0#8VgD�S���_!�ޠzH#�IV��5~���E���P9�M��r�M���r�0��]u�(W���]�e]5���P����
p?�b<��0�z|n��@�F�D!�c�&)Ҧ���eU��uN��nN�6�&�ᛊy9�v�<������0(s|a�}R<��SDB�нG����$�/ʓ�T�;�تף6="X�L�k2�rC��v�<��d���(�$��.�/���a|�\��I��� ^c���뗲�|�Լ�-�A��8�o�����]=�{Ax�%�:pH�=!�qQ߬.�ޱTdG���D��(�f>lO%��cxI9��L�	G�Vp��<g���4���x��W,xB����:~/����g���N�Kvz,��;u#��_`e!�눕,�k�F�NP=6*q:���?#�D�9�
�b1(����:�4��6��T+;]�UpC�~8_�hAG*��0�XᯮXٌ� ������ZSɆ�R��U������O�s�wG�;b(���z��o�+a�n:|ݣ$�g>�}��&E�;�\��I.�P[؁�8P�]���0��Y,�6�CPN�|.|��#��S��A�MR~ls�0񏨴r�L�-M��.+SG�i��k��o�	*s�
�7�[���[��aj:l�5R�m�p�y��fo�J���~��r�ɍ���*�Xz�<5��������F�ۘ��Ɗ�JNV�B\6�H�����yI����˜ճNx�ɽ��T V���Sص7�Ljϵ�ѝca�Y��ho2�:07]���ޢ�<��+�T7 �V��d���³\�Eoډ�V�Ԡ/����ka��\1��>�c۠�