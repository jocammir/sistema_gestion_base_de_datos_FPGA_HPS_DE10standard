��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�Bd���eE:��ce����D;����m߰�I�f���#��-�D��wbrGm	�)���h�R8�k��rj���[��u�
Ml@��#_!&'��mN�F�	A��G&�W�5���k##�L�
Q���]X�iV�b8G���O&1
��l� �TN�z;p�@	�z�u�vH_E>ƫ�s�����"�b\a�GYy,�#�����F�j��8�����,��J��>3�f��e�
��q�Vm˟$���ǚ\�:SSH7��2RZK����j0M�q�k�ȋ/��Hձ��okuND�8.m���`F\I{L8?�V;�4�]��"�s_6@�듐B�d#�*�.�G��n��J�b��r�E5���FG̺�+2C�'_*:��o�W�4�̂�v��NTq�zܧh���p�����~[��,E��o^I�j.��uJ�\%e/XI�]��	�q(4��+����6���#��S5d$DN1@�m�<m1+>����x����k2���3�!5�������5�IH���gZ�g�Z+��^�P�ڐ�K��Vl.�μ|`��P���; i=M���U�&v�
�r�]lt����K�P�%́���U�5,R	A����,F�}������'�a>C���V�h<������4�!u��Ə͜Bp'�k1vs������<#�Pz8(�Zv��� ��:҃nά����j�qBO����鉥5�����^ʖ�"�w}C�NfREm:7Ɉ��qܻ;�ў����`#���+Y��R���Ʌaӷ:LW���G�dc��TY՝�o��C�t�hMɄO�5!��?hci��B Z������#����{e��ء��o��ŉUx�x�&��o����l��.6}O���3}�r�I�9d��s��Y�˱Q�p��d�v�è�>�S�`q�4&��f���˾U�����j�T��d;#�?\�_��_�@+}[�웄銯�d���}�(6<�)*2�~�+�U!�4Յ�]4�)?~U����'r�2�,���N����$�Kk�h�f���(�ӵY��因��U���N�T��J����G �����K�w��~�����(���������Q(-Q������^j�ӆ�2��{dU�#4m;����6t����@��ݳ�L���d��M�
   V�u�ǷM� 9◩Q���	 <c���%�6Ǝ`��Ʊ;��P��ʦ�ORWh���3J�O�Uqcص�@8`;7驥q���A�6PK�TR��w�����{DX[�U�ѹ�˜kqz���t�l��a#��	?��QZ��|_e�uF����w��J���\g�T��=v%׷�X��*x5]2���M�S�Kq5w�,�Tc��B�9-ب�n)/a��Q{�-1	��N_E	�~Lkb�ӥ����K�d����T�	ʒ\��=���()��m� c�S���@��&lpGG*k�,)�ь_�*��U|l0��w�VE,��iL�eұPd`$=�����6+!ݘVdQV)�[�����	ca<���N��>�,�xPrKJ�;y߹6���$�px���#�=hxQ��"��Kn�$�F�D�
�AY�� ��_=.$T�B�T��m�4|Ū�%09�+w^�І�C}&�����Z�e�H�dX�K�H~��k�Vu��u�(E��<Z�܆��%�+��v'r*��i��[��=�|�E���\��v���6�\#B���a?+���6���/�V���I�.�� �#�j�̶7A������H��qqU��� .���Dro�о��@�N	lZ���W_��=����nS� M��;�sН�Ե��D�W�@����޻��F�9�?�Lk]u����Ip]I��������$�l�5n0��1bW�K)�j��(�:4Xf4���Q�5X���3Q>dN@�2f���k�t��uф�^�Wh���q5���q���[�
�q�g���6H]��h���G<�����ک?ULV�_9H��Q�!}�7nDi��5����@ s��]|�K�Yvcbz�4���R��r������{����ŧz�k���Ք�x:�^�&'l�#3R�v�$��w�A�݌Bz����<�]r,��VU�T�r&�c[�[��.〔��<;?H�u.vp��3Y=���Q[����b���_=���5<G\�O�7�:
�&���g��c
�?�C�;�w�Ѱr\A=�/#�d����V���~��"g��f��_#v�t�`G�Ui����OИ��x�l|�G΄yot���z�#h���g��t@�oh���DV��7X���. �����撳�6�%~�O���%�h��&���d�Ḙ]����q�^IV��8�Y�}+[h���H<�G՘�Xv��
:�H�#�a�l��hH� ��F���.ё�~�gW�Zm�$�	�p�mғ؃���nS쭰Ѯ%�ѥ�	-we��b���AҕQ�FC�j��v����EQ H��/x�^��2$��0�kb$��IÖ�����1�]N%l <Ɂk��Z��*B�sH�`�S��w"L�Dܦ2U[
drM(c��iz�]Gn����!�fwD�d�v��n�R7C���W�W�D�T���\w_y`���=�Ƽ~�jpEڍM�Y�I�����%ñs�s��dț�*D��(���V�SQZ��֪��a<�SV{��ꟷN��;޾.х��L'����iq�|��:.L�f'�BD穢Q{�d�hNӃ�,��$xPy"�a��N����PV������}�LR4�E�*����>�b�^ �$!��Q�߶+�#���0��֟J�O�	�����x���p���JN��*#r�����;+�v?���HL�<rݫ��r�Ґ˾iUx^��Ofb���|yl�K�+��Mhn5��z�q|���ZbPO�D�tvo������U��Ǜ�ln�蒖�������A(��*����zґ��T�3��H�1�f�_����48��d[@���ÄK�$
�A_ҙ=e-�Ǖ�y�@��-"b:T)�x�Dpz���z�����S���[bN�:a�q`U�����~�B�<��_X�Nr�%6�e�J�p4�#�e���G�U�+�w���M�ɬm5��f����ê�1�y��U��tE�pqS-�+"^/\=��)��R��An#�Wet��Q%�y7�$�G�x�)���� 4j6d�9���4��o g՚>��p��9�_�1Q�
u+L`�;�k<��42���{�EF>8����EZ�����iW��!����Qc�S�����G��S�Hk��G��rϕ���>�{g5�u������ֻ�(2��'����Շ�-���w�gT�.����L@;dB� �;$��"�}-���w��<Em��/#PeB.�jA`���`����}@ޟ���pT����Ѳ��=�R9/z�$$��x��?��m2�*�9zݑU�1�Of��k��z���
��*��|�lCf�V`�+����s~��~l�-��@z�t6�E<Y��_h�M(�F$$�j�'nq�An>�f����S|�I��f�X��V��	(��c�nT���X���ȕbtP[(dUz�r+�_������}�V�1 N�c�j���9��U���c$��zX�����������.��D�C=^��aD��R�P"���W���쓋w�ڥ8��X�H߈ ��;s���jh3��𣑈kl�)Ӧ��2�6�*1>�����R��7j�o��s������R�rg�}X.���x���pt��40T'��QOJq)*Z��e�S��W g�{k*�7fI�������ݵ�8���
YI��@@+��&�1ȕwtXO"���Ϟ���<m�u[��Wː�5JyJN:���i����+vuz���;�ه�0<#q 4S7����q�H[6�$_(5;���� hO����N)@� �;x�绛Wʾn\���P��ϛD�8 ���X�=�*���ŷQ��.٨�t�-�k�&p�H�bG����o��
�9cZ,)b5c�"�P�y�8�&X��[�n�LQ���0����'4���d�9w���]��tl�DqH��솏�";�
����3 m����} S�·X�!�OZ3�׺�
�lW��퓆��){�ѧMi11��g�0�vq�DWd�CPF��OC 'm�g�/�D	���c.�3��){+�7>ޗ��z�H�[Wy�|rcp��v�\�c��53X�䙄{1 pO	��'>t[A/+ ��_����,Of�
�q��-��`����
�g[�������I������`I��U]�6��IB��}C6,7�m�4kU�כI���t0��SwǦ�P�9i� �C���.	>4��a�_$�"OJ�H?#2�c3�J���B��)��9b� �cy��V�w���J'S#�ÿ�]�:W��}��:���ۜj�_��ǔ���tN�]��'�@q�&�o�;�ۨ���3���d���|�S��f	ݨ�q�L/,>�R��GT@�o��d�ͬ���L��q�5:�Nv�1�V!�x�%�! x3I�5���>f�0�K-�3��;�]�4$�Pt*��&�^>�fl}���3���6���������)���o,�{h(��:�K>�Z���Uwc)����Ȩ>��=Ǘ2S���/��x'�����Z���ݘ���}k�*��E�VIX��v��"�6�2�t)n����M�1Y�����ĳƫ.�}�	����y�u7��S,�/0Z�Ĕ_>.�7.��u�g�`�1���SݱmH���}xQE���ºbP+(���y�׃��o�-�Y�]��f�"���
��/���OH�6�:$�������ʝ�'�-QzǃM�89��:T��^b���Z�mڽ��K������f��o��(�A��)� ��{鵞���޹b�G���[��Cl��݃���iQq!��C��F�ߩ�1iI���G��.z����p[�nh�C���]n�5��c�H�D_�� �Δ��c��|�o��@�/M�˘X�=�Y�a����"h�x7|>��]����I�..�#��h��)?ŷ�'�y��ӿ{�jyd ����H����H�98����v�4�{���b���ݑ���-S���*R��'Q�"}2�T�sa��I��n�)�\vm�Օ�����,~��K/c�I1�t܋�¯����̠9�L��2��knF��K��z����"�N�� ��։�4$z,(bL�vo�v�D�{o��s�t�k2���NO������mY,%�^���W5�T�������[yI�Y��0LO�IB MV�O��wd��'���L�wx?���:Jȿѣd^�"�J?�$,�a��DI��@���!# Ԧ��a�T�J�#���.3� %-�V�݁M�5���X�-�@f�7� %��#L�.@a�D����X�^�^hqF�6�1"M:���`E�}��O����*~Ms���/ �iG�)׃�t-Be^�x2�@���]u�P�F��g vht�ΐa��r�z2;��������"��|��c�=x�T�� Q�����o@�,S7t'^w-�9�0�G�ꐎ�� w���;�	t��T�ߧ��]���x����jM��J9���[�Ώ�Ϲ~���W��y�YC��u�\\J� �u��=�3lՍ[���h�P\���)�8��F����&c�	�)\��ƺ�#��q��]rN�:y�w6L�yj���^Ƈ�RQ�x.�cB"�'��Ll��auL�9��@
_�B/{Я0��7}��S��SrO6�f��y pg`��&�����1j'�WҮ0G�{,\�����c�kՈ�j\F �ͧ���ϑjT!E����s�	��E�����mI$��i�r�¢�F	�Y���a0 <�8��ѹ.�{/Aʩ��-�	�4�2�4 Fa�|8��w������;^b��75�Q�E�Dxu`^ͽp�����i�b0�+�	)�}K���$,йhh��)���Ŵl؂d�l�d��<�h���r'�Wn�|��1�(��RH�v�X@�+6 +��ok���"Ys�cC�e_JS�� ���X
Dy�����n���8740�(�㌒�������㷂��e���8irྨGa ��^�<YJD#
�c蕲p�g�o��	�j�ޑdٳt՚菅�0��ҭ{��!yb�}u��yfJHhW�x��S�����7�ՙ�î_��GPB���?@�xj�.w<o�l[%�������F>��P��plI�q~�X�y��F�@�5�'�#�:>�vw�Z[
A/�njN=���vbc`c�撈��]�_;O���>d	�8�Y�8��@p�Pe��o��[̭I1J�j���fD9��^��S^���_׿�No�J�i!Z�;�¢o�lC[��q���# [T�\��8��9�:h��/]��c��{8عp(Sx�3V�eUR��s50�}�3�{_�q1�V��b�M��~�F�m���ݤ\V
@�)�빂��k�#o~��;�@�
�t��\�
ݩ��z�tc|��B6��$4%f0Φ�iBؓ���뱼"&��҂?��*g���?M�"�B��P6/"��k�yمP"Yq�@]d,#���ą��MJ�`�m�h�Nͪ-3��_�#n�禝��־��~��Ǚ�V=ߡ�}�7K���3�x,6�~0��k�Cȫ��������2'6�'b�u_�"�"=ԉ����E���H�H2��D0m���a��^�݉����8�V�!;/ǫ�$S�xh-A���䌁<�\�'��ŧ���U�'�ˈ����C��o�WS�ߥNv�����B#��n��W�5h�H7[qn�C��R~IV�O{5l�H�+�/�l���P��1���*j	B�a$0����W,vr����$PӦ"{j�� ��q���'ԍ	�Kc,O�ED �-P; ���L���+��5��:4V)�@�DXyP'8�)�)?҆�n���7�2�St)�c��`���[��(
�W�B�����T
�c�~�̓��Ɛ�;�B�mOd evs��X�X��P���#�����Jo��8<�"YD�J�$��zZ]?�dȼ%�����b���a��o�L-o���lMa��Z�4,/�xn�P�U	/nbvv���ݤ�F�ӻ��!t�v�s��j�e�L�H�:Np?ڻu��H���mS`Q��}�VV"�W2r>>�F�c��p�9�z�M{_J𯯶DDܣĒE��/���}�14�A�0�HZ�_9�;�����EZ�[�oUU��3�'}���̏I�^��j{%u�x��f9����b��6�y]�T�����;�R�p�	�� ���)����l����]�q�U�>�w�I�I���5.�F���VjM ؑ�X��>���_�]
h|>̫^��ڀ!}2�*�9��2H^V�wj��~��M7#��)���-��{�4~����U�l�]��#|�4)��k��7t��ɝ��vy����DjtO���U, A�c)�*�ޜ�'I��-����124�P7j_��}	Rv���i&�y�4���«�NoJ��,댮\�q�X�3�L��v1>��=3o�h;/Sy�=e�H��{߂��4cל��$�˺��fٯ#�j/�հ+0�c��i��Aҵ� ����_7-9	�"S+,a�I���Y��p�������^�ڧ�I���f;Zo�4�s!_��h?*P#*�#��Z�za��G��@b'�X�W�8�ҿ��<4=�i���V>g��?�1�d����!4@XM��}���X�d��XĠ�rc9�ܬ�K�b��i��˯Q����z�k��/��;�rݔp����0��T;���
�ހ���K�K�����L�������QZ�\��V��R���&���7��q�g�H1g�����4��N��:\f�jK���fN�98%[t�
����ZϷr���S��I��G�	�]@)�~I����s���!��pht����0�7�R&����]yZ0r��pK���L��a�����N���_P�r��%Q�ɸA! ��C���o��TT�c-e}0�Ԋ'd���;�? ����]*?5�h�� &>��B�4�IW�߈����H�$eg�0"ԁ�]����<��D��5�ڲ�W��s@�h�j��2FR*�ݕ�'&dm��5K�瀨bѭgK�j{$�8kg_�������nŌ�=ssK��
n�/�L���b����>�wyo��~����La��m�k�ŗvtG ��*���k�(�t�s;l�sBA�)d�|�<w����w�<(�����j5�4}V�̵�)����G�;�(6Z �rK!��Hp�OgL
#R��/��j��̯|���,0��J�[)Y�?F�ĢUN����j/�<>�4Kv44dH���du{W�$�D�b��?_:���LٶҒ99R*�p���?H�
߽^�'sh��&���:�l�Z(V��D�tcHƬ!�$�e�sJ���@��{�����̊;��hc�|:4��{�Ґ4���p���'���pu�E�%�-U֟t����E4ȑVA3{�9fQ!������
x�����f�9��#�~��fl�Ò��|Y��H��ċ�%c���ݺP\\��q>��n��OH�� ��1��h����(�Zlu{(Z����(��P��c{��ѱܪ�ӫ�F;�x*#S�XY0�4w+��O���	�p��
�w�J �=w7ibZk]d���^�j�6�^���!�i1WS��Ռ��%�[���OBj`�������ia�,{�*��G�Q'nD���R]�*���\���+�x"@0�.�_(��g�D�nў�Xeĺ�b��tT����|�97Gի�A���EE�=n�0\��8��+��(d����_��{N��m`X��`��軽*B\����z����E�輘�Ü��ݵ�>:�t�G�!k��ݮ˭��6�J���16JF���CY7?�V��V�<P��� >�Q��#���Kgc�v��,;���c�Ob���|`>g�̆#XC����ak��`����AG�2�!��w�d]���?���2pњr�X�:N�sQ;Gx�������Y�� �)ډ��ƕ��x�א�Vjw���!�f(��\�2@�_�Mlk1y��r�3�P}35������̹�6���,�㜎�-Z���ؙ�����GH��^/�����ə�]��満� �*����2���\+�!�'�����-�"�]�I��e��q���w얆I��	���D��%��ڴ�����d�1+Y���=ŝ�8׳�X[�R�M�(��j�	'�)+6>��0GӮ������*�4��"�IV������%�Ɍd����f�h����A�x��T��o3W%�l,�7>�X#�����Q�`O7O��>����E��>z�s�r���K��[h�^V��������ۡ�����3-��i1�~�p����2�1~(^�B���̹�lq�i�JA��.�C���?��peg|O���H+z>F% �9<�
�3��u��|}�س�x������K��b��$,�Ϥ`q!���p|LO�z���X�1���*�$J��4��u.��Y�:�ĤۯDi�roP=�b�;_���X�~h�ٙ��>�W� �'����6��z���"9
��C)k,}ؚ���U�L�Z�v� 4�*�

��6B��B��K�O���'P�8�]��CJqz	�;M�HXlC�3WI4�����J�AK
a�*q���y�B��]4=�[7߉l�y��֙�uH����T��;.�Ίu��/�����&��!iJBn���� �NS��ֺ�>��}��QӜ��M�	$l�k"�]����,sNw�Ψ�h���t%�$T�	(Bo���g�.�͜B?� ���.��i/����6��	�iP�zp���Mb׫*�����T�m\ۺ����\�!qܖ}�
eB��X{�q'��Ro��S������OS׀p�v�~��+Xy;M�ե���Zr_2d�'��y�s`��'��N)� ">P��*PC���$�5����$jsy�>�����!�}��w��5�ƺ�t���w�/���D<ʂ���I-c�f_Ň���Y��u�UY�o��¹�ϼbaO(�V�q=ul�n7�?�K�Q�(�at�E10��Rq��TaŢ������(k��8;G�_�hO�;��)AB�ԫ2n/�Y9Ź��/Z�̦+�	�b�L��r�#�d�h�r�I�f[��1�l0��;��{��\�Ǒ_��H�f����ޗ�#��y��N��{��Y�E���P��Tc��yo��?G�4K�ʟǃ.UJ2)L�߼1�q�H�	4h���:�0!��N���B˹ Y���Is�^Uߪ{u�
O���W�+��n�߃�U�f�F=OP#�_�9Y� {�[�+�����	4��J9f牪�/xg�$ ^<d�^D}��L�\E�����lQ��R�b�;��ߗ�������ܛ]��	���9�6V�k�c*2 Ł��c~$���+Aڪ�IK��p'���	�Y�տH��� !pU��Eda��o(��JD�y!ݱ<��G�_��5�F�{���I%̎�D�ҁ)QF���5 O����*?1�u�1?����Q�s�����ј���_�+m�(I�' �#�.�:ԉ>�ʎɒ
H~]�)���p�YA���)/gQ�	�>[T�
}l�7U:��m��cG�����'k����;�`����8߿��
�gT~���<����e*I�3���[��U���[Ⱦg?��=6����!5\֞륷u��`\)x��g������st��� [��3jBlE�V��J/��b�IF"��o��a��l/}c��C��Y�2�_4thd���br��^��{�`���鄖��~�!_��	�4E�h;��^��ހf����� &�;�e���(7V����
��%�+T��O��ÝB�o� �
2fu�{qWd��D�4ow���@���QƏ��}D���TJ��0ӹv�cmaJvpH$�T�~���Wv^��K��t�J2]p�a�g��������ޗ��� * �/�]4�:���q����(��0W
�Lۿ���S s�ٱ��L)���a�ž)���:P���2�HX�b�Z� ����t������ǦU��QT�|B5�C<����z��Ǉ�N�'Ŭ ��o�u�3|�0�iܹX��� FlpXv��=���'�b�? #m^�1��s!�DuƪA�~�����I{f�oH��ya��m~ܧa��������Yf�ʥ,_b�\�����j��\�O���O.֑D��BO������u��v�i��q��J��=ρY�2N���uT�`�ཛY��l����&��v�c/��*O�����/����fL�&�c{~���z_�g����H�_�y�*�O�����:� �$���i��dH�M������l׹L;��(�ĕWN��Y�֒��DT�����m�Ķ���݈���D�	����+
��R)�&u��|����ʰA��� G��7n"X�X�C�h�z�E���ƽ�"&�`h ��|���I��e-GբG[�E��%�OP��Q�!�]㩗����A�N�֑E���"+5��ֿ2�z�˙�4]��u��y��=��g�7�WSPO#�	�䤉v�e3A2A'�m�8�>����AQC5E��7����X�<k(X�J�}�R�O��#���G���-.g*��Uʗ�]=��L�K�_�\8x��kd�b
���[������{?^ߨ�(��?�kLoÍ��-x$�����k�bA�ۍrV�TZT���$�X�;>����a'�8�
����*�\��I���$r��j� k�a�קD��c!���6�]CGf(�S�� ^�-:;�;�	t�y,� @���,�N�;�A ��N����:����)��$3��s娦�A��8Ge�y[*����/���U8��{��dg�O��^UT �x��e~s_�L8,�Ll-�h�XRd!��e�I��\Ff��T�t�U��+r5�\��'H��50V0�% ���pK�y������:7�d#�|v[�-��˶��֝DV%���7��O���l�8��me�ے�w��a�ߵd?��_�^"߳��PC�lax�*Ր:��T:�-ڔ�͉O*)�CyC��:h�\z@�h�;鰂w服�RҞ_�ӊ�6�R�/al�N�� s�7���$ܟ��O�m��� ����	���ګ��S䄆b����> ���Bڦ�0�4A�~Ψz&��Nu�4��|�P�Y5ݚ7p��ɋ�#��7�
Dq��.�� nxj��W`"r|�0�d�|�㙵��2����nJ>	����_��e��y���~3��xGU�Z����gM�L�|ψ��F^���5ɍ�Y�1�6t��,�;�y1����M���q��=����%�� �+�'d@3�Զ���qd}�K��iM#9��/�-���� iw��#-MM���R(��d�}��mѣ#�����(۞��-֛q��EEbgG7��P{�4���[�ό�����S�ȟ\\u+�2�7���T�f���7�JO�DN|�K��0�:��J�0J��Ⱥ{��3{n�~��1�އ1o�cWa�
-m�W���L������3�@��(�X�C���X���1��A��]
��"��YV��n�%�l1ܳT���9�59
"@���2����c���)�?L�T�-�n\W�\��Ka�3OH�мG����?����ST��2�i$�\{ຼ����-Xaʪ:^ý-��p;v�1���m��A�:ݒ�H��\��J�]�۷M:����/�ݾP]-���q��E�H�8��g�&� W���7�#;�;�EJ2�l�AKe[,T[N���Q����ؓ+�ًC�φ���-|��@�.�.���&[Mear&��I�j�7u�>p�L�}X��A�Y��n	W�Bz�K*t~�����C���tU�S,PU�:g�ӯj���1� ��,�'?�Z�ͭ|j�*����|�. l}�d��*�[��� @1�{�Og!*Q��D�^Ul����)!A���=���R���.�[���6).���f/~J���[��Y��^�M�ڏ'&7����Lӹa�]˅���|^L�5-���3O�"6��������k���5c�Z[��PNsWO�!i����8�w��l����X��p�8�{JP���HM7��{���4L���R|&D�iR�)���"3~9��%r��Ͽ�����K+��<
�FC�U���"�o*@;O\��99�4S`"8�Uھ�� I�#Ԅ��^^ނ�m�E"6���%�œ.v������A&���E1�	U����V�N��j�`��s� ��
�҄B�<�Zk�i��6��'�C.�V��}?�uP�,�O�P�ZFv���#,[���m���T��(/�D@o7�:������<
5�8�7FRh
��Ct��#�{Z&2�z��:ITj�y��%��tG�o�:A�@|>�W`�*����0{pi;����E�鉭�L�s��Ю)�t���H\�u(��%鵧"��̎-��ܜWFֳ͘/����j��&B%����ѥ�/��y��qV��T� ꍕj�͸d�#ҡ��<�[��ű��kt�iZ{�`��I(Ñv�*����W���6~?�p���� �4�ʺ؊Uj0t:��lP��;��xl��̯6�� WX���T��?�i��0,��.�e��
R��|�3Z�u��<���Kt������j}�� ��B� �{w���5��t֕���w3�0������.��WLJt����+7�}/q�A����r���+Fܓ~m7��8&��}QF��1���-��	�lδ�w&��,s�3db��4ٚ�Q�B��i��0�� ?�! s3hDM��ӽ��e��D�������`&}�
�]Ю+>��{��o_��N�[U�W�T�Ӂ�0-0L���-;_��!4SjH����D��M�s�&����O���@Y�1���$�.&�Y��H�����*}�D����k]n5�2{�=�,����c���ng �7�c��~����������J�TP���Ս�N��Ǳ�m8_�g�,�� �v5QRfM<m��Z�+�
)�`�En1*(�ayHy=�P6����m)b�F�]����W�����u'����JY�H��}
�l$a`�z���W���='��$�`pM�uD�����9�}SQ��N�ex�ϟ��M�Vh6���=mC"���S{�̅j�K��,��ױH*�{�+��6���H�z1�]�����W@i�C�~|\yx"�%^ܚQ5�R�C*�
�l�Do�C>#�n��/8ڠ��l� �{h��XEՉ��y@����b�-�q�4���z3����FJ�[h_�78�S@�����5�M����[D�/�"��<�{�^=;k��"���YW7�D�Z��(��Oceb��]��Lբ�VV����l��̒!��t#�����*���r"~ގ�A�,��F���K�����߫IGǛD��͈�_���p[ѯ���1V �-L��J�ݙ��ڌf�܏�+yZ��������5AG����%É�8��`���b#�;�#+�)$�'�˘��u���,G:��an�]�g���$6�u1���bUN���Ȓ���ğ��&zF��tRK?Q�� �e���4��E���%â�rr����X�4�$&+?�,\���N�O���B誘BȜ����V�CCL�!�^�nq�]ӑG96���A�i$M��?�NҬ��UysN_���p��)��B��&X�[�f�߼l�>�|ȗ�W�µ�]���9J�3���T3�B�Al�"KЅcT�_��d����2�O���El�I~j®�.l��3j㲡A#?^�կ-4W-0ŕ�;�?!���I�v�����#D�koKz���E	�9w=�yoMz�9Y7�CL`�
ewD�5�LTS�������p�-�����~���L���x�>��Bߤ#e�>���A�}1��t���h� ��э]�i=w�i���'"J�`B�1IT�T�p�rI5��Ե���I���ܨ���a8�^���bTED�O�U C����V�5�h�i���օ^�;u��ð� !&�hy�db�'oIUg��,	�~�W�!֛�9r���� ��63��2�t����`�ƫֹr��em�����uUb^����q�*˄V�����?�)����N)�y!0�0	�yZH��<⑹̸_�̠?i�ZR>�-߅C�?T9`��z��{���ܔ���:��A��	,md�պ8�Gl�0p�������D�MDG?tKP�l=�3��I� �J�w?�����~G��M}B��0��T��<Ԃ����c[��-ށ��9��m��� F\��wI�h�+G�v t�h�%�Ї���S�.�e!ͦsI�q���&/��Os��N~���T��_���Ӎ.򪤥s�Nx���䯋�%Z��-h&ú�'�BaaB)���!�"#Z��fϾM��U�'��BC�-�/2�m�a��_Z�j-=���\(x��
BoJt�N�t�Q�U���mԶ��N�:�/8�&pW��m�������8����bw�����1�=�~v4�f�- 2��_�E>����-���p0f��T��K����N�	xc���ٟ����L1Ky�k|fZ����1�Z!]I*�1��Q��@XyJ�E��#E��q�A]�Ƣ�D�i�֌��-Hf:��>��I��8y���+ةƬ��+1MDdݍͩr1TFX���O�,L�������]�ʡP��0p#Vu��;?R!�0I3s:�t�ǰQ��ƪ/M6��2�i'���0��ߟ�l���{�ē&E�L���TM�
a�ؙjR.j��"%bsr枟Y=���	! ����w+Y�[]F&w����J3�:_�W~�$����v�,Q#}�R���Mjyzz�N�����P��-�eTV�5{�^�|UW��2�a�~�4� c��#��E�S]Ca�R눬�m�������ӛG�v���OZ`@(m�H/�9A^�"媙`��>���(���@eAv3ڲ��ʥ�ǚ���,��W�"'X&4�K��6+b����*miڳ���������s�z�,�+�Lm8�x�\Tظ�ic&N!��F/�l	L�������S^�S����ݓ�v��������f{�S�x��Ŀ��/�3j�=�U��9�q��/����ǈiS�;�LC�lc��g�U�9�?+���̚�R�U��}/�^��×��h0�R��z��VTf���^es�����|���wXg6Q+��O���.�vF�
��p��#+���,��q�����L�x߰�f�f�HKk�?ʧ7�E�H�)����h����P�C���o�\��T�
�Ȗ����R�� �����4� ����=>�{��D�����g�\��M���*g*���_* ����,��T٧;߻���:x��\Rn���!90���Pql[ h�0��)�,�I"v=��e��'!�~�ޙ��`0r�Gb���V����VpB��	��7[���h`��9��*!���� (�s�?:^T�%�����N��1!G��F�wϫ�Y>�g�͞2]��ж�U*m��'�kL/r6�Ӎ��1��I����Nn�$��1@�p��b�1����m���8Ï$��q�|�5bsr�Ls+m�%�ݕ��M�u@�ȟ�j�,	�����`��e�Hg�D�^~CsŽ��F��+Mu��ӷ&_Q�'����D�Sw��P
?�|Y7�b�D!�<���������\�K>Ҁ��?^6Ѽ1�8qs��3�������f��ۄ�0������ͦBF� ��!<������t�ب#�3%�����!�t������Z6!=�r�.��ڤ���F���,����˻$03'����Y�r? ��J��`x<��8�)����)����"q�2��u���u�vB1�����+��Fi�M�F�i�����CI[|�C2y�r���m��K"Ԅs"~ZY��!M$7c��l\��J���6?i�EGz�,�a�l~�%����$�ꏦ�N��ӻ��BB9p��ˇlϨ�EoJ+w֜��c���Vv�Ul��ޙ��<�/�v˒�bP���n��$��P�M���&�YG�J�=��Ĭ�ό=S��O�����h���Ͽ� �}��y��;&U-��v$U��&*+y
�͇7vbT/��1+?7���F������?4����9���~�r��鯱#��-�P���s�i� ?��(/;�<@�����(s�v1Kn$�j{F#�� :?wZ������^���3�V �i5�Bz-���Þ�@(v����,M,l(n��R���ţ��t�i$-�� Q}H���p'b;(FLs}'>J�벗?HTh�d�n�@ϰ�ZW�i��/�j%�<Q�k)���qS��l?Ů�*7l{�����s�֊îj�s��ּ�]@�q�}E*�A4�Y���vfx�{�@���Q���{�6��Jx���D�{�mh��	�|V-�uH2��n�t�Q`59�T	#�9󸫭)�? ����Y\S�~>��T�H�ݗ:B��м�ۍ��ǌ(4=l�KiTwF�n3�}��zZ�l[U�v�\�*��zb����6ɫ���$�,�z��x�\������bA�)�直���ט+����Q�#�1�=��9K��\0�٢�5e�saL4OI�.�5�-�M��Y3��*���7��:��v�>[����(Ai��e�l��/�ݧ s;5W*v�%!�\��>�s�~Ö�Q��V����k�#wA݊��/P_�Lʹ�>���zP�?Ց���{�7_%�>��������p4�}���YҌ@���|gTL��xu�,�B�z2յ�Q��� �WI�����q��t��4c��	��nɢX�wG�9[�i�	�өZ��5gX҂�,�9a�r�?�p�-�h�V5��q�2VY�-}����Y�+�`k���*c5��Ro?��[0 Jm]��f�<��'�
lթ_���K�����go�i����6�ag�ޏ�5j%D�:�n�]�y̴�M�m��G�� �X�
�4�\�`,MU��	P��{��Oi��h�`�Tf����WS��e�W��(~;�<dz��H�lMָ[�B���޺e&~��/S`�xLfؑ�Ï�����z�1����՛,��"�`�J�A-��zo���T�.t����g��aq����)�hYGɯ�"	�����}�^s*i��fXr���4F��-R�?�`�xtz������Ɖ����AtJ�i&�h�ki+�#p���Cy��-uq�p�i�!z�p�����}Q}4��Ɏ��ׄ�4�$G�S��l��,O'p��ÃTm�r�ѱ����8�i�p��c����A+�ߴ��k���oڢ�Ցȱ�.d���+f-�=;�4�X�[�_l{��h��H^c�]����?u�ҵR�HtD����ϊ��>z���?�?�m9�f�2��Y9!q#�4�ʩa6�㴻�����8�_��.�ǩx�M�i�:���B�:pB�s�TN�1j��ׄᬚK�/�X�:4d�p�~+��б&<<�L�a(��O��üI��fsj�P���]ycF���ǅ�/�1���Vg1�{��'j�!��<�y̝4�)�k�o}x�בU��f���Γ�X)	�dx���D��[�-����K�O�8�d�~{���A;�O� |+k�R��&���m:�n��c�\��0���'���(�J�T���qN�N����\H�Xd��ooX��5�
�8�{U4�>{�M�d�$�0͇J����s�Jqͩ�T;�x���jc4;�S-���u*$�k�J/�ǎd|F��J�C����rҿ�Q�'�z�PLˠ�'Y�ӡ	L��%��gQ��0���[wuDv/}@'�F�\�e��8�2�<�o��a��C�@������O��7W�!{��L�_��n\L At��RmA2��M�3;E�tyI!�nN��4��@V�浈-,�i��/\�"�J�pvpj�����\�ձu^n������.4�j��n�ׄh�����ޭ�53�[!�������ۻ�k7���kt�7�'���E^ ���#�ܫy1T��7�n4�)V��u�@O�ɴ�ǩ�R<$a�Z�c�|9���@,�8�0�{y7=v]%d��}(�Ȫ�퇪�vcY"��
��S�0��� IwRf F��gĽc�(��⸹�9 �>��Ǵ�p<j�ڃ���;��l��7�[�_�ޅ�ԄJ���}g�˖H�_HR�Vb�����n��g��b�{*Z��(B���{��s�;����JH?��C�{"~P'҉��͌}g�\�̗�~ea��g�
��+�Ɇ�04^$��<�͗�]��-C���U��Ln;�(va¾<{����4)l���[��Kg��e��������h��:_�O��hVu��30�N^��9e�󥜓'��L�EْĄ�sӗ~�&��IZ����rEV.D��Yj�<�W˲F�s����3�^��m���`�_�]9���$�a�E������>���<=�sҖLhOt����ߓ�c��`�b?��ݟ�K"/�i�b{��[�3�B��G-�+��N̗=!���W�%-}�^eP�b,��W��'��t�KH�|ʬ��y9B�|ad
�>�^�����t+�}[����E=L�2��(qH��,Ά��a�֊�J�.W5x��O)<�b�����n{azX>F�'�I��M�Rt�edA�]�\��dZ�Xm]�?=-��u�3�pM�k��sC�x� 	��6E���E趜�xI�NI\��.6�������z�d���g���G�=���#����Lm�E�t���ז쩱n�U�� ���b��#. ���#�&�A8�k݉U�sXrb;�Ԩ��g�8�j)������e����T���,EN�N_m���V�Q�.���	��2/��������8�k��Y�+�9�N��8z�[�����x����rq���X�ctƨ���^̗=�)#Y)i��b�Q����)�����tO��H$��&պ�_�z���]�>%�g�<�z=��e� ��.��֔�E*���ì��pF�����U�<�<��cV�]є�A�օ���̕�8I	��6r���1!�9�b�f���lJxG�-H����E"=gM�7��i(�7�P��"���Yn���.��ӪL1݆zȞm)qb�ϭ�~�b�]	V��0d�e�;>I���&0��$ރ?� +�����Sx�-��!��/�������L��zF� �������s����o�5O�i�W'>�O�Ug�B����NLQ�IS��k�б&��q�F�~2�C]�e�K�PT��3�K4����J����gVB:��ɼ�#���q�B7�x�	�l�3HeEk�D�l�#���o��L*���F��j-�歎�g�c�,�*3���C�xc�bs8>n[k��)z�.�j����"�C�������u���y�{q�"ù���h��i���h���}@B��&i'L;��q��C��U�$��>�X��.F�Gn�aE|�8��j��_�p@g�������o��o*�`�l<nٮFɒB/�߈W�w ŀ= a%�E%vQ+@
gt��Rﭠ��)Y���FS��?a�g)�����Xa��}3?��6m���P3��YgI��r�4!��t����w3�8���I�z^,:T8~U�\b����0��:;u �Ne�24���� c_˻Z���f`�9(�H���rw�P^v���P����CB}��-��P%��(��ҡS�('j_1m�4�j���������_�Ӣ�ǣ�-����n+N��E�ФA4�d���;5H{4��7V,3���~����n�q�|��*�_���[��ǃiGT�cV~�@8ܴ�
~�e{N5�ї�F��d��Y!N����_��\CюP=��ƂV\��җ���cL���8{�-y8�z<%ɿOm��ƌ5�0�s����L����]���;�awN@��a�.��61:�\�&�O�

ﶰ0�΅qW`N$�\�x��֫���>lu	���@|�����Z���2@3�wlM�a`<�6��FX�M��$&0��Į[@-�� �"A��
��\���hgi�p�/dL��s-wms�͛v�!%\�l5��I������H��Ģ�T����m���G��q�i����y͝ߎ��>�ƴ2YJ�N�O�ꥤoT������4~2w�T�)�A]�d(+�;�n�����E`L��F�����)��6.�K��-m��z4��%�P��^>?��z��il�����V�Yxv�3�B֓a�����g�=������(�xO߁�$�|�"q�.�r�%�KO��h�qGmה;�g�^��@��m�Mr`�xx�jj���c7ʞt�w��"g++ ˑ
K��f����fj��J�L_��<� ?�#4o��/���]H�u㉤X�ZfC�U�GDw��'�A�g�	��R��Jv,�u�,B��E��c��Z��8l�>Kn��
:���*\4� ��ւ�{n�4�}6�hűZ�g�X�gv'��N��1����z�孥7�/!�n-Z- ��W�=�������=����\^Q����u�\t
�f����C�T�6��L֌�����cm�M24m����*X�6M��\�C���="�sn3U%��L\_��sO_L�����s��T�h�]au��F}�m�MN��Iu[��T����IV_�w�l[U�lk���'/Y*;�������x���^�',K ��I_�i�ԝ�iK����g(����uw��Q�(�3��*�q��O:�gt�u�����y����ˊ�3w+I0�@H��� �����2�7'wF�2.��G#{�Y,�1�ʡ��^A}����bҬ�e,F@�,V�+{�s�� # ����o
w�$^����в�hX���nbMgF'�O�	���>�"F~��ѿeL�rz�~�r!	��Ln�`lc��^�s)`��z�t�����]LϏ�[�(B��k���^���|_�g�{NW��K�	�f�[����G�Z��rD�u�>T�{��MHFG��1�!uPl�NVs?��a��Da���D�6����P�RG@��7�b�Ǯ�:Ns�t�F�K��z�,;5�i3��M�{��C���^e�����]���ș8K�[#�t%�>���jl]P�'c��;�٤�"=��|�zߚ9e
i��>;��I�]w��k#+��r���j �.�u7�u�RS0�a��j�Yz��ҁ�W
�9?J7뵹�h�j��JvZ*@�F�>tg�띇?+y���E���} �qSZ�&|���HQ�%		$�bb�aܥ��)6y%��^3�컁Wi>��S!�
�-\�ߟQ)I6��x��_b)�	w���n��Ɣ�@�i�~8�g���?�����ba��KE���Uᔕ8��D���k�#��&��14}䝦�냦�����e�,i}aא�����#WpQ��N�#^��� ��<=JX�~�/(�A@>ڵzB;������6��Z��mþ>Q_���*\[,��|�B3kz]�-c���c�F]t���_��uh]�͉ae_����C߯ f�u�ė[*�K��\ ��Q�9R�ʞ�w�	�v�Y���g�)�6_�.�j��K��(�m�'ҁ�؀a�mzr[.����;�/=�w
U��&�Q����E�5�c�����&k���$I�ai����akV:˓����)$Ą��P%�T�K��Q��$=�E@Z�?�ĥYW�b<�n�-�� �1$VR�d��l�@������;wU=�mJ.s	�(��5�;p}�X5&�:̬*ƾF�m3�#$�����ҽ?��Xyk�$6��Z	�U���+<(�(��蛇 \�(Ȟ[~�,�E)S f�f�w���P� ��(�����K*�M����X)/��$O-Za��~;�S�XE�,7�F,yGj�T��:��f�^ɏ�p�2�UmQ<������Ud	�й�f:�����x����pU����!v=rQx�4ڻ}�|c�Oq�n7�F�3��>azI`���}���l���,Ԑ�:6j_�N9��Ƚ�Rg����Kp��ӝ���sq?@�~V�utl��,���5Շ��_��({��yo�^�?��VLZ�}Q��ݲxј�3+i���hH��ƜCb_tqq
7�B�42L@��ۉ��&m���;�B���!ukHB	���D�%]I@�z.�j��*o�6������_�0[�0�ϝ��|�qe����.�-m�ǽ�
o�]�Lry],��oD��	������SQ.:���]`〯�d�����x�������gƙ �;��qRs����պ�ZG�k=�ǆ��BX��CS}jRc��7���h�I���`aENg�0L��͏�LO�v��6F�3�����N-�Ƹh?3`�r��=x,�&��eg�%��m��Gu\"�{��ӛvT�L1��5����
C�!��4�R���*i�tǟ$��*Dp$r �!�����f����)�^�}�e0��s1��K˞x8aI5���2��gr��
�me��vs���.�wy�7�!�ľ��d,�������||��W�����k�h���u�Kb�w�lw1I��q������z�H[�6Ƌ����қY-sf�{��Q�/����i�|y[+o�a�h�U��K�l�/T���z�y\Sط�5�O�i^T���,�_P�ii+$X�P�?�b4��+�զQm�
`��t��>�m�;�n��L�V-����>��.�3�����tF�PV���b�o8T����'r����Ȍ>ӡ�PC'��i�O�E��;Q�wwBۀ��	��̞3MF+R�4Kˁ�,��4�~���e5ҘS�x��@���s��5^�
�PO.ql��P���$�/�2�HBs}�1�����C����Op�	�b�����7��qo}��xy�uR=I�>��n)nϿ	�<�q�(}�ߛT��w�lo�ϋ"�r��y�*�=�ޗ�6�p�R�,)w���Ϋ�CZ���>��;Md5��VJ�/y���4�p���t ��9�=m?sYc ���.;"vv�^�k߽�Z��N�f����,D¸[r�iB],p�褠e��.�5Y����;�+˕�ixk�I� �7.I��
]�4Y�����-<�;� �k�� ���7?t��o�j�a�̴�PgQ�@�3�1�c��$(jb������7�9og��3	�����}�z��(�8��K���5H�"���W��KŚ�P�1'O`Q���gH<!{e�m�����2��a�Wn�D�#S��+2�w׆�ݘe:�>A�)T�l�'�
��jf��ٖ/�R��3�&;^��U�N�R�f�c��#t���͉�Gky�Z�~F���uO����gJsP��'�
��_���Z�`֦��n�7+6.G���Eɉ�!�8Eۤ���u�x!L�3����\���&j���e�4����(�h��H��
���k��Oq�.���S?����0�x�`_����$�q�-�W�����]�;�ԃ��CP��� ��e\1p�4��i6����M���3������^m�L�.������G���N���V�N ��/"Rք=)��E�AW�oB����,�X����]8�D��:���%ϧYd4������O�>�~�y�V����W�v�1�o׊�7��d��X۾�v#~�kX��
'G&6x�ԬM��O8Gi��]],5#���p�ۅ"��54% ��"	������5�7.���t�:uE�r��t
� �Uo�Uc��сl�}�v�f`�v�OI�����v�B��É���Դ?$ukJ���O����Vx�6�Y(<�PG�,��ta������u)��GG�!m���*�J��N+���\�K�N����Д����-�1ʊ���֗�eo˵��Z�O[��>�5/m�7���9�!r�U4k ��N�?Y�,9�A�P��W`s٤
t���C��ټZ�n��7�o�݁�vxG���}��K����s�(I�gڅ	�v��c
�'�`[��)?6�6�&���.�ag|�1>�[]��T�¬Qm��ȼȾ-n�:�yDuv���	�����\ �b)�d�=qI��	�f	KĶt����r:u��`���~q
o��ޠ�Ɯ'=}�Rs�ǩ���l0a�f��@�l��s��=m�0!j������S�YQ2yLH�6���Ԃ���I�����8�����b>h�47���i.B-�؇v ���J����l�#�h+�I?�s� }Sw<�rN���#�z;D�����J�\��,��vY6�t��D�EQ��bE�p�&���R���$���1'>���m�#r���E��>���,;1����q%�: /����G~`�_�l�ʉT�M��ø����|eC��Q+Ě�I���'^���έO�6;��� �<"����k���ZA,u[�4�X�!=��bڈ�rӑ�%�٫���z�����TH\h�p�\�����˷vh`�jt�������b@�
���-%P����L�	�-���'Y(�@.O�޴�x���t�����:�nM���j�ӽu>˧H����ұ����Џ9�N=�:�N|�ߠb��ZX%��]F|Y"������7Jitr��L,���z���>�������2/�^Ɗ���S8,g:U�?������o6+N�����s��n�W�^-?tD�2�������Oݲ�p�D<�A7�W������R�2����7L��5�Do�P�]�h%�d�9�Z�KF�!�]�����V���5�X3L��Z2�9l�\��.銟�l�����a�'�1/������ϖ��ߝp���8Ir^_�ґ����m���z�eT�%�J�����[�غP��H�B�~5���������p	���Y($P5�����M�* (==�w�Q�SM����Dתy��d���f_�)5�2���h}`�S��f��Hw��Z�XxD�6gk6�A88
��}�7P�)?� �-�4��ϻ��$��ȅ�>�H���^����1��}^���,�d��'CP��C�:;t y�K��<�e��'f~�(r�IWtnn�������?��t��ˢjkU�A���Z��n5g�$��'���sE�JC�ꎱ�iZD��`t�.͋�7
�����<��am�iϓ����� �>Ze��GdG������7�۫��EWP�<9��ֲ�ge�]q=��'p�.�f��bx��(s����["�.�=��ި���K��H&ՙ�������E�6���n��� �Ȟ.1s�R��(�
��]� .B�LD���Rч�oA(�������o�m~Q�x-b�da��ƺ�M��םi�8������jigB�����0-�8���,p��-k�"0���� �����ګ�q�J,W��E�װ>�|��a�qn$B[���`�K��`t�[&�f�;#���D�n���VlϭM�����D�)Sc8\T��1V�X���A��/��Y;�B��w�3���)!b1R:�"��[������r���$�Û+�f��9K'����yV����G����Ų� ���¦�v[������k���_~�|������������yk�e����ì���I����f�8l���>�;8���K ���xvۇm*��f�}P���t�+����s'��^�YP\<J��=>.��*�Jx���*��/]���������E�Vq�wC
10��%�*���qB������+r^�d���� i��z?�?�'����ǐ�=��*���0 �2KV|�����>�D���1hx�M%�dxZo�"��fL;�ZsPS��I��FSv������t-�k:�����)u	a8���St�z�B5
��^�@ٷ�?+���¨��?�R0���)�s�	���"�9�Du
'o�ĐBBMd�#���	��,������Vb!�C�Uѡ���y�u�YxeºG9���?� ZO_�\�"����;� �W�ڏ�����P%K�Af)/ӘK1ڲ2J�B�]�i�u`�|<�򈞅Atu��� ]�ٖ"j[t�j�
n�i�	��Hř�w��p��\HO��72@���T��tS��[�Q6l[�]��1 �Tu�
v�"˔I�����������J�郗�Y���!�ʿJ_��%\e#���F��XY^�G��5���kk(�����u�[�����r���\�߭�c�Ү�18%U���,���h���� �Ss�h��iFXL}�%z*�c�t�XhL��!�ꙡ�Q$ oDJtXO��vF�&����I�U�r4��v9���4�t~05�y'���y�L8�L���"J��o$$i��`ݾئ��΀�2��XU���K䍳��l������qzDw�q��⠾"�� ,>��ݙ�.I��ڲ{e��ssGu���ƪIf�?k��[�Ϻ��$aQ�V`jpi��o"���|��]��7��yp��oZ$�6��!�>#�	�Nn��0KdT-3�q���l�=eϷRd�y�3?\RY݇*=a��z��X��m� $� ��O<+ub<7|?<<Ɍ�\u\�m/1ϧ�i��߂@(�j�GXk�	��o��1�b�K�+I<C���#Y�T*�OQ�W�L�o`��d�/^��^S8��;�u,Z�ct7g�ϥ���~��+H-YE1�n���*�JR33$[�
���{] ���?�Qlh	�u�]���:���a���$;m
�
_�cls�ɺ�Gƹ�w�#9���Z���yY��Kz�C�&�-�+1���~�8��B�*˛���+38�n ��6H�\����^;)�ϻģ��$�\�x�'/��}���Œ*R����gOGP�$�'ĚB�fP��zoV���w�K����6^1�1��"��H���v�dQ��o�(�-� 	�.~��w�
U�b|W��mE���?��s�98zMZi3�	r7��c]��D����h�XB�,9������}��o՛Q�7��QN摕��3V_S����W,b��������bC��O*�Ϻ>c��v�5]���s�X��d�עo��_ӌ�a�U�}��<]E����p4Z���j\T��g��*f�R��5�0RK�q�fNfAj�O^����zT�m�߆�=z���#HCγ�g���k+_�������G�f@f��NxXg����I�N3�u�0��MZ��Ɛ�'�>��
��N�f�0UsB��I[$]������27��'u^w���?��E��?	 >�@y�tޓ�F��t��Xw�����"�c�/�����%�A(1k�m+5H�\4o:�0=��v(��n����$|3���@[��9�_�+ ge�)~��Y�.�&�����RQ�ʬ����=XCc	�%��C
�[k���r"{Ў2g=�#bO�$�{�˕�U�|i�0$%��7�{]��r�/Ja����,��؊�-
i�e�bw]�#�cV�Y��dU��.Wհ�+��b�J��t\>��nvc��D�i�Yۮͧt=J~%�|�ք�Ih՜0ͼ������xI5���5q�x����g�vE�����Ë-;Qäl���wcVcu�W�o��fR������&�F,���,�\W����<�P$�[-H�ɤ�_���U_|�� 8����F�M�jCL`���zS�'�0��p�l��Ӏ �M�㸼�g����껂0t�ũE60V|���8'Y���<��ʠ���#3������e!f6���A�'���j���:%g�����{�۾&��`/YF~�L�\Kz�f��X�#﯐��1��SIYv����=�8�R{=�Y��t�v��m}�=Pϫx�y�%DM�-�����zFX�x{��~�T��ł��}�+G��.Td���n�I���T��H>��8���)�,���Ft7�*8R�0���7$7�Ϸj�p9�9]���9 �}�U�#���� !M	s���:���@��#��]r�Ɠɳ��[aam �0��kR0Cj�J���3DM\ѯ�y98���+٧O:����R��
��69A҈�r���)EQ{Kj[&V@h�m�K�Y�&AnAz�%7ڵn��L-Q����ڈ�F�*�SŁL�P�JRJ�䓋�PU�oI��O�����>��^���M,h� d<E�x+��N�E����X(8�t��CjI�fh�je���t�nV���k}����[`x$�gd�芬�	s�yzyQ�ƕ��R�y0��ߧ5���a��Ϸ|M%�g[���L�:�c�۪K��qܗ���E��A��غ�y����v�]^��s I�+���l�l�W��+�uI�g���F�U��Wq�M�{�{�O�=f��m���rX�B��	|�0��df<�^Dy	����,���<WmQ��W��}��٭o^�
�O#٥�<3]u ��a'���*����rTR�"��.o)_�_޴����BS���w9��c�?c:�9ZZ{�QY�d.��C}Ī!|���Ǯ&��fv�`�L뜆�A؎��Σ�v�Xđ�/c#+6;����q��W=I[AW��<V��?���|�Cb��+�&�-t[�,��b0���a�C��N��Q�X��O7�违�Y�'�d�q� Z���Cd���E:�ضG�p�{o�Z�h���S�[P���R��_gD⡑6�5w=+�\(����$#���&'$� �7|�*gR�HV+r�R�Ԅ8�:����Be�/IN̙�vdVٌ`�CcH�.���r��HI�! ��1Q�}�ʼH��Y6�:О&��[��y)71���
#f�tx�>���w��I�J/��h�-<�'����-�!:(l�0��\Ԛ�حA�;�[�e$%���� �R�"�3��[��6�(f�hB�.G�#�!�0����g�^ȈiX�E�N�y8�aHz]����e�����b�z@Զ�y�-�k�����p�$۴��ʣ�8)�#;�0����~l�8=tXj��>9_E�y�xv�>Ӱ;"3��c込p��;
�\'�+���
��g'���O�Cv;�*92z��lƴ�U��+uR�D�N�бZ(��W�p�v�nvঁ�d(��{w�N�A.��������m|;"?�K�θ�k~���b��Xb�Ϛ��(\�)����ۆ�?�����e��O[$���8Ԗ�=R@e,[D�	s:�,���ќ��`*k�/�p>��$�c�t徜T�<�U-�?{�J�e���3D�<Sj��B���6g/݀'-?��&T�z�1~���&��b �{w^���������!�&�9�A�L1�,�s��S$r:B�7�GI��˗�2�'�P}Kr��2}��@BCNxR�'	з�5<f6M+Һ:]����"h�$�҈����fl�G����V#����=���]O2)X�P#?�(B	A�y�x3;J�\�"=�_�ٙ|G�P �?��
g`LNy;�$�|��C`�.��_��/f�Q��	f��G���s8mpeYp4"L��w��ϯ${򵈫�4��Ǭ�Tq
�ߌ����v/
�����
˓������$��6l���6`���`�����[�i���ʓ�E+��ҋi���J9c�F�ޑ�Fw��-���F��H�Zh ��2�ݤ����-e�����M梎!�$�XՄ+u��@�Q^n�RE���9��k12l5��<E�C�!�>G�=Ev�����'-i[Q����-5�g�@��D�/�}9n�����Z^����t=HHî>�P2+��l���z�*#�'�[c_�%�y�J��D.��)�A�%ee��b�]E�P�d��˧��M����גּ��(��H�c�q,�5�q~C�X#R����j�v&E����68�.�4[���z�*<6���ҜDS4��9�nEA�6����y|�g�ODoW���q� 
���<B�=�m��HN���!+p��r����3QZ��c񪹏�Ϝ�iH;w��y��]�K{�	+i�W�R��j�|z���sw�qK�,rJ/������Oإ5˖vMAG?K8Ț�%o,_���C<Lq�:c?�r<��:5L�-r�w�㕋��-�Q�g�!��w��2|�gGd�-F6&L/J����d4��#�F*�X|ȫ����r�	u۴#���Lq��S�X�U�+�|IhwEM�j7b�w��{�ŧ���3&w�aܷ6�R�(�r"�����i�̛��0��Z���I�~k�&8Va�q�{�~���J�����:�jܥ,���_(QOQ��{�Zt
f?���c�jn�=yMM�	�Hl�Lt�Q�g!�&��pw\��!�4���k�p�P��a��lXeE�]-��F_��I��^�L[ox�rm�ƍ�a�6lR�lC���3���򈻋q�ۯӑ���um�o,���˫hi�N1��4|�Y��z�M�R&y��͚v�1)y����U��������'Ǡ8�k��s�&׭��T��j����/���(��}�h�S�ix�
&�?\��\Cz�����-��[�.D�4�*�Aͻl>�dT���Ӎ�V&1/!��$���,~p-e�/s���ǒ������[��(��U��9ϣ�S/�߷�; %Z�)�S����LJZY!3�ʲ��iH��I�4Sp|�Hۈ��W���i��}��q�){(%"�����U�$�Or�:�Z2�T��-���p.���x��ڟ�jU(���y�Y��y�:�r�9;� &L�q��u��S%�D�q��N�(X$�eM 	v�� �xr���W���H���Y/�$�8��)�(���M���c�������x�+�鞠��b�ʴ�&1߶����C��6��:B�����Z.&[��J��t�Z?l�M�����lr�FV����*������֟v�֭Aӓ�)|��R���e�e��zɹdX�lh�w)�0c�n��0�v��Q���}���ģ�^���&tN���r���-��D0n=i_"e�a���x�[;���Y�-�|����
uytr�TԮr*���_��*҄
�t�M��}�E���E"��{��]�6��V���X �y1�KaZG���h�[�(/uwY*��1�c�Q�i�G �B�dP���㾫����F����x��u�`�>co��p꾋3� �6�Y*��=����m��S�w�Tڷ��[)�"I���x�c�Lq̓0�,�s��#��G:�����~x#o��B���7��h/������d6��(r8jb�z.�ڦ������][��
�� �i��}�[/�_�P].=x��,�{τj�D���5e ��Sx��k��u���B�V�=ym7���3�0j��6{Y���JR�TY��B�J�)��`�۸_����Cc�%�-B����\�D���'BE3� ^�HBA���S;���]�Du��u3�u�����A>v���وT��w-��AX��ɫ��8��n\�>dyO��Lֵ�jG�6W���b���6X!D���`I��κ�'��;f�9���v��Зk-��c�y<�9�Q���bk��n�5��,�oo�M,����DMg4mt�)���f�[d+�@��*�3�o�}0���cZ$_q��`��/ؔ��^�(Q��NU��W$�4�`��E�	(D�����Q���U�y�H��5;�C b-���0Â�?�u�*:֍���@WHچN�v�e�dQpq��1C��}u@*��0���/��f�t���s��M���S����a�4���f���)n q�`�?ȬÈ�#�R�7U�ОE� =�Z���O=��]�DGp�4��e��-�g4��b���k����&�s��x�"2v���Ҩ����L'Թ�oZ	�-@��.��[͞I�����K��Ʋ6
\�����'��ϋT��(j��p�Ms��&�"? �/VJP%!l��]u��+�U~z1�݁��� ���@W��E�ч;e�1���Ql������0��k���D�ր����u�}��w� O��i}^𠯐��P\��=���V�0�s�!��vl]�k_�9�1�T�ݤ̬U���G�:�:��v�prqs�1�\i2녒0zg�i!�fJ�R
�_jV;r2f����9R�H9b:8�P���E]~�����"�@4^N��K5��{{J�3U���C��$���e?s�����mA���4�-}�<���%��گ���i��[Lf���#l�up�����tlӭ�FX�������`��1GS ��/�T���-tEx�}Y�[Y�)���R^<\���Y�K��ƙ�B�0-7��P5�?�&�G��D�L�Hcѷ?�BAG�+�B��Q�_Wp]�e��K-4��L�jiRYw�
O�s�[�@��h�����cg*�� @�#�Þ�N�����-�ƻ�;��۾���ف�Y�[�n͕szZ�l*�S�OV ��ŎH�DI��j\���cqRB�r�!�o�?Ps�g<4 ��P�+D�!�	��l�������e�. ��T"��:i���y��l�������Y���,^�D���L�e�ACΈ�^�Ї��'�E�n�K����va�)~�)���d�\g��RÓR��z.�wu��(/-��.w���b�C:���kޛ���t8��ZNX�zX���=�ڼI�k��{Z�#�f�Ie��_�ߐ�����߶~ �>�\>��m�<O�M��ڄ��mlu��Cr��B�YH�i�@��@.;�(�~��y�F�mj�D��kv���6%�*��^h����)�a��T��$��
ʹ}b/(���P��Q����ٙL�"ѤO9�aj�Ur�#�n��v����[��FuM{Y,�#�o�����PD�f�h����m��7·.KX9V��$�R�T��\�W����.��S�=���an缙��C���}pw�Cu��d�]츢>R�B'�I����"^���s�*٣�j�Qh�Ǖ&�u��pI��i�x�}�.l��YQ'��(4lŨ��o�kw�Ι��Z3�
|oZ*Bu֧s���O9� I�G բz*�\R��?�Z���-s��F�l02tܩK�ͨ/�K��l51���o�Ӝ���K�.A��bEԼ��,� %!z���ǉ�ֶ�b][M������]Bb(��m{b	{��|����D���S��|�y ��\��@��q#�s�.��f\l����[�=b��qU�x��[L�(��g,�>�%�܆Bn��y'��=%���*~��!>Gb�vh�W>�2���H� 
�����|�c�����f��4��l_f���-�3!��ԨA��i�z�VIX�K�~�i����v��Bڑ�%��E����%�G0��F�� ��R���Aw
�5����2�ꮪb�|Hzw�y����5�fB�5���O��˝;gB퀺���ۋ]�k<�O�J{�{�r�]	�1�H>k�j��y���5\	�$��9UgƔk��S+���ذ�\"��K�S����Avak�I���?�Ӣ�
Kv�w�ѷ��OE)�X����ND4,���YO`ΐ_���yW��»�`q�o^fI���c�|s�	��y�?:$	�#�rj�'}�ЈШ��te(-�1�M����r8���[m���<���u,�Ѿ5�Ǯ�%ws���BNy�_f�Iߖ�� -&q��|��&$|Sؐ���](�=�n��X��`�b�mkHG��ဲ��6}�t|��v@	�a��� �*D򥇀/T��φ��s>�C��$`���!��5�	M��#��VE��l�3�I�m�<�r;�k��t�Y?󮪧�X�{�A9⚪�'���^��VĒ�$�j�������C�ꗐU_z�k��8��0i�m�S����Ұ���F؞(l�J-)L�a��$�P��+I(�i�|��\�_�C�������4���?������ʠ���Z�BW=xm�˩��!a�����;/t�%t0���#��8���C��-���/���W�{�Ou��b��R��`�&�;�y�sN������Ɋ9�V*&T�����tk�����?�Z�4�0t ����I��MII��:\�9�Sr�,g�.�.��
����݈7z+ع��6�S�Z2p(��bm�Vz�4,q�n��T�P��0��!�pȗ����7=���c�E���ta�����k	��3߉s�[�]��Si8Z���������S��p�U��f�x�Y۹װ�Sb�*$;|�A����ΐ�T��`Z�(=Ā��AiJР^6C[8�}`/��I��3���k�o�B�$-^�#ݫl�߱ɪ6ՏGd�.�3��:���� �����y�Y�]L��[�>A�jQ������:�76�o�-�(���6����ucnq�>/�Y$]���Y�A�s��ڢ�| �(��'0(�^a�`ŔX�9����L_����80}6����2��[�x-l���'8�%1�@wJeA~ ��jm��8L���̄�ǔ̚�cT'�v37�����x�
4?�8��%�٭��x0��ٰ������ph�}��g�|7g �7���%�����ۅv���-�`ʅǅ�Zݺ��;8�>A��'#�2�W�|�����^b%�C��??0rӞ�b9^�g3R2%�v�3a��w9��#_�;u�����&�p�;���|���3��� 3����(�NEŠ�K"o[�N����@g��=���|�t�/B�z�\�x���4���#86J6�L�$��C#�ѣz���P��@r������s�qcߌq�=_��(h�^��Ȫ��/���j1��d|����+�ȏ ��%w�ӃSgk��4�U��ز�����bV�e���Q�F!xoi��}��sT�P!�jN�V��\~j=� "�y�fj������yά�M��<����N&����h��)�R�U���Х�����V�IH�6�u�0���k���1�������P��׽��KC�3%��c87���D���=�K�M�������I�6�\��z��eآ���c��9�"��0b-���F+�&'[W.g+��3�Ssx� ��p6�����#L2K�\.tuZ�Ӊ$L����4Tn8��B�L�<�y����u�$'�mEbbKyw1�l�`o+�W4h#�Z�������T0��x�ڠ/��ܞf u�����X�
�jjgRSU����r"_���^���w�B#X>Af���u�`�{����$˻}�7�q�j�&D�\�K�-h�Z���DU�V��ҫ���cK�M��:�����'2���\��u�(��1���l�ǯ����w��M7UzY-��8P0�	3Wq$��qϰ���~3��mUm�"�WI"	[��p�~����/�H�>��W�h�E��JfG���������e�l9h�łF�Ό�6��1�ȭ�f��nD�����u�<���� �L��}f�tӁ��j�b�[l2:��)_�h�F^J��ګc�/5=}������G��`ɂ�@��S\/��:
��D|���ٞ��'�!�!Ɨ���7��G�0�,Z*���5��mVr��َN�Ƨ��8'?��p�ޥ*�a�Z�zt����Ǧ��S�`�Sb�������0����&������ �,�K�#8T�'�e�0kq��H)���RV�7Ϙ�Z��*w�D���yk�)a�{,�t�KhpX��\��I�L#(f��H�1H7�P,G� ���\�k�8�	2�i�I��36q)e�݋���)�����{����H�#���g�BC1<̉��r���	��^}.����b8��a�<�W�&	W�S,͗&-i;�EfR(b�O�*�t�������R͕����1��:��sî�ٽ)��](W�~n���\�9��XQw�6Y�+{&2=I�'<N#�uR?�BU������j�G�w��ʀ�ڝ�8�O�Y+.�۶��'�}��hو�b��C�j	���)7�
������!j΁d��U7����1�@L��JJ���l���8@�
A(�8X�+p\�x�
C"����R�mЁ���z>q��O�7�>p��� �޷~�G^h����/�����,�*�?I�<���TdE�NCB�+�2�3W�GX��0-ٌXOh��;���m��o$��`D�6���0;�"�2�|��&�Ź#*���?(;
�	�2�!��c�!5��p���m�d�-(��ƌ���]��Q�y�T@��W��_��DF�dλ�y/��&�q�XK�Es�p�C�+K�A��(�	��Kж��P�&��?o��a�C�Pz������5�)z�! ��M,@��F��ej���G�-P�<0�w*�$8pRX,P���Pm���X���Lc"N�]Y���f�����2�Bb,��Ss"a�;4jn��;���a� *�U4�]��n���"��'��j��)Jc�BdI�!��U��	c���,�$��k�d0� yJ���Ǳ7i-�w(՚�\�Uq��%=��)��D���U��+N<72�1[Vadi��bݨ(s�$��K��������|��E'<�{���]gI���c�@�My/r�Ks��њ�V��Iv�{��7e�V�(��;�>�x��i�Uh��d侈1cU/��]���V�4+\�W�d�C"�e�g��f~?���M8�G�`5�֙�D�G6W�qua$��[c�k�����-�É+R�Y������[ΛH9�������R��^0簙���ǜ�
���%�k�0��V�߆�cY��g�k���)��"?u�YF���"�)Cr��!x��b��oU	?x"!�c��L�������C��ӗ��Vᩈ��/Ї�� �4Tmm����a~���}�F�<�4a~������4�3�����dP4�����5�l9�o�T�/�U0��X�G�Z���Jj���\F��?���0��%ZI*)�l��5�=�C����j	+��N�����`�v��=�&����M��f�gz$B�*��8�0��1�����lr$��
M���)Z�b��fmXuN+p!��&�A��woG��؏��K���8��I��w�/1���$�C�o�����M��&�n�`�K~�'-�͢�5*J�n����o`l��a0^_�n6�}�p��;�$T7��:1{�3�����W	z��}�8:��X��ڲ?��3�lh�>$'��P�f���9�,��qe��i2�=��.g�7��W��ŧb��z��D�NM'�w��xQ9�<(І7���Y Gdz3�)�e]B�Vn �+��5*LX�F�`�d��(�&��P91��'9�>"#�4�4�R��#f��*����JlA����.���������,�*��,Z�W:����08�xȵ�+u6�)��˶V@ܕs���x�����_02 ؾ����w}�N�P�Aݢ��:R��8�Űe�&��`i-�?��:tx�^J�B���l�6��,�ݪM-�i����UY�c�]�:�}^�1_o-7�B" Yr����5V��Mo��w��(��Z��w��rf�to<���Gyz�	I%8}�i�L�ٖ>�rϣ+��g�ʂ��[{�~��7W��%��������7��5(EC*x|��PO�6�㞥̧�R�onP��a�e��c��M�Q�בV6���4Ѐ_�,��pr��h7�#:؈��4��"��|D�&
�ar����5�� �� ,�c|(�R�eH|�?��=���FڅN���_@[\]���"9�P$jY|7�'�8�w�Te
��I�!�+�;x�n�q_M�d��^u�#.��r�����p��}������Ie��} w/ɱsuYp>��ޱaM��w=�	���Ut��љrx��3�+�iQ�\�jJ��VK7���s��g���+�)Nl�^ ���̿�"?;f��'���Ί�n�Sg3r�`zY��ǢP���f��M����n�� ��/��L�R8�_��F��|��[Vi��q��'�~�4�Ҷ{��5?��
�9��,>��Ʒ�٧�2��v?`�;��?n�"l� X.�30�l�Ri���~`Px�9ଫG��F(��~��xI[ y��U���ݾ�u��D���-fQ���}�)p�e���ʬr}���惀N���.5ZغMc;�����|r���@\�k���-G	߲���_�޻7T�#S]� �������-qO9�	-u�s�6��^u���t�zCb~��/^ѽ��)���L�;ū��	�/����$?cւ��c.��USR��ZR��B�#ܼ��n�����lk�ݕ�H�]n"|�\����==���x���� ��8�ڠ)F澀W�]z��M���J�cC
��!`?�BJﮓM�-��	�	��	�8'�
�EͲ�{ //�+���6a�m�����X�1aHq�4�1���$���_l�NI��k�`�K�����\CK���8N�q��b}��yc�>����.�.lV�0���4����4�1��"q�������K}k�ʳy�-�!�#ʮ��]<ezz6"�K�=�S�D��#�Pf� �~�A�t�NF0g���J������RnQ�R�&�yo��P�q�tY�B~ưƐWyN���ԉ�y�ѭ	j�<#�yT�h�P}�Ϩez�7U��١�[�>u����1��~g�'�O7�����c�n����zr�_����	(F#1���#�?���ۙ6k7�֐w^�5-[P4'�L"ʌ����1K	Z��bn��s.!X  �N$�]w2{�V����_L�xW��D�#:X�
�̆O�{x4�}�3	n��/uD^�.�,�$gQⷌ�e��6<���ƃ(tHSq�)Y^�0%qxj�j�d}��8ܲS��A)�������FN[q��La���/�)�G+&Y�EA�� (7f�Q�H��^�J[�nVN`�6�����8�}@�j��˷b(�����,�A������]�_��t����nh&���7`C�(�$�siiBs�>SL��|z�j}]��H�`���}i&���p!�@���;C��(Y���k'�S+�+���J+�U�o�=�Dt�e��/P,:���;�#S���[� &y,�=��k��ؤ����y�?@m��2Xr�L����h�$�r��xʎ�Uz!�hb9�g�FֵT����P�	���d<�7<�3nT̩��4��+3���H� �TɦF���Y��m Ύ��[�0�3QS�)"5ɦE;��.�)��������������B!˔����B����
�q��Z�P�����8}�R3�>�7�*(�N�T�F������xݼR�Y��O�[�w.b��4W�'�bX�}���:l�5��,m-�J	D�\�:��"��`N��_�2��S�N���:�S�j��nݢ5�qs��ˡ"�����o�����D�!F ��r&��n�ײ/��� ��n[\�����C4���v!����ࠇV9�\�7�h�\�~ ڷ3�߹�Q���W��j��^�B8��_F��Ak�������	�1�$ݥ�J��S�b\X��#%^ntb,GC�b��Ct�_zI�1��G�dYs�ކ�}	\�T�#ǥ���b�Um���b=�idiYSD�KQ�{j�9^`ru;�Q����`��2��#�+�F��kOn�_�$�����J}Ο[!G�52F��^WWy���e34�>��\0���WzR�á�H�Sh�,S�1Bu��9AJ{ $�]Ғ#�"��~Έ&��&,��5�-,�s���b�H�SDso����.H���X)슨>�!�L�Ƭ~�s	�ߘu>�F��i|�N&��r[�#l���[�����b��yiJl��7@;�py�
s1(�gf��+	#-�b0ʠ��|���=��P�y
E�'R_ޙ�K���t��]���}��Q"/"�)k���*~>e�S�9[�(B�7A�\�yl���r��BbĤҝAk�$��蔵w����G�y����,q0���
����%�x ��&�¸��+#�TtZ��;��9{z{(�]|�x����6��v*�x��J�+"2uQ�f5��.ʆx�N�2=�k���p�eV=�#��Mo\ �J&�!��В�k\��
2��J�Vᅽz���Ҿk�ͥo���*�L%���0�Y�2��:���4���`�� (f��%�-��g�V�������S�+1�������$@�����k޽�v3IRM�*��?2���4;��m� $0����	!�sC��Q�������w&���_?�2�/|m��(�齪�����]~����P"�Ҍ, o�Q�G��.z�?D	᭔�|�añʾA�(�W�0�u��j�{zW}���_8���R��3 �%�#��]b=���͉p�d�W�G�~���FӦ_��ə���&���)��Еƴ��?M��޺<X} 6�JkN�R,k���fLSOy�����|m�)Bڎ��V�w�;��m
�F