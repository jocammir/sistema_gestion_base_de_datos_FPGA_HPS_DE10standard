��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��Nڭ�	�����B�#Z���?�4�j��0�ΐz�A�y�[��I4�fB���_Ɛ���-����B���M'~��k,���'zf���]A�� -̭���ҧ���D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0�����0)v��H=u�.�Ƙϟ�WyM��Ә=�E����~��H�fF���1�5Q&hY�x��?d&:������"��m|Q䵱
i�m��%!/��L�9� 0�>�ɴ�&4~��H]* �ګ�V.�%Q�_8��Ү��t����5��jiI���eI�%2�q-kL8:����H���2P�+M#�̈�����҃�2�P]�b��1��F����9R���{�-�ǲ������*��[3~���W�D�B�$}�t�B��s-]Q���O�D{���5�r��$2g=M��R�M��
�Q��dc�$N�C�r�i' Z���$�g��[����C7��^�1�v�W,�=e�E��Y{s�pѬIś>+��	����Gu���� �����|��K�{��h�̀���c�Btٕ���z4TYh}v��4e����*�]��c��;��8�g�?@Z�Є7K��|Bl7�ֱB�����7Ɇ���%���q{Z,�c��dPN�<��԰h�͡Q�,�%m�,+���F�?��#��.�r��Pjkg/:4����6O����h2����=��x�@�c�IBT��8��Y5�n޵��Fů�Ѕ��x��,�z�륰�^x?��W/!O{-��_��̔�ڵ���B1�:�����|�@�� ��E��9A=�n�ㄦ�������w�3����߲K�(�܈�e����0;��lyɆ��Ǻ_��<��������A����oAc��gy�"~ݣM$;0*�����6m�o�~��eg�S�K^pѮ��KM9�����K��'��>Y��s6���J�h���P����k��3~?����3Q���Ȟ	�PA�c��n��M[p�k�P��ǧ�	\��y��T���z�yH1���LP���F"m1���Sm��蔪m�qթ~��9N���*b7]D�e�e�����!���`?�I��DK�x�O��\��6����mFS�����T�x�S���N}�S�â���A*M���7���1C�z!(��i����Hj�xY�5^��Ґ���a�%Y�*���M<��o ��i#r6L)+�I�ཹ��9�6�6�#:ˀ˱C����M%��<i�+$�H}�_/��	1�n.��rRK_���9��yi�B[�Tu���G�6�����"�H� ��:	u�85N6�ۋ� �O,�AВ9焽��rkd��i�}�#����YZ��_R�~��H���M.E�	���bsL�#�J��m����s_6I���@dEQ�B4�
N��?�.c���X�v/��y��\� ������w?\�d�Y��
��]~�H8� ^"oc��o��
�x>�"JG����Q����Z"�nG�Ik�_K珜Bq��-���љRA��K�W8�}�}�{�^��Xxĺ@<��Z$-gM��_��M>VL�-��:�!�A|0�7�3X&��p�x!��n���D!����?�(���vM;��X:��7���פ��m��)^��ôRv�gI�����C r��&�:���'RJ#ц5 ���|<#���%�����R2��dLdhS?B�8�����;��cD�;n�ޥ����9V���q�1�U6P��'��=��t-U�t��Q'z?j�"6�����1!/��b��y���>i�d���Kpr|�t�oa����������ԥ�E+�4$�q�my��
���4)��O<%���̊f3��Y�%��8m@@�5�1X��tJ��>m��S�*:ci_}�UMe�s��A���<߆<X~Xb��D���7h�)\`�����]E�����[l��T�xʬޙ�y�h���d�z"�U��;��h��?�m _o���,rD���!��'���կP'�����ؽ�r���ʛ��M��8��KP�u|�_ف6S�p�9���.�7>+A=�@��I��2��^�"��oA ���pf�Z��
s����I�Sk^��d8�1m����$�u�����	V7�4�u����2��B�-9�|��E�,5����rbؕ�˪	ĸ�}����)��� zti.���ʏ��n��
��R��~���y�ޠ��cV4�7�8M)u����*dߪ��Q kY��^c�0�� l8�������K�	<V3�%cL�D�w#H25�9=�2�AZ�9�RI��!�T��c����MTg_[ oA��O�v���o�E�V2+��39�T �[:�c�o��e_h�=.�Fohԋ0i�3W�����l.cA�I#�o��\��j�5j�0���@>+Ϲ��`&��r����	D�\����GAK�L�v��O�҃!jL�=O]jvל������t��9�YA�*ھ͹+�h��j/}�Ur���Ow�*�vSyC�H���ZAw�Lh�E����f�4��Dg?�F*����XN��G��!H���-���.@��,��H��L��s;�Fp�P����X���n�Z5��v/.W��o��zy��}��ڵ���*�.���v�wg[��[�\�� ׏�V%�o'\��V�Հ��	cX�7P1'�;(�1�� �[�D�p����Y?�r�!��I��=�$���t;�}0�G0s�E��P�d������sN���q#��E��>�F�[�W�7�Z�R*Fq.:c��!Kf��V�ʂ���7k&�E���v,#�HS+r��*/!n�ȏ>Y�BpO�Hǫ�zPӡ������
�3%����!�RHKpv7�=2�2�jFp�oG�2:�bi b����������%w)j�E��u�ъ;�(���s[�В Ԙ����Q��
+q����
{=�~1�cǳ)�@� ��uΠ�γ�ٯ�i��FS���oIt`d3���R�5����;�=Q�?��4���~5���Y2�\~Ij��=O�ڀM�.�d�e��}eIXB)>It(<z3����QB�"%y�R`�,�>eZ���`��6"���)�ұ��E�_t�ՍȎ�״	?��;00=�E)�P�����x�.��8�����$���(�?���9�4�Z�[��=�;k���� ���R�5\5%[&���@�m�#]py�Z:��i�aH,�,[WXt ���m�B��*]c
�ݍ��S#�P>��0�2�g(}�~)~3�|�1J2l���c.�*F��L�TopP�:eS@5<1m��H3u�2Zk�- }�O
`O�p�Ջ �-�:u��7����&`s��p�I_�!��̞�g�l �9�&��u����RlBR	��!N6�]��R�E������O|�2�;�n�[j��/`����0]����p=qZ�R����Vh�g�'rm�s3����y�B�)񑊤��U�n[��5�=�V༁��#���/���[^�~�cń��Y�څ��T�i��J��%&��tŲ�"����=��;�nA���՞wC�A�����S�F���0��óW�Z8Pϛ����<�˔R�{]���JyDa	��-���s_��O(j(eɒL(DдjB;
:�]�����#��w:���b4ߊ�2���F��ԧ/x��)�W���u6*f�����Me�N�UP���1��=����N��X�!��Q�>��G��N�WqB�1�2|����2nտnQ�0ܖ�{�FC��7�og�C0tܦ�z����h��V�J�-�6&<��hGÃ�t(��\V�5� ,k��<�u��t��
?�?O�B��jU9v;���5I3!x�N��Ů]pݚ��B�@��߆'�f��L���l���
3+gN�=�k��
:�!�Z�Ho"�r��h�L���n�J��Nd�P-H�
�N����@�Ss=e��uJ�	n���·��ذB�CL��*f�W�Y�wdp�	��p��,\�6�h�M� 7�V�B�
����~��d��D?�&��"�nD��P�mq��_����M3�I���1w��*�7S9�b�g�� ���!0��6�s��7gbc�6�H��G+�ї�~��c�DX���)��O|�+����`�ۨ��f�2����:�3��8��.�/�K�r*m��l���
)G�H��� �g��.E�)^N�T{HԎ.��0w8���`ӹ�S�q��>�؀��Hɇ���}�N�;�
R�V���#��>?�#*��SA�6bS��7��M����)�߰���� '�@��}�8�/'������N6��M�c�=@�g���V��+.�y5���7��ѕ	�J*�;���c�G���**�fm9�g���^��]@2����B|w��z]�|�-S���L�Z�z���S��6k������ɨj�P�t.�L5ᄆ�;��o��*v��\��ABO<a)�K#V���_C�3:�,q����|��MW��
��Q���aJ_! �p(�x��2�
���V�{eQ��hM���/�>� ����c���������r��������
���<��#:,<���ڲ�:�ᖈ��"�vk��\�Z�q\B�t���vS�>�b��J�U���$|0��s��K&	MbD"�[��m���p$��k����HxD�ԛ)�N}Y�2��y�)r?�6�Q�4D�$�8��*�Qv~;��W�S��A��A�,��O�?�Mؒd$��s��p�HjE��ލ��i��֩j����*�����PO�.��s��9:Ibrǆ�X��E��&�5RȄ�:���NϨ��S�Ը��;ȑW�{���q�`a/t�u��]���=��dK��wIx;?4B�>5l  N�����v��3��00sR����C�����I-��� �`�yUl!��!>��ۄ�hD��oT�&n뚓8�)�6�Qnqܩ�Fq�;�00É ˝p>i��L�!ޛ}�R���~��(-�Ɛ�u-��/��(Y�fW��@Dn�)��õ	^¾q�5�U�N,�p��J���e�e-zE��/]IK�\�6�!�-��H��(_�G�쓻XD�� �&��%�����w�f�3,���ԋ����J�,3KU��}{�p�^��H�@�$���~��Db	8�}��
=�z3l�ݜ����Xv���(��B=����L���N�[}��uJ�ʍ���w�l�\��Y��G��4��7Df�!SRI�ND̟��[�ZU6�o���V�_ !w��"Q� ��^{ihk�9q����s{�����;	��W0s��w@�9y�휮\[#%3ɞI�w�bW��4į�n_��[i�a�6�VX�/ET�u�^�K��n��*����t�S�|��y����`�t�ѫß�v�\x�=^��1|X�V`����GH�{�!�n$���"z��?�a,�}��<�c����<aý��7A���É�6�J/�@PT��<�D|x�P��E����.P�Rߪ�%���B��6
$M�Q�������rycX�|me�/@ �ȓ:FYa��q"�M���N>O�voڋ����Vx�
ńF�P��mo��*dDg�t5n��%ɴ��9�3����kj�3%X��[x��/��8-(0a|�r��`����Iu��&�V} �<��+�B�­$�L���y��0�d�~��<��Ō�-����9��et�H���P�F�mkz������0�r+�.t��N���j�n��	/V����+���j_���Z{{�����Y���;x�k�)�	p'}%�CkÉx��.�T,���9L\RՒ�H��#��}��\Z鴼�u�W�z�����0ʝl�K�����j&뽈t����郩9�t�5W�_�/އ���D/Wí���$���2�V<:7�V�u�拿�Ȗe��C(f��	�k�T�;#�iC����n�r]��UA��Gvk���H����(�,��Q+�я?��x��<6�$�D��A{۹$�&B���[��
���ۀZf=I��$5$�c57���(w���]�A�M_�W�=D�!{�o����;]����u��|FG���#N�h�
��)1�w@�S�������l�%�)�e�r}$����ǭlZ՘������ۻ�O�q?K�����7�6�r����2��I ��#�z�B�d%I��z��q̇i��I�/Е]����e��Ӂ�O������U�.y5j{*����"un2�y���m��҇q�xUp���c�g\^� {��ΒH��-��D��,���l��2�n�O1E_e�%��J'PQ[��+5��JC�����Q�m�wF��6��������B�X$z'�}hߌ4&t���%T[C�G�Z���{?��v�g��xG],�IJU�Z�I���cJ���B��
���	��~W��D������#�g�h�T�����yt‗��1$��]����s��T����j(���R���R�&%:�]h*6j�Sr8���� �be�W�*�&�L��Ք�~���@q���-��̺zm�lpN��u�"-���!U���Q߄�=(��C�C��E'�u�o��FbY G����ͯ�*A�F���.�9�QD�)�����k���D��|9F���PހG�#�E�z.���L	Ke�y~�p�s٫�����Ss��i�U��'W�yC_e�ѣ�n��B�҄
7��b�s�c3�����$�jk�t���GK���!
�#�c]��)x�'W]F��I���h�i�C阱��'��Pq9H�n"R�:\���=V�����b_�����=J� x�+�K��ă�]逋τ�`��؁ޣz/�\^Dg�����]�Ǽt(M ɵk�橁�s��8>o�/��E$��]M���MZ�4��i
U��Aג�?��x��ن���5�P 7�&4��L�N����^�W�|+���R�E����A�F��X$C�����CQ�ͼ��(�ߩg@�FQ��I3:��N���ܙ��5�8��S�.X5�C����Jl���F��'�ogO���D��r����1l��ݖ���pp�@S"�_�f�9���� O��u�ڰ�xy/_���
�����G��"�)*��]֠�rg'�����o��Ū�:�x��)j}���B��#?��?Հ��ǌ�5P��%w���$sqoZ�a�BѦ�&_`�_	�%k�z��"���/˂ܟ��=G$8J4�Z?��B��k�ZҎG6�(��>�y;d�5_�%f`Í���y��>�|�ی�Y~�F���(�1��Ѥɬ:\��v��䡉�H��(l`�����9ZvC��"A��#?S������0�7VU�
*�M��y>�N�q@�}\=�'�_����~ѕ���;��%���4A�J�u�ĉ6�gj����m?��6J'6�����N*%E�p�}�&)R,�f�Ì���k�7ᚣV��p�v�c)��-�WuES��ysxŠ�b�E�ɼq���ZBơ�u��K���6{ՔOPٔ�Z�t�{+��
��1������R;J�5�:G��N6�q���w�8�0��x�;f"GR��[�[.�n��J�Sm��n�s�n��)���Lq}�x�h���Cy��m2���Jލ�ɢ-��E��S!������0|����pt1�^���eS���T�-�M�g�!�{T�ޑ�a�9J�ӜY*�Z��M�;R�Z��>pi�֪q=�������ǘ˯��R���TXR���IA�C�����#��FY�PβC��'�X-�4'[��bY�z��j(|
�U�����eQ-�uv�Sfﾈd}Y���:�BI�z?s� h:�[hU���$r������	p;(�fk֩bS]NQ�S��ʌ�H0� чnn�?K�L尔�����QԎ�#�o�'�hɸ@WBJ�%����/�OW/T���9^�dܰ$�L�٠�|og-P-S@�Φ(��;!j��Ƨ�^��]�"�	Vq���#Qe�����5�l%��.t�8t+��%�l����S�g���Ɨ��+En�P�/��[���嵱vJЎR~.Ys���l�m4k�?Oހ睲1�\�Ԩ��g8~��t��3�7ȏ�v�����vS��O�aڜ�z��)�l�Y
$[M�z����\rT�S���\M�����C��\L���:�� !�0�=������Y�4!��WJ�d�����X��t.��h:��p���G����&K�p��s�^��O��\��X���Լ���j,拝]7���R!�2P 5+^z�q
V��ܞ��E�ʞ��v��h�H<m�YB�#�h����tp՚΀Ī�{�8�R]�s�Td��Q�K��䑳j'.'ܾ	�y��[�O�j����yh�6vL�j�	V�Ap|�;��zj���c�^���m��O�AkZi���H4f��~j@���h<y�6K���A�ԗ�Q����|��L���N����{�0䟍[������ҫ�-���ic�|5.*����7����b�/h���$z���;x/�@x��K#&\��G�f��7�l�i�B�ZXlg��3)������z��� ��3r��f�6���1�>흇?N����v9UVw�n��w�d@�����I������(L8n���Ҕ��u�U�~p,z�.w>�Z5���_l'בU�f�U��3��Ţ[̐♎w�E?���?�����M7lGP.�jK�ifK; �5��#Y���D{C~�0�ۚe6���Y�X$�;3���dc~��x�l�~���sIX�7�,b1�������cT����]젎A͸�a�Gl}��$N-'���[K1�B>�(Z�}���?�r�6��7
A*��Q}��XٱLNk�.L�5�������ӈs2]<�
=0��!5,�_љ�(�ߑ������{�ͯ��f��F���>K	�҈E�<v��q�'֒�/����e��IGb�ƭuM��c=0|�����,e};3�c}钠���T��$ew���_�Yl%]�%�D�4*�N�}sZ�5��LZK2�EK
�F���&0������iF��w��)�î�hr:�US��>I���,�Xx�蔏��~�5v�ѩVDh��sR�7ˆ����7,@��F��ú�H���4J�rM���
��ē��ܞ=i�Vx;�5����j����9߿_��Mؙ�
�	6��e#��}9�z�˄Ź� ��o��+n�]]n��/����ʈu6hn�y�'�Rq��
1J5���k\�f�%�sI#`?ǝ�,�c���m�b٥騃��0拫�3�%VWl^��Ⳮ+tߌ��H~H���~ޠH^$��(�b��"-'ק,g{����C��&�MwE}��t��w�Ȫ:t���i��eh��������X���@���C��Z������L[*�3��ߝd����.�"�}X�&��������f�ߣ�wƧM>>���e�~{l�ߊ�f��!.��/ �ΫGk~��m+����S��ܗ���m�X@t��i��2����t<�22�y��Ӿ4r�h����l�#��]cU�(uD�W_q;�"سVy��-1��P����2~�:¡��<� �qK���^Y�dڱ�H.z��T�E��τy�YE�Թ����ձgͯ���������<�=��
�Jٳ��)Q'F9��N�d���g�
���^��Pw�"�����>�UV�����\t�1X'�S��ҡ�S�r���QFw�-�~�Ip_��Cl����m_˜�������
)��T��Z˖��^]�ղo�mk��g������0og`�[$M䓭0��Cxm��!&���RTQ�Er	�Ua�=G���8��!��X�N�aJz�����"4�_�T�OUP�����F�2�p�[EMY�tV�P��x�qsxU��e"�r&A%ސ�Sz��gݼ@���|z��!R�L�?�����&q��wӯ�Vdc��{�!K�T���6��y�F�@�A�/�ؤ#C��z�+�vf���B����lY�\QD�>�������*�x�/F���?ו)؂߲����G��G|i��)A�>"���vR�߰�n���ɽ�s�%�Ə�_���f�O�[1����^ws7(v��;jO���y#J�ɠZ���)��W��6�R��˄�*��c�� �Mq^Qm�a�p|V��䠤n��nx ��ES�"i��5��@�9�a�h;!�$ҙE��6�G����W��p�MM�y����W4��xM�s��N��fౕ~&��p�j�+�X�+@pp�@�;��td�Kt����q^�ܼ��Z�jP��}zĮ{6���Ҁ��=�O���ގK�A�Jo�"^FN�����J6�g�h�A���Z` <-�u�|�G���$S�p��3E؁�Y��x���rI7��4���W�z���!�b�3�}p��Bi�p|!pS ܑZL�r�aC6:�����M�u�,�5�}x���O�/�m|��D��Y�D��?�X
,�	�GER�R7��mk�p��t�H��V�9b5�U�N�������1�� ȶ7 �i@�������׿���2R��(*.N���$�꾇TL�!��b)���%�Mb80D��
�OL�D@���� �g7��6�a�]0s�3?��)�\��llƼu�@���RMè\>���$���c��TxQH�"o����­YG0����Gl59мf�����3ԑ�%��uص/�2˼�Ro|�~�w�R�N�/y�h��RCэ���̑��U>��&N��>���U}T6M��b>�ۅFB{�u'$SqT��D�V�]H�Ԥ�vL���C�c7�)cfҞ��V:�^w 5k�*�l[�Z������+S_��fw%���{��1c�����9���1�|�;x�t�$��D*��j u�i�,���"銝I)�d�5
;jP�7t?�=0��Pr.�e\�[�rh���$J�%���
��1@[s���E�t���6
���ܭ�|��th�7�ye���#-�A��ʡM�_v�?��o(���?n
N�WY�eu!��@��-s9Ҝx��������k懀�)	�u���eó�����9�����&��V��mi%A9	�0���0���A[uK^X��ŔPS!/@��v>7��>\2���M�3?	�LG��s���swe���a	�ƳM)Ӧ$˘:^��t��dH��9�����!�1�SN���t"D�B�Ǐ�ӲY0�D
ـ�H	~n�+*�h;�۩\�W�Z��(�*�A��弐�`���n��|����}�l���u�T|��b�`J�f����=�E̲a#�_j�zy��	"�� hPD�>���o7������6Hb�'b���;�CQ8��E� �P�������$�ޜV���h�����&
OUy�Y�5�h]Q����A��#1a{�R��>��CxzkD�H���<�M=��0kpm����`���l��3Wăa�	�ހc�1s�D�.Qa)IaD`m�lJJ�!$R&�%���I'�2w6�i��a|,3�t!����T%��e�8�x�J����������lf`:������d�L�O�Y1��s�0i��hݣ�N�<�����)Th�Sx�=4Z��be��NOv�d��M�:� }uE�~�>�������	*���f����۾�źlo�i�g3�߁V6ϟY�fT*쌓y`#"|`fc��ޗ��zG@��	�I.��y
M-J�k���������BSꪔ��f�B��c*���\��T�K��jG�{:��6u3xf�"a�֛c)�"��;8d��'q,+���?���n��Hj�3�:����'�`Tٝ�B~Ӷ�&:D��+ɸ��3�w��q������?���(�˕K���a,k/�!�|vՒ]��O�1���
�7\���7چ��qmn�qݚ-Iy�B�՝�>��gS͹�dV�O���f��qk�Qש�� ���~,��Fh永G���p2,:��!��vs��+Lc���8RP �@���i޹g^K��l��`��EQ��Z�[�A���cK��=��
%�slkl�
vB�ޗOn�|aţ����+�f�����d�R�@�;U/�������ʊTd�j�x3L���8@;�Ū}�>@mE��&�iu�V�$mOX�4�a@_w~A���,u�F��+��9hs�����Ͷ�޵ �r?9�-%k����9&,v�rS|����IU��u-|����_^+y���0V�B���:�u���F�7+�*��J~@�(��:�J��y�]�ڸ��1Ȯ�"<����C_�6��`�p�j�C�q�:^G��ĵc�nw�@ui�g�V�
g)�yWSJ�p��a��@�4�{��n(��P
�*-J�Q(?�g����{���ʚ��`+#d�nR�$Mg{w���&Ϣ��&�5����3R�,����?Lw�v���@��5�K���Lh��0Rvo�M�����!��Y&}S KDEHR�¥VN�%EB��4�5�B�0,�v��-�睫E�0�/��\����B�|�X��"2`h��,��.���k"6�S��4�s�]��xt�R�J2����|������F!E_��2cCbBx+��' $��N�J\]��(*��oa֢z$t2A�=�l�52	c�*�E�#�q�-�����;]ݛ �Ih�M �|6_��S�/����RN1D�����C8�U��g|f����ǫPpx�fۍZ�
��Y}��h��τ�is0U�-}����g�[������Te&a�U��V=���) =u0%�#[*��
ߪ�x�׫r�%����q�*#��/�'O��bG��R]-iC��x�/@������M�b_�\�B�I4�d̕VӢ�_�����v�c�����uo�����V�y����p�_g<���.x�Y7p��~���,�_�m��"I��w߃�	XϹ'��8�d1b�����MK��\ڗ&;8�8ß�t�s���e X���[�ˀ9�Wk?�(�v�)�E�u��	�gFٹW��g^������y3�.�� ����lU�ԁ��0Y��̕-GJ�܃s��[P����3�=I�jz�B��ҁ�QR�'w�����<�,?��NY\ޤ�R�.���a}`�PS{M�����=O,�ד�2��tB23&�5����r�Mjnu~?��%)t��+�ǂ��
{��]�8���o��-%���Jqդs�-ۯU��T��At�q|��4�;#�.�:!��1�D.e�6,��=◓\����M4���xW�}T�����wt�%(8���DN`[�J��U��Fr#e�=�P�T�K��`��H�(�.5�� ?gK,(l"���+{���(�3�,>l��NO�j��n{ n�o��i�����cS��9wgk)'~�Ys8��"�e8Hᐊx�N�"�
��AN,�o/v�Ly��m��y���6��Tiu�$����m��/�o��t0�HF�+ӫX�9~�����&�D ۬��Lf��G�_�5y��GJS�b �=�~[��Z��ha���ːR�ϰ�@g�
q��w��(D�+e>��X��K�S��lR�0����r�_d�S��AL���+2������{P��!X����y�\�D�%%�g�ե~���M��+'��Քh�W�w��eU1�@y%��-y�k��1��a��d�Vm_ƣһ�&e12N4}ɮH�b�\+rbi`��Au^�/%%���7�����l�6�U0���"�?BYA2#T�&E�c*���`��
�[���<�	�����f%�"'�.o����@&���ǝ�O��x�S�/��SyhG]�vy�H��?��>�pP���`t��yk�	�O���x���Vܭ�(�#j�0��D�(�h����s	F�����mRe {���0c1�bF{kA�S�Md�<�����E�����/��Llc��WC�K�Q�ÆA�iX��n��O�1V*ĉS�����u���Y	�tS������
�_d�d3�vD��� ����;��]�a��Y�~Ahp�(��~`��8'�&LQG��g�0Յ�4� J�l̿���\�E/�S�}51��{W�2 ����a��5Jp�)���H	�!~��qm�#��;hZ���';�)�%A�'��=nR�>�v�B��ˀ����X��3�B���.� �������_�R燦R��͔"r5.|�_�L�����g'_f�X�$ɭK�}���zGࡏ0��x�&N����'�	s�,$��V�݆@�%N��@�;虖k��u?X�3�/�=F�o��v�.��>O'MG5|���@ó@J�Um���Hw��&J��ZW���+S�"_S7�90�K�*�&#۰������W�O��P�sI����d��\C�z�/.fv}��G�L��� )΋%l�ɭ�.l�2����-���S6���^k��e�;����?T��av+߻����{��l�6)� ��c�~�K,Gh=;�\�$�W���;�^�\�|ݳh��p��k]����6�x�;,�}��|:C`"���~��y�O��$���j�x�� �����O�%
T�Q�[���=Z�+�a������l�����A��宒�~�*��0��g��9�� ��us�S�q��9�K5U��:B�<��Z>������xs֤�$�Z�Au�:
X���z��D{��]]mL��7��ƴ�b���������չ��J��!Dg�MK*��e�,�*�tY,�;�l�Iw�/�7j�=/��R=�۫�S�"C��oo4��)bH����?m֐��~��R����d�%� ����Z����V[x�v{|N<����(��p;��C���� �L�g�)y@�?�+��p�j~j`�S�y�#��O�P('�6��p�#�UTR{�v�� ��k2<�p��,��R9��i�}x��k�%#"I���χS���ͧ]4}�MLş���i���=_��8v5���@>�gD���df<k(y7�~�P3�z���J�.d^:�Y���$�]$9c�V�Ѐk�s�gZ���a��p�@!�h����1�� ����sy����_�!��L���8b<����rv�xx�5�Y��'��&Wqr��=H=U �T�N,gL0h@V�r���9Z�Sc����h�b�l��x=�?��A.%�q��l?,��d���g���xQ�=�k���<�).�¸��X���;Fܘ����=���K岯���Y�N>�E��ʞ��cP��9_j����Hs��iK�B)񇤿s�����YR9sn뉙�A5���T],����:��[+E5R(��=t-�pd4&�M=� b���F�u&�n~z7�h;�w>�f�)ŷ����65��xIw�'�t�|�'h�[�+��S�"�����:m����oH�s2������p}h�!擸g�V�W��㱪��L|D��o�d\{�#�X�ȅ7�������A�I���г��|Ɓ�Ub��t۹�D���mf�g#G���`����@�a�i�Qs�]����PVi)���6$�ႈ��=�������,s�&�*�JX�Im���O9C`q����I�<D�6��B��)Nݩ��z �pr�s�}��B��7vh-��}�\�HXu�P�;.�o�eq�Å�a����T8��L��-�~�]�{�'&�z���8�Q�*Pޕ�������"��Β��T.$���C�7��.Vҭ<���)\�X�x�yN`�(����r�1�Q���U��ؤ�����.N�Oa&��U5�j�E%ɥ?�Pd7�d�E����O�i�s�_T�4�I2���E�y`5LHT6��#}�d����n-P�Z��nX�F�E�u	�	\��%����	 c���IPŌ���yq<��7Z
�7h�~]�{�vӜZ���9a��մ���'�������hp(�?U�;���|J�p61���SHq+2��䊣�Uɻ��:*��	T��ʒ�hST��/��[)�ډf���h-��[%l�u�$s�#H��!�h6��B�M��"_ё��t�7�S/�"E�T�ߚl�D� ���8t�����U)�.wJ<���ا��
&{`Q��K��^D�\��S�Ԯ��5u�(B)h晅�_�uz��z�,�Ev�=������&"Udq$ڔ��ҟ���X�V�ݴ+�$KHm�YA�����bY(�>�D.�Qf^b��dgUl@��s�-f؃"�Q[j?
�lxY�>Jl[�cJ����\�1d��ǖ��])O�C(�X��7w2Cp�-��:�^SӁyQ�k���2��7�6֜��KQ�jE׃�n��^��zY�t�+�y���_y�L��ybz>���Î����X;���<�D��#���s�H�����2��Hi����y�8�G��k���G��eg����|Q�xY6�c����q�g9��E���D6W�i���Bس%l��%��mHz�V��`U�x��Ǿ���L&a��aj;��s�(������:�>"+U+�"^���#��2:+^ٞ��LkK���mF#����X�@26��I;!����Q��l�����$����d��V��`�F�3�d
���_��A�i�R��qg��nu3��VV*��9����POMﾃ��E?�+�.*�쇰1g^4ț�����0�S�v.V��#;�cWմ2NC������sÿ8�f���VYO�}��p��v��&8C�G"BCy1~��,c��ޞ����
[X�0	�Z���?_��������g��]�Ο��{��d���3��[���
O0��$����!�)}��e���_�a`��N��Q��ͤ���e7�w�ֵ��)p�-�'dBX}��&_�V��O,�W̶���U;*%	j�H��p�Q8�}�κW�^s6�
��k��g�-���kW靶��ª-P��&��!�~Y�y�
̸o��xc�l��i�F�"m	1�u�Q�i�9�LJ�<Y�h�܃, v��û�"��g���z��;��6�s	{XU
w�(p5����N��@�2S����"J
!��5	�KOJ���q���ydk3�س*h���G�:`���ۘ�Tf��7)����G�XJ�5щ`U&įZ�GL��4��ׂ��$ʵ�#��8����%�ᷴ��v�l�el�hN���bUЎ�N�Ӗ�&L�v$�(^����#e��*�nN��i�����ё��y��K��{aMu���Ɉ���0s#���˾7b����K>�1��űi:9��]Նw9�C��S�ͅ-�zs���Z��Lq����ˠ4$�[��6k����G[����Òa�x?*���,�����r����G�Z�xO͏NW��>���;��y�ŀ.���2�,-)���� ţ;%���T�&!�I���n? ��/3`vgu>-�.lY�|b/z�s
��$/���'J�5(u'#�4"���a�L�f���i�MfDJ�F�+����
��[trrQ<d�,ev����Ȱ~�T�`��:c;�[9�!���\�co�i�WiPzΰ���ct33�x�c쵢��R�t� .�m	�ϮF�0,�k����h&n+GckҫEU�!���bLe����2��|/m�Е���q,-�x�������)�Ho��P�y4�n��t���3�avLM,{��s �3Dwi8�yV���F��W�2�*�=�<i`����*8��Ǣ�i?2c���
��}�T���Yj���l;J��]��ÅUj�}��y��g)b�x�ڲ�W�8� ���f��A����Is�9c$��v���}n��Rt^dhU�` �w�i�I���F���Y��|�ٖA��[j��Ș������<�:������+�Å�螬V�a�n~A4���B(-��)��X?���y�0���]�|��]td��
�0�����,�؛�C��h��N��K��";��1�Ħ���l�"���ޏ����!�sC�璁��K3���}���r\��i�~��"*\�����遇�r"
�]g���R_�NQ.���R�}���ʞܒ)5{������%I
p=k.�ej�����5�pf��^��ﯗ
��ͻ�K��(��5�xg-�ҝ�r��V"���e�M�UPBT ��UI�� ���>��3+g��B�$I���!�a�1�?�8����A����Π�������H���	 NFI�NvJ#������TI�$Sw���I���/���z�к�{,����[|��Pv��t���D���:	|�38Ӫc��wB\$�hHp�|�ӻB����?��S@�p���aqk���Y	�J$J���|�̞dNM���G��h���o������'w��b�g<M�T4wRcRȉxM3�sai�Q�5J�w<0FE��O�S��7����Qg3]_K��I[Mr�So{. ���#���#.Ǣ�֮��%�"0+.�@a�Q�m證�ɳ�h�dǄ�1�I�6A�����q�gQ�8���ޅ�n�@��¯0�9��3ǖ�u+hK��..��8[Kl�Q�_��T��]�d��و	��Bk����7�;41�s!e���˱���ź�--Q�)��5�S`�Lj�h��v�P� �A.T!��Ј�s��Vc�c*9J⁪G�����a���m��lߑ�u!�� P$���~���E�'2OM�z#e:^��і?�ŞR�{e<����ق�;�t������)��X!�?�ur��3��A/�r�Kߏ�չ���ܲ�Y륯b���}a`jI ��H�e%�����n�4��T��lq�g�p(-ǡ�%�Mz:���n-G�A������Rh~�`ʡ����� ����ل��M��Pe��so	��!�]�<����OZ,��>��TI�LZ9_L�)�}��0A�"X??�-u�(�B��IV����\�.�PR/���6F&L��yӋ�9��ܩ
��gg=
�ũ(��Y�\�����爞��p[�"�=��&y��EqtsHGw}V�(�,�PR
��譲T�A���h���PD��i���[r���1�YE@�Փr���_�5���Z�nC������T\�"=p=���_cnwM���p�
Ǎ�R��v�C
cah��h��F �e o�2W._K/O��,[$�"����6IW��95t�� ��|uݍ��kc��-}��߁�g%�>n�i�.� �lc�5Ƿe���8�(�9�NB�� ��ix�=��F��y
 ��Y���u�4N��Z}[I Z.\oeA.F+	V*����2�a9G��*��ϑd���*����է���Nz�	y|��b�BdǞ���JX2WU�q�� h�/�V��	)0O̙���K�^�Q�j�[
a�:.Z�Hd��椡rȦ��r���"xEG���b�v��_�P���>v�b`8S�5��I���(l�f���^���*M�늎�/=t���k����w�C��T�b:�2̜'C�����#�V�!���Bٙa[8F��]��m!/ CY�(�S(��� ľ;u������L��{Fۣ�:���^g9>򚾸�8���bQY�=�\�T�U�;B��� �`6��w�;��a�n4�fd�c�0EG�z�ϲş�Tb8OC�k��F�Y���2��p��GeG����&B�(Z��n��"(�$���7�����A�� �
����¨�N~d�x�Fg�d�Ao��E�Qf�������M<#�T�/Xc����l����������d�O�|)T�H^	hN~�h��F9	&�G3��Ǐ��("���蜁%o6C"�8���e��u�6%���Њ�YN��sH ؊p-'
��k\���+����H�i��ޖ�#z�'ً��"�Rd�l�Wk�6�d���M��O��W��h��@���ҡ�V�c����ߑfLI�.�������WJK<�>S�"�����l�򥚭��+	�E��/�Jy�f����{?m#�A�_�B�@}����c�����.4�����R&����&]����(���_F7-bO⡶���Ef�d��r|Ixtfw!�$�A������]�0�X�zõ�,ތ�Vt�1 �����x����h�?fE�f�C�4��*�5/�2Ti���nͻ��r�HhK���x�
��?�"�7���$C�<4�;Z�Q��a�&��:�(�>Q����<.u��~ZIH0��+��T;��F٢NoK:	�r��?
�C�؉��Z[g�R���"	�%!d�i���g�Mmc3���~g���L�03�����;F�_��Er�bmF�^c��R�%qЍo���/(�������E2D��%��D|�^jga!�y����3@{��X(9D�<��RI�uυL�?�L���V�Gj��"����|oy		�(�8�-���>��9Y�ÕO�x���r�љ/�7dO���$PY�:�ܣ�\�p*q�;k���(�,����&,�J�H�8"�{t!����a����<&VI�v{+8!\���� Wc�>t]�f�=�4G��W�h�S'�.��)�id���ђ��IW�w ����ۡ��/�E�H*�6IQcd���7�
����?4�jV����,�����([�������ym����>oL{����?����)�.\��+�bj~@(��($N�g(5^�QȻ7�־^��$� n7����H*
n�h��h"[ê�.�;F�+��!,e�W ��B�$�ڻ�2F�2`����͖�{	���#��s?0:�II��yQdc�e��#&����	8��N��2�ڗ���~�O��1XA�QA}<� '������V�
��J��Կ5�,�͐�������L�5��j(��;S�{1E�� â�}�sA�%h !^���9i�RѴ����U�U�9�3�����ɭ4�#�L�P��N�A�8%�O\{\�	!X���\�nm�8~�v(ޑ ��ʡ�*�Xm v	��� �	�6��������a|���V*]n��:O�ᮊ�9�"^�� �9��(Pý@�
���xnxd{�7.R~V"׼�h����-�p�'�rϜ��/�a��*��t0��^J�C9�m]Z�U"�����L-Y�����[Enr�}K��X�Rd�r�riu�S�kfRv]q�.���D��؄��m��d�D�b�[V�=l�d� ���4Wd�Ϋ��T����;��X�*�z"}�s9��i��͋��QnYw�@�JO����!��N�y�߯�K�&m���\���]1*�)��yt翷$?�mq�LkQH����$z���	{_�݃b@�vGKf���`��ޠ���Qalބvg�=��h�(��y�Z��e�1`-K��b�+T�L�;P�&���;�wΏ�p\�fC�/)D�:{�I�E��>d�/1Q}h�bM��!�>�3{��n^L=|a�LU��!���#����df?t#|��&2�)�9G��4�QW�F��.��zϰ�YQ_ 4�Va���j�$o�����=Y����U�^�7ʧ�v��߄P�+KC��L3hʕ3��H�z>$J`ŘKNrhF�����gU�Ũ!�X֮�)ܨ4f'm F�����-4Fè�Ӄ��r�`�ꈕ0-� E��Ү���HZ�Aޘ��xL�PN��F}�W�P�	Jc��eU���rAX8'
���2�P-	��2p�0K���J�q����?�}O�tk&?��R�����Vy,�ږ�y���cCK����:g�,���;�?6�2��S�Z�A���y9�qq�rsI�����2eKC�*xaW�u�*� �A�;�C�Ɲ?���o��ȣUD�!䁣�|�ӝ����ܮ8`�J�|!g]щ.1~B;�N�L��T�"�f��Q?D�q���������j��� Tѧ1�n��F�M;�:\���:�r�����;��!-�����v8��n��n��T�JD�z%<}?S�
b�p��8/�t�8�LD��/���&nd��J$�P���XM�0ci:��o��\ާr���9���ȭ��S������Y��w��~�^wHG9h$p��ݜ�'q�bK�j`��%G�jzb����Hu��y�p���wR���#�6��0/�v�>ϽZu�1��n+�Ԛ^��"��=ة�T�5�C°�@�Z*Y��$��I${������4]Deu�z�,J��*�&��K�TtpQ�<�'f#Z�0���4=����{FE�xnHG������R\k%.\m�&yk�#˅��GÌo�� 	Қ�
E�h��K��tst�T�Ɗ-8�LR�4����?��P���M��/ۓ�nT͍&���맸�Rť��_�?�~�2�2���*�����FDx
q�6ԩ ��:�?�Lj.*$�*����m�I0,�r A7�.΄��ݽ^!8���4`�pS�'���c���ѫAt\뀠fݎ�)�M� 4U�[�la��Ir){���2�4��R~Ls����D�O�ݢ��цdU>i�J�]��L�{�� ���h������VM�"�"�=`y�G�����8Pi��B�\�?x�>���}��;�PT�V����'���_lQyyl$�|����x���m��w��&�wb���>���і�#�	�0�~(w5�[���5�(�r�����2���'Uܯ�	��������Όes�������KͿq�%?)�V�J>1[Y:���p.�C�4V��iO�D��fLH��2Ȃ��w߼���b�cRKf�^q�{/�I'`�Y|TB�f���fO2�u`B@"��R9�5��v`��Cr��Owk͍���W���/�
�8ka:CԫAD�j8_�;а���M�{8��c����8���t&O��c���2B��@"�x�A��v����X��hG��u�]D�ͲA2���,��tZTW���GC��?A�J�/IkUe\�i�䗀g�*��/��7g�Qa��d{�+	��5SV���^�,c��z;<R��%�r�N�`���!5y�<_�x~�|zM�p��}cN�!�R�p��0y��;$\��B��C��IQ^�E��Z���lh:���<�1�5u��	�Ysn��"���!�d�����Z�ʝ [�K���7�r��*�B������V���6!e��of�s�XH�ͤD��'$^8��u�f��KB?R��F]�R���|�Kb�2)h���dL�8G�-h����uM� �X6����9����3�~)����y��]y�x�:[��%��+[*ͽ�6���,� �M`W537F�ٓ6-@@w�Q�v�B�CH������A&�Y^�P�t	����lkp�{K�D���L$������2:U@U?G:�����E����B[��ί��㦓D=#�_��N�������m��i����m75�=p@�엋%��,��t�@�>γ���穤吪y��P�=՗h,~w��3���.=Ck�xc$<Q�L���K����P5x�ԓ��1���T{�����Y^+b��n��o��V!�cO:�����x,'o��6X���.�����h�Ľֈ-���|#��cZZ ���%�'|/+1dh���V8��u��;���*�g���V�nQ�f�\耲浢t��ܱ����ׁ=�t����n36/�p;I��j�ȵ�iFbC��Yr���
��Jy�|�_�z�a��K��JzY�y}�0�|x6,�J&W�s,V���Pz�c�<�F�8瞋����e�rw��~�Pe���|줬粱��2���)3�r��)j�c��M�	��v/稆�����0	�E=�/��.�����x'����x%T���d�MG�P��._:QQC���="�g����Dwb�}h_���J%K<R�Y�oA%�	�岓�a��3p�����C6K�pl)�����c��Xژ�i�P*[�w ;�@��\?>kY]�����b)�s���9�A���PY�Q�@�Qq�H��Z@�gM=H���e�I�u��Rr�1���䣟�Ҵ�-�L���'��K5|����6�2'�^�*�(��`˨�k��7��x�8����f�n4���[�3����p�bk [G���Io*�!И	���	M��y\k~*�X�)�#<B�1�����͗�#Q$g�d�����`����Ur�ޅUъz��VP$�H��YJ�c�y� c.�!f�޲��W�(c�D���+-^�d$�+��_�}jD�@�;���i�(���Mo�i�q�A#�s��:�i3���Օ����+і�#��F��/� -X�fN�y����p8ט�l|���بa1���l6 ��o��ĻU��(���<.����<���=���[V�hAB�@�Ž���=������B�D.�G���2с7?�6t�gs�����.#C�"<����wVϽB�mV���W�>=���B��ϧ���Wdm:���І��s��N� Mn"��I6{|~{������OF�"ذ�JB� t�^��B���y0�+좪�1��;���X��M ��q��eq�YJ"Q-{�.�@�'c��A+�����|���9�+ү�nq4wF�i�RDqG�k#e8e�T�dǹ�'�T�/xY��/B�v��Vm��)aVb�X`�h�;��W[[�A�N�z��TE�"{H�ï������tw��@C�>�x=<�\@CR�\Ql��x���*n�N�T�*@�t�a���8�r����f�G#� �Hj�u��kc��mFiWY� 7w��@� �ςU���%x��c[�tr��gq{�l���z��筶�L��%��}��9���R8��.k<��g�����.(��7�k���c�7k	�_̂��������;q�5`�ٖW��[ 7�P�5��z��*�V������;9J�C��IW'�i�����Ow�m��N�M��&��O�R߼Efwq�Cy",�]�=�D���UP.LL�C�3�b�����/P�����[,6���J�6��K)c�Ep�˳<Sf?��a�uF`-v� SKH1��(��i̗�0�8�䴪��"DE`<D�Xt��N�T�Ĵ�����{s���'�i�)Q�J��`�Z���!�Ar�("t����r���7'�vJ���!λ�r/"���O���1}��S�4(������� Ίi��UZ7W�($	Xm�����d�Ό��:�5B�q%)aW��|��Ŭ4S�����4댞ZMZ\�
U�ɠ�<m�A�mHio$;z��c_�D����%"k^��	�hF�q�q��}�*n�9��N�Ǡ�����VH�S/p�����_�b���J�+bx����^]�����'��!.�J6�vq�p��TJo߂5��A�ʇ+��'P���3�eg�سG�Tϫ���YX�k�´�Lt�":�ZL�����P,5��Ѝ����ړ�r�8	q��M�B��;%�V��n+��.:x�8��ӯ��Qzۡ����z<Z�g�r���)�󑁝&�p��V��HԢϮ�*Ă�b"�K^���d�����A����XZ-�!�����A�Ut����p�7��8��^r+O���`k�ǌ�fڲ�l���ek��\< ��Pd��~S1�ڤ�	OBs.�=yr^��^����V�D�2��r6�T��U?^tzː����G[�v)�a���2��ij*�~��̥�����?�^tIl��Y2�I����!����*��j�����|��o��e�
־���Y����K�"�
*��%�}(c�0�ؖ����[��b���������3� r=WL
�63�i�[鼺tހ�C�����h/��lў�Ct��P�JSӵp��	3�̼:]��z,�݋�Oqi:��e���R������t���}�L���i=N�W�6�J[(�����u#؞FB��ZD{߸�ߺF�ү]V��"���N�B\i�!�:��禜���N���/�G���ٽ �nu9~�B��Ϊ/~$�d�tF�? �4���:�F�+fR�$�����TE�q7s���H _D �i�~w�/�_6=L�t
ﬧL�>�Sf�ϓ.u.]C��`�/�r��6������ϽpI����SC������t��V�����fpu?LZa��3��Q�.�"�}��.T|�^b�%ʩQ�L�0|pg���8��"#���Ӯf���T��"�f��>�m�t�D��3��(�i[C 	���kpI�)-�^��u��UX�����~7��Xr��K ���1J�Жw�|�,�c�^�7g����Z��-��U�����V?;R��*�.O��,r��D����"|���ע�cNs��q�J=܍���6�8^��I��a�%u���Y�	A�G���!ų����'{r��S�hu�E�����	F���畻D��8��g���@�AJ�֣Ů�^��x�F�X9��!Z�E�ŢR8*漛c�dh`��*Y��àd�[Ut���=u$��@����E���3�[*�~c/@���B1b�P%px��9ZA~p�����:O���㛬Y����;�Gk�,<3l����~E�[�U#~��Y�.MTf3�����B��|f��tyj�jy�h�q�5*�D4Ied�����Mtv�7�j[�0!�4�!lA��C5��n�Y���i����_:i��	���qLM����v��p�Ѻnh!� 6]~GDT���Z�'�P�3[�����F����\ݞ=Q��l�8��w�$���V�����������|��vk���ݛc	9Q�XV0�S�+�P�6�Arw�e�#^,٦ˇ�H����V]+��E;^��C%t7��kw�hHQ�k���Z�nԨC�s�V:0��]Zs�9���
��cY�.�$�\[��-��?�f#Zm�pOdW1 �@��"R�~:�}.��p��V�T{��CU�/���?E�8��@k�7Ww����*�G��.LK�Y�)�"FfS�@v<Ƶ��`w�8Z�����b�&���/�u�V`�QA ���F�%���(���?B'��9�xq��;fX��};J�٫\wIOP�~�.<�فZ�T%��U�.O��u����Ow,F涣TP^7��~���3k"����1�I�L����&�M��{h����� �!�mv=�"_z��}X�藾9�߷ʌm�lי��(V�U��!�v�@�ׄ���ߚ�;��x��"<��5�ˎfn��e��D��������D�`*��л����vs{j�,��	��H��RJ꓋�k�Tm	���u��;��M7���s���L��	�P4���̙�]jf,�0�\O�̶'�:�+�>Xv���w@�ě晔���9P�Q��'=؏��Er�u��Zk0��=����C�vڧͧ��S�Gl��A�Lz���Ɏ��5��d4�:1u��[��N#���Z���~;����?_��|�ѽvh(�o,Ǭ�wMe���'@lH�`1�7�=X(�[q����r���X�Ǩ���y
(��D(��_��H�N�a5���'48>j�������	
zͤj�X_�NUm�f����鬃�]�"���#h�z���r����o�Bd�$/$2����qyn�.�I�-�����^z~v�r��.�*�5��'�.Zx"U��DY��bAJ�lԴ<�͇�+�/S@�S��� ⡒��̄2s=��W�2�o���?ۡ�S�M� ��ZG'L�l�]�M�x׭�}QkT�"q4��/!�2򘨛�TJ�d^�d�[��~�s#Ty�)�wBc��_���\�����&�)�øIйeSW�e�?��tC��*�Bx;v�l^��B��/���,���HN̴������O=��m�{[5��{x�c�q���#G����_P�5�4���!0D�f�����f���ۣ��H,�~���,�e���֔9���B�? �>M�+s�A�z?�P�>�z�!���dxT&�}{RaZkx�Wb	�eXx���j�}b���T����d��NE,��ѱ��y_��n�=����D>b�b��_��n�r"eռ=�T����{�⢢���w=6-�H[�nIW��:L�юҬ[�X�b�B(��s��oz֦��d���AK�O���6/~[z
m`ӳCp�ɡL7�r�Y���1'�����y���F�>*�L��m�z�{�g�;H��!��P�&��}'Uֆ-����F������6W!�
�FЮ��c�{@_`{��@Z}�m�W��'k���k�y�� ;�$�)�h�PQ�N�(��&���1-�H��:��<�ә[ur4	��j�V�^��VS����v��g��_C�d�^n�z��C��w�杧��+�|WLƿ��x�����j���"�s����o5=����Tȋqr�^d:���	�T�y��
wEjJƥ���R�>�WZ��#��.f�-p�w�Jع�1�/7:l�L^������������ &����+�z2��n��}8JUz;��`6���@L�G �l�/4_����'x)�AZ!L1*�1)F �-|>a���%���9qMK���J X�q����b�2�+Z��~�? �Q]f1{,_�aKw���՚]�O�܇'Aҍ�g8�e/�%���J�I�3��	BD8�-wP7P��1xu6}}GS�+-��`�;���i���{Ck<����ó��t��j\�ĽJ=���*�'P��1	,V#bA �-�������C��<X.���j�R/7N�d���n�Q��I��?vz��l���$zY��"<�[&��L�k�W��7>��u�2_�g��1�8� �q��sͪ��'�V:0[�� 3�^���>�C�����")Q�C�O�������(�'gZ���u����X��#_xE���㘶�ͬFCxC6���SI;G>�D�"x"ٜ����;�Bf�op�Z:K����x�������C��@�� đh����YH��F����wҴ����r�8��K�Jcț��Y#��f\�D��o=���m�m���'tE�{�����ٕ �(�R�����Ӗ��<V�Ok�6����*�&��[��Nw$YL��RU��8�*,�]>4֒2�,�TF��g��@����/z�!<_��N�%pԥ�GV���?F,!�,��Ġ�a�:
6�N�0�z\Y�#4��X-@�{��&`+{Aqu����X{�^�����S��m�'3��l��|���`����S<Ϡz�_���e*G��b�K��]1;+Q�#��ҽ��%�z?�Wa������!a���V��O�n��[��ŋ���-�U&!1F�!q�:S�p��<�X@�F?����gh���./�*�*9�5Q.[��;�ĳE��-�WR�6��)�����j�3�̻�!)l��T�V� ���0ICI��y�]����-^͉(8Hr3�/o�G8��x�����,����x>f��P|S
YW�g���F{-�֛��V�l�se(��C	׊U����F����/9
��b����óz`&l71�)�M*�8nb4����*���UMb��`T;q�D��U�i�BM��C��0N���V������ȫR�0��S�r�� ՘l��z��7��7����8����|�J�D֓Ye1-6]�h̏b`��fP}����F���1*.@�-o6a[��J�`;� �<�#=8ں)�,1�le{6���F��v�y~[u�`b�˯��B-�N��h�F��p�(���R�h���!��^�RF�<[�x�A��-Q4U���JnI9g����v��i��D(��N���$	���?�����8�;E��z�����;�-ϻ�n@Yc��+��:
� x�E[�(0���&j��1��� z�oC,Gm���E����0i >�u�^�
�.���j�{��k��Z_�{XS��d|�� ��PNz�8�B5k����	t��x�����/�.�՞{�(�ؐ����Lj����#$
�U�e�ʇsȀ.��R��͵wIÚcfyH�Be�A\�+�0���A*&Y��2Γ	6���{6�U��)�I�/�f;�$>���}8�����9gGSA�5p�Z��h7�}��y�N5�՘D2'E3�J"����e�E&6n�Z�7��Z�/��o�c�y�,1�j%+�ྣ���	z�` {��\�>e��h�Sp�{
a��Ӣq��@D?2�C"b48'���)9�G�Ҙh�r�d����j��>t\����/Á�񮝆��tz�����Ǜo� ��u&3�|��G��
��h[��͞H��K�|�����;��E���o�T��`7E��O�*�З������9T� �i�4m�^c[ak�kT�[�1w,�*% ݰ#w�c�W��}�]*vU�� R�!^6�`I���[�L/};Ur	�<�S�d�J�p!��@�G�"��H��,Ř����׆+��G�`�@t����2O'��_[��H�x��#��׀~uy��ǵ,��������`���qwu�
�xO&�)f���`Q�3Ӭ��B1b׊l����\[l���o	�E)�qGp������UynX��g�E����!h�G{��J�����%�qy���te�J1WBs,��I]�V=����2��٫鈳=���^.9�����eg���N�	��׍<���ʮckđ�Ϣ�%K�1#.p,+��,�������Obk�$��������m��ţ�_�}��W1��jt�rQ`�}�|cd�<�ZsB��䁘��I�M*x�_-��!iI�
�)�{�<����ݑS�kԢK��q��m@�>(��.!?�����{����vdo'��U�ͤ�=�v^?�6^�%�u���ȍ�����
�����l��<�[h�\���d�&���V��L?G}H)��� �O��y��(�a���]���M��h�n�����z�fM�+��e����/��A�ֽT����}���
N���t�aTݍ���W�A譻�R��M4��MUhWd��K Z�,��<��mn��R�����H��o�s���{ &���@i�=�D�T9�~GU��Y�ѣ��1"�M2&��פr6�?�<�@tr��Q����!?��B��m�Ʋ�ot�?1?b�9���w�X��Z� ��cS��e�;Q��4��d���O��^�����~Q�G^�N�{FfB�Q����ʫal�ׄ��V�}���%Ib��/ȝ��)I���@��k�.~�E���C�*��0Z���&�|+9Ĵ�~+K<��A*�dp�tBa��M��v�n �~7"CmM���������� F��?s;���]�ࡰ�I��&\-3��s��9�"������n�Weܼ1�)��ʡ*ʹ����g��
���.�r��ԃ�9h'V��[�+�@a�cM��(�}�Nsa&{�pJ.@*�8�%��[����T�?�ǢG��P.�H^�����$�� ��9�˄��a֛��xy�!<Ž�Yϓ��3���E��'E�]��'�g6��`�B	�t��c�w�e¿�*� �(�+��R�K�
sS^�������|҂TK�έ�H"�0��w#�G��$\�l����%������(�3�s�ߔ��t��qfX@��M�z'� }Md��P�=U�����\:4}��1��=������� �������>� R�]|"\^lqv*�?�^�Q{?�N|�	3{ ��^Ea�&��rMd:�ֈ%��8�rM&./hr�iՁ���MT�:ļ�#�z�mܡ��"�ۦ`f/�;�<�ݲ�v�j������'����p��޼�j�P�J�Ale�n�P�]<��Ij���0��
��*kC����u.p�>���r*�B!���P��Mϝ��6�Jz��,C��~;�s�q|�&s��������{1��.p�ߜbK��%�*�߭�n������͏W��;(s&E�R?��� �b�W�_�IƉ�e���OzT�Z�]�q�r
�.�Y���攳4� ��n��Z�2���>4�|r�UY�Lvp�Xm�/���h�J����r���²FEP8qn|���Y08���b���!��p ��M�)���<����H��f�#�v�3���A��I[L�5.�W���z������mv�s)]��!�W3�ņ���k��ڻ-հ��F��^��X#�����A���ۂ�QmUm3�����
XZ�͙� M��/r�4���c�F�`Ϸ�`	����;��w�Ӎ��Ry��y�#�7���Z�;����z����%���/��k6͂:����}�=lI*p�rsc}}�"z���yhc"����� c*�JQ�C�Yz�(]�P�;�S�m��FM�¸0�t�ڄ�c���B8��l��0�����v���^�6ց���$�0���7ŉ#|JݾgF���4�A��3J�4�N^�<R<��\���~�˿1r��q�4��$��T�~5����t�Ek�$��l:r�W&| ��
�)-c�|5���P��p�?a�_��C��@�A=��uĠ�P����<�kQ���L��$�e1�9$^Ɯ�<Վ��B*���"b���П�z��ş�=��dp@	��HHY5�UI��J���0Gj�x�����u&@DXaM!���zB�w,��~}k��>��t9�;�GN��Vs�	��X��:��?Mm���X�#��C���vH��?��n�:�X?��մ�3T�u�U6�^�vs���N�MN�4��/Κ����z7L����G�S��u���{~E6�_h�̡@]HK8k\�Ϻ��8
�����T��8K�F�rDo�_���9RgUƶ#�˨\�����t���?�
,�F)����u�;��Pi�P, �E� hGŃh��t�w������V��/tNb��9=.,!�(�@TbV�6r<�ã�e�#]_��3�9��&�����7��u!.����h��F0�;&�QU��,�l����xUC���xQ�x*KԏRHݲd�b ���s>jο�g{<��b�J�d�\���2u�^]�����8������z�J�$��>�܂D�k����R7I�L��u�Q����NK�Kůqӽ[�}a�}�|�W@\8���B�n�DIX2��;x���W~��R©{a����,��;>蛤%��K�a���BU4�^��䷪���Ot�]�B#�c�%��|���OE�?�S{�αJ�/|��̂w���~�CM�ղ�:�M
pM���9��	���Q�&C�ۜ�}}�	����" �����=V�X�Lu�����5�&�>��Dk��D)@�}��Kn$��ܔf�\V��*z��� ���ƶ2��f����b(d%n6��L�0����wd�C׼��C@~���<>��X�1}�d��{�xZ�������\�@@g�'�-�Y���Cs{z�����Y*�)���]0�b�`�2������Ll|j�F��Ǎ���V�]o�QV����1��ǾXO�CWdb�B�F�ԗ0f`�8��q��}�Sz�����w�3���< Iی;�_D��.�ڦ,v�����f�e0a��F����밀�,���-D>�h/gh�V<� �O�7���J{8t���V�,r������.'.���=kb�C�F���*��d�A���@���� n�o7T&��׾�Й-�:�fB.�F��3L�(���Z
w�4�O#otmlqЌnA���c�rX���z��~�gZk;�JK|� ��X���?ש|Fjx
t_��>���;�-@��c*����k�@�]�+S[�J�[H��Z����ku�����y��"��!sͱ�k�(��GѯO%A�
�qr#��'[-�ɮ�c���Tr�������U�c��}�ʥ�ɁX�{�T��l�fڵ���I8s��B�(o��ݷG:sH��K�k���b(�1-��H%�p{7v�U�[�Pt�Ё��'/9+ };F1�I��Q�35�׿�%���{�0LC9�DZ�<ӳm�o/jQ9�ڈB}s�����h�C(k�j ޘ 9�?�?.:��W�+�(I�2 ��/Xh�Li���Hd,���`��Ih��Yo ��@0�@ԯv퓽�Lиj��k7�R]���O9q/mq�]:���5'L�`+��Dv�ʹ�T\��
���n���e_��b�_X�i��Mi3�\L�Y_��,�df ]!�U�r�Z�`������O�X61�&#x��l���`T;TX)>���r2��/.j��������^lN�-�+�3,��:� �$ b��i;i��C2�K;s���P���^��R�|����?��鱫�l��A���1z���J,9&S�9;0�� f�]��2��~:׍/"N���R=�e���_��:u�P�lC������;r�-<���}|��V����w����j@[��%���Ev�e"�b�I�4v��ri^���s-�L��R���Qeŕħb!��z�2줿��e�0]��@�ѵ<���2�︚2M��j������'�S�	�^� ��O͏�
��?�����Q7��ұ9}�n�m�.����ۖ�.�b�P���6�H�5a㧷j�/_hO��%LA�L�s6�Ll)�6�$��2�����
��ɮ�:���k&V�,.۸g:������ITL/�۳[�-\q�2��܃#c������(8O����WJ�L����F̊���~�#�<�k���뚪Z;��yG3����4�3<�*�΁h9�4�i.W�).<��=��8|^��4]��.Y�[z}H7�#Y����(1v�� �^���S�1,�\<,巹١���W���SZ@���E\�4��s�U�¸��)8�N#��rڇ����A貺끥>+�N>O�8NX�;��p��6������<>�5�#�����g��s�+�?���Cy�^�[+@	��X�.W�Le��?�2|j:�L�0(� [1=D����`0K��>����bqft�g3 Ġ7m�ݮ�iѮ=u̧�׷ū�а�w��G��RR[꼁�%zK.�
<H1��j���Ȼ�[lp�2�����_tx� }�3��2m��D��~��/*9������m�l���O�Հ����1�L�j�U)�ah��A2$����_f.�b��'�硷P�
[���8�؝�ձ^i�m����q���/j���ul��,�J,��<�FZ?m�U��y���0���IZ.�����H������OY���btW�x�H�aD�~�5��ϿF��Z��AhѰVt��Q�n����jC0:�Ԇ"A?�$����hyl���OF��?��a4�G&�q�>xa�86���6ⲍ蛚��r�	�A]Պu��$����W8�?��i��y��V�c\�`���F�4���Ҏ����P#���4�jD&��q&��k�d2):�aGKB	D�D�ήvQ��HV���SB,��~II#$3����<��!�p�cCҶ�c�ω��q��f�\��}?M�1C`x�����V��^�C�6�?`\�Cx�	�G��컬��Ѷ�B!�!.���w�e�ά�S��*?��@Ra-�V6��/�od����[u�U{��aQ�[3��|����U+�Ơ�0�5��^w@`Q��)o���%���0��q9�zS)
-���E��e�RoU����&���u�!_��F�tV�ß[v}�i����g���v�����DG��z�~�'&S���w�9�����
��'ko !�I���,$ߞWH�w�X^��QA��>ݖ�)����كD?�:r��H��J��`�̼O\�a!��u�k����Xe�__кF{�8d�Ve�"#m��*�|�U!p�&��:x�c?���dt�<{�ͪc�5����;P����������.�ͣ7D��L���?cDf;:��7��}-/�bhˍVkL�.�3k�k��x,�Ģ�3gV�%�E>���o�X�hYG���,m M�3����z�$N��j��(K�.��М"ˢ���)F���u��.ؤ�.S��ܠ��[/�k��v`�f�N޲1l�����Eg�lbVK&\y�w��������'y���{D_TEcP��l?���\�#v� ���KE��Y�!��i#��5;y�C-2��g�2o���)
�"�Q<ɥ��<�>��I>xTi�U~�|�"�;�8:�l<2�F$�u�Aا�S�m t2".�*q)��ީ� �������Ǹ(ֺuƥwZ�X"c=�َ�瘾A\���Χ��V�β`K�[�.�<�W}n"4_���� ��ݍ�>e8l�^MU������D�(��1�=Ʀ�+:�Rn��������MMW�萻��}��x���v���m�T1��o�I9f��ˁ��%v��IKb�{�[a'�����ᴝf7��b���┟j�
$[}>K�E�FKܳ��^{Q���2�c��x<���*�B!f`0���z8Q��l����PEoMo��>� ���"�,�G��֯x����f`�o��H��j�|k%
ؕ�i�Df�qӽ�3��ؕ4~d�7a좭e�r3Ξ�Z����q
9NO� ޑ|Q� �z����kB�.�^, ��ή�g���I�8���d�O�/6ǿЦ��"�W$	�5��nLߞ����+\���3=7�#>s��.��1c,(l����,��-���t�]�g�ԝ����Y�vc����=Lj;>�!���x�q'��^��-u�gq"b���Kٮ<(��t��t)��{�ub\x1�f�Ƹ��%��Q������R<}��r�OcG��>����C��'m&����,��7Xzs����/����_��O��D;s�Pn��U��&qoO�4!�f�-���K)��E�ɪ�{35`(⧴@�������JQs��$r�x�B���������
c����Q�d:??�J�U��%��uSq�S��_i�oTN��a���Чi:I3F\�]�:D�#��Ό�'�q^�V[�w�3 1�ͨ�s�Y�` ����5��&Q#��w�2;��A߱{f&�� Z^���=���̺���!�m$�'¿��"��4ޤe��	�
�wh1/
��'�ܴ�:��g��9ޔ��~ۄ	=�����5����?6�n�����\ŉ��1�Č�I4���h�c������`���*i��a>1������[c�Ӷ[\u��S��yI���Q��jG��:���^�,S��	m���]����2������L�g�>����nЗ2�6*�tA�m[� ey�~�qx47ͣo�Y�i��6X��༨0�ǵ*o�Ϛ�i��Ҡu���m%�m�^�uvhĔ򉎇7O�'$X�n
��T�I����W!��7"�yO8'^����c��MYC��Ċg_z(gG3�QR��c�r�{����� gѢ2����>|K���P�N�l�ˇKY��1�#Z�E$���Gߢ�7c���ڛ��x�<�e��3P�*���!�h�c��*g���*ߘ����ϱ���x���Li����G��^D�V��+��%���Gvq��f�a!���F ��Z�+7yx&I��:(��iKm\"]�[(�>��\�Rʶ�6v�;��� ��q���Q���Y��>�O;
��a�fd����҃V?�1'\�W�%�x�S����I�4�65��=d���ןIğˢ>?��ÿ�eONF�<�m ��m>��ok�Wy�����ц?4���M�o�$���-+��D�/�<^,H�Z�����EiA�����Fm��h���Y��'i�Hh���y}�˻=�w��?�*=�|��"Jn�C�fNM%��J�,�/s
|���>me�����\jV�/c�m	W���"��Ĥ��a0�;�q��}g��N��z+�g>K8�)Q��1�j4�y���w`q��
7��&�ZcjT��nP}����t��M��d�}�`
�%@R���硸J��^��箫e��4�����]ʙ�~x�[�E�H��L{%�a�=OֱA�"3!�2��2 ��e����7pF�0�ZQUKj�Rn ��K%�!��[��K�͇���FD�;�����]j[�~���<);��8�~9o�=���.�)�AF~W��kت�u�B�5�5S���|Y<����@l���֜��(�BHz�!�����R`� 5+��4����|��?8�H��7e�
��Q&A�*Tg�GD�c����It��[�ձ�׾#��RN�݊8	M�t����p>+��ä́ӨZ ��ۿ>�v��w&�1�ʉ�'ڛc.9�fV���	�������Dq���s�?�Ը�� R�
�PA���4Αú������x��7�g<��Ht�α-��}��p�d�A�����	7���H˪�dyl2C�w-g�<���g=q�|&�w~׎�+^.i3��Q�
�>�)��4�[��@�Hn\͹�R���[�(z�&���ps�T4��7Ц�i�,ǕMj�=�H�s�CUXiy����Ϋ�an͂�3��Jtʜ-w��W�lY<"2��QqC�%k���\q�'��ͥ8W�=�1�U�j>Z޲����ot����֪+� $Ɇ�-g�@X��lY��
�����7�i�M�O�G�#W:�ww�h�QzO]�����u��ij��ѕY�xa��.�R_��P6��F��7��Hf�?[s­��^�h$��!,:gS�hRtKvCϝ�d]�e��q0����\m�~?���-��U���[�>
Ǌ9/&(�(O 6n>�t���l�>�;�>49 ��	2D��\ڇ�$�B�O	8h��l�X����}�THw�۾v�0
\-.�3^��O₤�� � �6Ě��6~�"f��F::tA�Z��P��F�ʗ��rX�d����j%Uo{�\=���z��0wR�z��e�N��ӱiz��$Gވ�b�^d���'�*�#!800�>��N�hyv��>�}y�>=0��*�;�:{�s�܋,�E%��N�ԑh�;�mZ�Y�+(-����~�C;d'�>#���_ͭ'>L>�DX|Y����X�̕�I�,�������vou^��F�������͢�{��t-c�_-��H[H��ls��BJ7yč��/���J�l��Q�������t�G������*O5nt�D5H^�Z�����қy����oj�Ў���y,���Sf�.ҝ*���"�~ya��7�n]�6ӚBST��j+�kXGo����#��!��7�lUܛY�(��nBj�ieh���=�Z��F@���x��&�� �Q/;�Q,���`��V��S�]]��4#��+k���O��{��z�U����]kV�Y�L����W�0v��M�c����0�6�b��8��������3й����i�#��zI'�z��>6*�K�՗�^�ێH�r�ן��2p���g+���wA����l�v�����yh�ΞF�3|��,^75�����"z�E]p6D$Y1�F��M>��m���;�����&+�f扞�i��>��;���1�0�d�@@~NDDC��OEU��7�Ů~]{1��K9q���/����\\����$aӵ�Z`�g�#(�jd#o��I�Y��%��=�Ȫ�Z *J�n��{��L�,d���m��g�ir��e�6�ʬ�ڢ< Iez���Ԭ�D��)�^nڞ�Ϟ l�Rݜb<��}�v��\{d�Cg�>�lT6A�_�z�K7��l~�)���
��6�;�5����fb y����EM����TΦp���
�n��O�IuE'�Ń>�X�B\&�����x��1��EC$�{�>>�X��&#�S
�g�( ����j����A�8����\��>L)���(����rS'�i��f���ua6!�3^?��E�g�7�F�J4����tϺMo�w,��ts�IE�Bs�N>��y7��q^�*�9���z�d����ʍ��:&�_�j�P�'�O	�d�C�|��x��x�y͜��P�l,<HX��t;��f�M�2\�F�@��X+��� Էt}V��ŎQ=�ch��R���0Nz��*�G����;�"d��� ����P�T1�7[j�+�D�#6�n�e����/w<�wum[+���
5�j�����1���cl��a�j�nK���$���.��v��*;w�H�>1�9%DCFh�b![?؇'����=^5�l�T\���(��s0%�fF�Sγ��//]�]�qT�
�������2�Z�YJ�o�s[X��I��g�UOb*�|�� MwA�8�V5���Z�rVz��,{�Q�m���Ł·�V�^�mUcE�ލo�$�ܕ\׉����љ�G�M��\��[wi8��OX;(�m�>g{#����O�[ͺ�Q���^2��Gr������Ƅ41�a�����?�i��z�\VdJ�&�9rj��'#j�W��(1u�U�Ճ��0̮��Nm3S&u6A���
*?�13>�~��q�G%���&��` ~�.�����@o�pqG��P2�+��ݑ�!Y�G����n�}�jݩb�]·b̹�?�||�l�@ڂ�Z2��y	sucĞn�Up��Zϙ��t,�b��F�W,���l��d]XD<!]���WٲL��{ɳӃ�]�Hs�;��0Y��õgXl3���><�$`��J%c�е���!�ق=�tv�!���	ÆhCR�\:��p�'�����Za�qz'C��������~����d���6}�+6�jQ=�q뒒��قBͪ��|t�_a���*���c���ޖ͞�v}Жp���i"�$�?
_��A"e!7��v�dٗ6ܿ��r��!��)I��Iؓ���B���&��愿���(����Z�N����jn�OcS��~����W���t�"i�|��O�ٵ˄+�s���{!4�ٖ��b"�*�Xi��fG�����ҪXGETK� E�y�'�N���.ݱefY��⟉�gjM�mr3H�0@N�-�70%�xAT(|!�րZP�G��lG�U��ZY0yӮ��i��AH'6b���w3$�DD�K������PUwف=]��'H����Z�˾ �������+a�߯�:��o�T��,����h��*�J�ڋF�?�M�C�Ɇ��E@EB��#r����с���JK̊�#����0��8%x�N+�`�8)�{YUSL��"�ܪi�E��ۅ�K�KƵ�f�?�\8M`��ߦ(j�>%���7�3��9���~��5Z �A޷#�!�n��d�Q��)L�҆I�$�<A3 D��v�0iWT|#M �I���Z8I?8D�$j�F�Vu���[P��6_����bz�IsD^�h�Z�p�����B��D?��ߎ�gG���ũ�aᒲ�{�V��߱ү#���Ͻ]��v�I_Sl��g���[UB���cՀ�p;F<�GӬ� a<�r�3������kQ�4�o�k(�Ì5mh��2xi��RϿ�N�|�<�Yះ��b����G�����q�H,�l�%!h�R6}��I,fW)��#+{&�\���h5;ld�Ks���/���~[ʆ~p���o���� ޒ �����Q�*\kw�8���k��Z�e�΢� �٩��T�F�Է������#d�m4��i��AG��P�'5�J[}�!�N����8��(~���a���m�0%�(^�I�-+��~^� ,)�L;o��ھ�O1�ю�5�A�P��	�d�+���6�u�>�vE����`�NL��v���R�xbw�g�ng�d�b0��@�bۆ��,X�U����V�~	T�ǹ����טzX�����'�_<����;f�&<��Yt��1(��M	��߫�pr`׌����䮳�o��T��
l��Z���c����ď���>\�����ܢ�ίa�v�g�4�~fR����z5IM�>XAW�#6���y����U����(�Mv�9�@u��_��§�J�����,���E�$�	�������D���z��܋�WX�H���UwÛ�d7��Ē�q�h�M}��%̟� X���ۣ{bs~���zL��J~}S���x� �o���g4�=�
ѧrVt��%�F
v%�4��4�	M9g�o��R�%�H(�%���������N-�g;�d�Ie�,�'�c0�^��}A:�6����c\�>YN*U��b