��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0���p�?�gu:���@�6h�S��藑��T/���y튼�J;:qD~�'	�r�n�ĺ�cy�` !*��흀��.�Q�h%sf���c��L�uo�s�\�c���y��J�(�{�h�ʥʓn�W�Q����1�Ӻ�@�|􋍂 z٤81����>��'N �Ds���hأ*��k�x/tK��e`���X0�*1�����Qw�A�
�w�3���m����`��t�u���ywM�n�bYw�8Y�
�*�|���/C`����*�
�)ϧ�0#���ӞN%2��Tr	�z�D�%-�w�P�����&mHnd�����=j�aA��J8��
?h���Y5�ɨ�T᭧/��֐'����g5Wx}���0�6x[Up�7RP?m�#�5��6g�K�9���4k�v�*����(�G Cjz���fV9�fx nPp��a����v������(�B��o�pD���FQ�9�$[�ą�C^y��#T�[��*�ޤ�M!d$�<K����4��I�D��t����NM�5*mCb9�<�Zm���N�&���j�f񉶘}R��@�[�>6g��@����1o>��� �h6�S�adKf.�{�N)A&�I\t�Fq׃��	��e���8�_��G�,�ϰJ�ǃ�~9I�x���="0�����r��Z�U��˻Zj��9��ˑ�����G��;�)h�n�_�Mnu_�+�O��"i�0�{�I��������|,ehib�N���ڛ�;9fjoAw�MBv����]}�(m���Q��J^�|7&��/IL��əW��i�1�R�C�3��vt�Z���R	����o*z�#Po�!��QѠ�K�t�v� ha�����g�̬W��3��\�W�A,��f�}~��8Na��f�o�A$b�0����%�����Z��{K�O����Z�9��`�TI��7[*�,B��	�ۄ�jFAS)�Ns�J!��A/	y��|��W��V�41=Y�cCx�C/��atng���ט�b�`C�1�M�7�Izdg5ǯ6�z�6�-�ƀѭ�O�=�甒X�B#��Lc_�W8��1�����!}T�o����]x��m3�b�z�6Vx;j���(�{���".P��MZv� X ��FG����ſM_�f}�f}|3�f��r�u�f�;�_�����D��(�&��ԽWk�z������͙�eHmS�˨���#焺�]�z���G�P� ��ւ��F�EY�AS ��%,tT-�
6�E*�ķ�V��#�zyO�,%y�'���>H����jG�K���jR�n��Ma�+ �nh3��r����nr��ho���#C�h�^��A�M��;oT*E��pB��z.�_��1b|:��˶�H��z"l�-k��4m�D�o!���+'6X���5�[�=:+,A�0�o�VF|�ҵ�l!8Čo[ �!�5��,�Z��Nw�"�h�[�&`ކ��i���d��2�*I�x�%\��c��[���1>8�ɢ:�-T�H�2����@���{��:�P��a�li�e��h{��Bw�����#�]��� d����j���A�'��}+βO��Y��M�D�<${W������>-D@�-̞��� ��D6�E�&4����y��Q�gr�,s+��:yK���cE�?�D�KSX�9��hN��\O9�U��&��Y;kѠu^t��z���/��"��Dx
`�ү��g�l���י҆J�=���A����%�����K8��?n�	�Ac����p�El�m��\,�d�$%�3��j���J���z$��G�����i哈z�Iw�ҏ.$� �n1����z���A��+�7@�\��?��W;��y�����v��f)�;Y/�`���bp7���� �l�CtN�Si1���V}���>0�x9 �f��M��} �����Z�|U�)8�A��A�O�1��Ʉ?h�������%�7�v�m:^r���;�7����$i��(�v$�[F�"�ۊ�T�2���I!E]�C��vF�X��ȿ��� �HzfO��`VmU��R:p�:R�أ��\�i�#.MC<кJ�:A��i� ��y�Mk(���$���	-$rU�ܧϗj`�{ۅ ��nWu�x��kG�\��h��sY��#�����ԥht�ރ�+i$�N��{�Ͷ���*0z�m�P���n��[&��Xi-�Bh[p)���� �O���0��D��x�Ț�W�<D��sN��?�j�y�r�*p�#�t����R3QX�u�ʦN#֊E��{lr�S�C$_���ǥ��I�	E���<A��p����:�ly�KE)�Sx6�q�xk���G34�.y�*-Wz�\��Z	�ј�y���});�@Wz(��������#R�x�P���<q`OcI+�_�+�p�ݩ(�K_BW�#���c�o�����!�=�f��P�����5Z���D����XT�7m.��s�V�_@�H/�C"q��)��[��-B�Z}奢�l(��#e���N����ߙz�-�0�X48C2rҭn)[��"ȩm�q��p��B6{P��׍�s�iPKM��'
!����1a	���N�a;wb�X��$J�z��7X|:0����)�#q<�o��,��ؚ��K�jNk�����^Y|�uQ]���b��S�������vۡd<��@"�dHR�� w^�C�ϊFW������+���fQ�yn����v뻬"�.��`m<D�[���G�?�b��Rs8Q9�ӑ���;�V���
��	mL%'Cqv���ʹK�VQA�$:��հۑz��4��|l�	�r��n;��LT-�]��'���_H���;������� ����Z���p<�8WH[iG1�[�||n|�:4mڢf`>�O%�՘�PPL�~��ӛ�	������R�>�G��A���x���%����h�G�^���F�>�0����j��p˴[΂���[,eǿ|�#�|j���W�¤*���'i��;����yXm��~�:d�������Xk�%�"�tz�M��Qߣ2J����Z����Y���&t�d�+I�ת���O��w� 
����[�[!T��/�B� �@<@��h��IJ(���##ϕ�b��8*����W���F��}I*<�6�nyhT�5Wo˕��ԒG5��F�/��`�<;XQ�_��^Yc��}�c�"���'�%kH�Ѻ?���򉄓>��E�J嫣%�1�����pp6{ *������w�r�^ČՓq���YU�\�Y�8�u �_���똨��,-V��������ۜ )��x���~~��Y�ӕ>)�q��l��u1�(=��3S�VPG8qɣ��5���YS�]���bc�8w�Ks������?ŭ])�� ����	�!�)�纜�ot%<��[��nJgb4�&��D�Vo$�^3��ݲ�cB�����f�//J�́B�ˑ����	�^O��ڧgkĄ��ϥ���ӯ��<i�ɥ�O��l�ie���
�3�\���;P�E�_�ϸ�~��q*Q�CV'֭	\�p��[����t������M	��0��xz�����h�7"5J��j=�a�.��R3�8�ή) n˨d���ز��Y���}��Trbo�!�]��GTS�`�$�7��%�b�����<ES���zIJ��P��4�8+@^�����M��s�l������GL�߭Ɏ�/)�/�g'e���F�v��L/���G����|�NV�PP�ꨠ}j>ܸ94ݨvx�%x6ct�
�3"=H��#�j��e�uᎺ]ޖ�
RhO�y���4�^�� e7��@�4�ٕ哂��,�����U����j5�p3(��5���73�/v����BUd�dP
?���y]�8p���5x%�t��nD)��U�p�շ�	O���5|f2���?<u9�T���]$�C�?婞'Q(JS�N�{"똜����Q���/p��y��v��X7a�ݭ��:�҆é)o������I��I��-���*���r�ޱ)p�۠R��r�q�J�+����M's�ְڠ��K	�،��M�~;�Hwo�T���cG�:�d/X���[J�*f���V.p�P�f8�f��C�y���N��?�� 4*��� S\{��sJ��{x�����~�$��:���a��z�l�D�K(�Ϣ^����&��%��4��$��$���a��&>�S�݅߹�Ș���5<ﻤ��'VG�x'����:&�'�VS�u�� �XC?�.]��Ǝ�c)�[I}(�@�:Fuҷ*ѱ/lU)���ߗ N���3�[�D+��=Z�`�#���p���n<�j��˧@c�*$XO:|t�i�Mv�"�É�B��~��W�i7�1|��料A.��S��aF�CwB���:�N���E;�T&��}���[Q9�]Tn{�����Y)����@���[ܐ�	�����'v��N�[�� �����}έ%mW �,B?�7��H���u$�z�}��� q�)#�dȖ���j|��O(���7Nr~f�W�K��B�����<$����J�n0��oaSӱK��Q��w�e���0/�W?UA�w�;�ѣ}�bt	���w�����<�_��Vo�Q�G�[y��I@����̦��~t'D���>����E~�����zS��O�Cp�/Dj�W�7X�s:b8#��8�/Ia�:�(�Zl�)C14pøB��~�� �+�z���=�0L�x!ɻ������X�tb�X~�26v;��E�8y�J�C�b�.������e>����w�o� v,E;�HK�TE�� ���)�< ��CB��^c]&�����$�ڸ��:�j���đ�҅�|3Ǐ
mbM^&��!����y�>�'�� ����}��FZFM�3�P��h.ڻu����5S|9i�n�퓵mLP	[��y�Ц��|4z v�j���}:i�I�j䷼zߣ�E�,�-�YVzg���zX��_KXF=���mZ�<cqh��Â	H��تf�U�Z�-�7mQr�Ռ�HG���W:��-�_�f��[�?3�
thY��WB������9�`�@�f�b٣Y)!zn��Vc�q�o��#�~�]?�j�x�%:}@o��=�M���Ge*��փ([ѡ=\֢��]�sܺ7�����#��?���?a:�3J�O�"��F��uD���G��.�,�F�)�(a��4��l�<�5)z�4�{�0�9�x����pf쾷�3�*\�/|�zLc�we�7D٭���U:��1W��+E��:�M]P���_)Z1E�Ԩ��i��_@)����K=����Ŭ�Ǌ5q���ís�Fk_�%��P���}��or7Ì��&ӝ���x��]��7���/گɿ������g�&�?g1{�'��' T�{%8*�W���'����np3*�Dt�C���X�e��.��5�t;�s4c���i��h���� ��� � 2=�mM�7�
wȭ6Mz�U^I�3[b��@�H$�Q�𹴘L#R����4���FW����V�)FtH3b�������Nm�%��VZ���}�u &����{��L_Zh����U�͚��&��6�Fph$q������[���O����2|���d��Hw���i3Щ* �ݤM���ŏc� /��	-ٕ���og��"NZ��5���31Φs�e���s����\ �H4��ό�6GE&<I��wԛwz.��P��V��,� ��Y�^���&G�}�Q��燓t���oT������~���f,S��G����B������ �f 
�A���Zo�I�����n�
�/�%���I%iz�$!�mď�	N���i>��C7�_��ùeɷ܃�� ����lY/K Ṉ�M���l�����N��J#�i2�3we�^��s�-N��4쓸��~��R�?#Ik����Y�|�|G�m!��-��!{�c����{Y�|QЈ �4�s?SH`�S[%_���$nY4��	���I��ag�i鉯Y�b�lOh����be��q)��[�lpo�U��A�ʱ���dN��:�u�C������b��uI:4ȐX�8"ރN�����ZJ���ׯJC�b�jg��/�Ƒ�����r����i�m�xmK�(�4�*��(nԕ'S{�=��A�X/�rqFv��my޲�w���rB����f}wݟ��J�����i�0��q�s�6} Թ���_p^o�]�g�Ɨ����.1S��Q4�s]��@hpA��0�y
��a>��p=YR^��5؜$f`]��J�J�l8�&����f��!�[εP�4_�=��=A}�J��v�6�����4I���ߎ�]�y/P=�̉�
PƭH`� A�s��5�Rϣ_R1�1y��zV� �iG|�`��H��ª@����c�֫�	S�7��Z�n+�]�}Vν�!$�����&G��
�wVԅ����/��тE	xPw�4O"�}�ԩ�q �ܯY.����6_�F<�+�r1=�ؿ]&��Ⱥ���jrb��oּˉ��а;�,�ӲU�cM-�3.�^^0O��D�E)ED��%4)�c�[��]���-��\�n{6O�����S�CK3�?9�r��g��!#�E�чB��)�y�o����'̊�cIq{*�$;-�۟���i������T���:��1�s�J��*' 1��B��n���G�g��O��uږdP��na/'T7B��~JNm��&�X�͏��	8�ߞ`�qr6�`�9qF�y��ؘ��rbG`�~+$�nt7�?2$1g���ٳ�oW�V�x�q�^���L)����<�g�҉G��O��|Ғ_RS/5��!�d��A�������{�L���0�{�g揸U���j�
k�K�Ӂ���\^��/���]�9�x��+_��?Dׅ�����uk8�
5 b�A��GB���[&�Y�d:�Y�C����b9�>������߼�� &\���r���I�Q[{r�8�唄�*!۬�_�#�6푒�lG�)7PO�O�j�ӻ�{�kZ�uƍU2�s�	��tsY��2O�����&y����5�e���O������{^\ƫ�Z���|�lL|�>���3I6PAW�"ܷ��S��_8Yۢ�ʀ�>B�r��'ϻ#W U蠒s2��(j9��L��{���z�&^u~?w4������(ȁbh����C�>F�V��0K$��:T�|ү�}Q�s!� �����z��%����<��u1�&u�C������kzO�<����g�y��������*�M) �m� /9N���վ�,%����s�~F��V>t  '5���Ϲ�i��@�+⾷�M��n�f����Kj�q
)?U;�@��G+��jJX���@����A�R�/*��o� �͒y}�5�u]�ڳˎq�YNbp��4�:�zq6�|�>��]7y�E�feʵ��Px�s��8!�]s�S���S/��$1l�;��x/��&?%�� �I�`�#�]<x�Ff�t���I�0X�-/�J�Es>m?䩑�耄�+)�O���Q�ˤ��@z�fH�0����ܒ�_��Ww݄x3�f�M�zpF�N��=�
�=���)Z�j�}�Q�&7�M1rUkxEM�w[��Wo��
�$!��I��O]4����.���C�J�Q~��M�)���m�{����� ��|N��k�����7M��8H`A�9�&���N�W�kKUF���sg�z��lƌq�m��m!@����C)D}Gn��~���w=��Z���j����b<_�f�r�̫��n�um�҃:*2��2��˲�&$s����TNGV���,�wm%-?��n@�Ud+G����0�"�kOTu��S�8Y$�����󥈦�q}-��
����f��E���f�AC�+����	r�c�Ӗ�]���b���\��d��E����(9-�n�[�;"of���/W�I�
�a�=3���� �#ɝ�f������z���?W�̪��z���?ov�����I
��� r�"����VF����2+�c�ye\?Y����@h@�KL�$��6�>~)C	���q��c~d� ��-�LL��L����G�"t��	АSFj����*;���ji�T�7�2�W�6QTa�L|X�U,52����$�*o������ۏ�|���]�"�-L�Z�J+f=�X�d~oK|{��6�^̊�� eʥ��۟>�s*8�H���d�0͡1m$�@�TVAu��X+2�?{�N�Y� ��D�@��J��+�p8T"�Kܚ���5Ԧ�	���l���3���[_�������f�&�<�/莃M�XoL���U���KS+m�Z�^s^����a��;�|z�mQT�;���?��ɹ�#�����r�a�ڟ������rl�ѕ+�~�BI��٦����)��i���ПT4��������7;\�J�0��^�QR�yv���=Ep ))l��e��	��ӓ�)@�&Ql���ݦ7��tK����%���/�`+��o����5���8]c������X�ĆFM�� ��$id@�N:(�ŬE��ן(ke g�nT�g-
c]������Rc3K��{F@9#����w�����0P�Yh����14C2�tElZg��@B9��؇Y\��sYmfC��#�ھa���� �!ȜW?��奘��ՀL�iG�76�%�dy.f����@�0;�w�QEK���&����xa�D��)��4g�MZrYgG56 ��p�Jǰ�]3�o�n��S�!iv�#d���m����6}�7�C��X��DO���6l�LMV.��j�ud�4H�z5��*P�3e]w������W�V�[lհH����%���M.��=�>��g�+z#K%�$q7|����SR4���_o���w��c@�g�����$��_��R�}��d�7�կ�D��g�n�rXM 3�T�2��s�-��tPBxR�5Gf����w�/k�e;�/��1�I�sp0$�����CfF�@j���I�⊂,�����|��cvq(��.��orUw
ӷ�h�7�2�P$���"Xd7����/ �~�x�{H�u�NҒ��!pl(>U4�.1Q�?�X�F�����)b}�J��;�U��`�V|Z|��*�;r���q������Q��.��A����N�|-T�2�I�k´�ªH���ҭ4�MRW)OE�Z����(��0�M�7���d��� g�t!�,9o*^o�"_C���f
	)�����xM�p���_����:�z-���;:!^�oo�[�[������zZ9��}��T�  q�3B�4U�?�aY�`�5��t�����F#[t�4U�/T���2=EvW���=ޔ�i�v��`
�\��=��*���h�Yծm2[u�U3ڡ%p)�����	����:&i��B�!����CyUJ9���2��a���5�f��A��O��ŧ�K�.%rZʢ�&Gj;t�!sL�$f�;vS���2����]'<I�I���uO��eD<1_�9�kU'.x|�"�h��oL
Y�"�
��>�&5/���>%�T �#FR�(�.r����:a��`A/����3���4E�nM�F�܏��F��΅Tk.��%�(� �_���kk�F&r>�	��9����"�O�@'�$���بϑH��wb�MaE�A����|�3=����|��O��Q����̅��>^�U��|�5�CDl-gh/*�ފF��N�lA~���}L�|Fj�à�nX�7&b�%�x����'w�)��7�c]bS�ķ��Ĥ���UY�S�z8�3݀ N��ΊW��f^���K�d�!���=_���kZ*�� ~��,���]�Q�|����N���;�?����3ǗNx섇��9p���M�ƌ2T�og=�����-K����,��u]
�,�[�sZO^�]�Mk��ϸ�rh[�^5��V�R]��NZq�F�1�7�/����%��ˀ�*?�������&���M^Ga8Dڌ�EP�S�����ĸ�:k�l;pR��f[q����d]ҕ�c��Ɔa_O��®<�')0�[��,ɡ�M	� �/���4�8(0���C���V�^ɢ���^s�aZu����'��
l����a�����ѕ���O�ׄ�L�İ�!+������@UЛ%��q�$i3z�j��z�l�d�4�2� �q���
%�s���t�E�)C�i΢&��NT���@��}?*�4L@g-'	μ�%������<5{�d�@P���)���TfB|�3����&�kC�9,��&*�8s���-�ڤ
c�*K����p�1[2��P��q�����d=l���]��?��͙[�"�:����׍�0�A>��m;@�;r3|�=Z��_�?��i�ֻ"���̞󗇟F O���F��%�^r%�ec���p.v���HG���]CZL&��D�R,��h��K>�
6@�z�sOAϻ������`~�R����V+-�nx���Ÿ�Xx�օ�h�l�u��ť�[�Zv��W�QK��C��L)���4��
DZBĵ!;.���P�������mנ�E��H�$�Ҧ�#ou����]�6�:�������
�@�}���I��1I+b��À_"�ӓ�4��p��¬1�p,��y��O��6��_}W��ӷW�n��$S�a�@r�"��T@=���#۴�8c����(���OD?]�aPA[ ��'�K�W,����j�܅��'�+�6f���n9�u+�1Ϩ�:�"/Ԅڔa֡ݿ Y���@(+X#h /�,�}�FHq��B獎 s\ch�*]���3���H߅�cM�S^���Y���q��u|e���ISS�S��kZ'�^�ɱ ��32�¸E5x1n8��b��9���j
H�e�lN�UJ*_��9���"w���쒆
Ͻ�ך]�;ՙ�d���o��L�\6}AjV�o��8]�_^���wݩ�6=Y�t�����J��=qXnǑ�W�;����k�Y*l�R4]�,�S_G��12h!3�|�\�M@;Ӂ�V7l_a�\Q�I�x�щ*eQ@T	$��5��[�盳�(q�"~�FR�P錳�.�&���(�N�EL��:��]t7��EmWۦ���b�� C��At��q��)`��t�5�*�U�O���~E��/V�D'H���Ϝ��|"�[�B�m��Iu�rfڷH�Xq_ð՜�{��j\���D!�'�?��2V���p���4`��6C2�M��Ȟ���Ԩ���O�z�K�WY�54���-�p�O�Y�Z���& �k��,Th�g�P����҃U�,�)ӡ��ԥ�^�����]Ych�(��#S�3��V�J��v ��f#���V�C�/��"Re��#>��t�����1�ۜ�1� �}��h%��<��ܠ<Q��'�����{�Y]�I�x���*e>Ps��R	���l�fx�A���RmKX�=�@��/X�֯��ϟ����U�t�dæ�.��&Oh�CA>����|d�?m-Ot��y,=�H�v��j>���������W���F������z�ߠ���������
��3d�$x����b������D��MS�����d�K�nK*���e�d�2uu3�y��s,�;ɦy��2mt�w	��)�� m����dc�TDI�\��B㵑�G�jB����&C�_Z����VKT��F@��5U"ۓY��߫��e�cb,��%c%6K��'$�b5P��P�R;��+|�L�|H��qQ�5oɺ��:����T�� �F!
;fZ9��7��\!�\H٪^�N�i0���-��|U���)�v�Sk+���n�X�9Z�<x��k�!ʖ��0��pÚ������(��+�
e���'�Q����QT�.y)���x`~�g35�`�~�8�n����2�,QЂ�#ݐ�L�r��(lڸ�;�2u=����0V2<�WC�U��Vj�.��!%��w��V���-^n�����q5�)��)0./3��I�.���?>�3, �e�'�R�>��Ƕ��¶�u���{�~P*/B��=���I	��!k���c����n2�>���r�:��馍ųk&�l�����@���ҮWYr�Z�A
1a${���w�s��.����Gf��z���{z��ArG��D�#p�笄��,\��ӭ�3���\�g7ᯙю�f`73}W�v�i"��"�����%�E�,�K�t�o��a�i|�9����E�|9��ѳG���R��uj�;j
����m��N�f󍬡��L�$��浛��M }�]�P���Z�l@�ᱛ%2ڍ�a�A��"*Ӊ�6�#�o�G�۝/WB�q >����xb�2j#����:����gV�]"��A̆�tBC�'d���^Ԕի#�jS	��+PL[l)9Uj7)�P$���la�T~L���!���? �8d���$y�L�6q��6�.D�_�����M] v�]��x�ۮ`���w���|ӥ�иc����n-�O�}�s:x�~_�5�1�6����������'~c���:�3���&�;��K �j\�-�i�p�NPmV�A�N;�����u���/�o���AyY�%��<�'75�8�d�e��#oM�੒Z���H���-᎜׼��"��<�)�����0�f�G`X��f�Jvs�����j/8��.���g��/@%�,'�ҟ	�{�;G��G�����d+��I�$.���B9�@�Sቀ�/�>1�.�[*����a��N�dOԐ{��)*��K�~*����ڕ�,�I30rw�����r{�A��Xl�k�� ��ϐ�lǖ�9��T|��|S��6�0[���Z���E�̬k���;�	,�	�&nj�i�=>yT�w�1�3��m���o�x�5ҙ���f�7��t�9
%�p>����e�ͅ䵮oe�6����kl���,�;K�Z��cI���>y\��������D�iX��o��؏BOϻ��S��?S�KLU��F3�3���*p#��lh����g��й|  nW�K+�X�Gd=��=k>!=�%�S�H�|Ml��r%v���@�:źԂ���֊A ����W�
}�\Ȅ��kNrN����B�W���ژ��a��������τ1}��µYv|&�����D�o9"�S�U&`E`M�4m�G%h�޾O��E^����T�r�x�U/plۣ�q��@.�G���ؘc�����Y��?��{CYBKݾ�{�r=C���u?8�,�ƨ��xX�/"�*v�k�
|��8�+&]]xf�t��<���"�B�~�#��mdk!�Bs\�-�l�����1���~K���@�
�<jU ,v�&
�ڻ�{���y�j?�-�֖o?��@ �-�|��L2T�OKR�<كN�G[�|�p�!XťiV�[z�����ۛ�������E���bG�������M2��?h:���~�DsZ�!��p��"�0^JPgqH7���o���f�� �p��B׎�q�u	}�RYF�z�׭�.��}��hVL�$D��0��J4K$̥4���Ӌ�������g�:_����_����[+m'宬(���"@Qv�w&��b]�V�P���4�cE���7�n���6Ug�匙��o����7���=JƧ�C�L���:��/�������9��w���vQ�sޟ������zH2Ÿ/�tD>]+���n����O2��GVG?��{�]�ݸ���T�/�.~_�o�b:@Rw5��)Q�SƋ�{`�m� �ӛ8� u�[�,!
��Ad�X���?/��q�����l$��X�����mT1���N�p0-�M��:f)V��
���C��	ɥ"���'��C���Ș<������?c�!o��h��^LQ���*�̅�U�o��\�${FQp��=j�Ҩ����1���I�֪%��2s��\֦صg ��VK�ĶS�J��ټD�,�(�%b��BH
~S�E�h��o���؉QoY4i�Ǣ�կ���؇Y�2@޺4-���Ꝕ袹�?z<��L:�����0z=:g�[�v�.�����J�!�:.C�ijV�T<��Lv���~1�k:t�mq(��^~�3d*w:�A �s�6_0�/)�
Ye<���e��X��	���+�'�؜yFN��;?��Y}����z��o�`M���d�_�u_���@��G^�����=ЖX�S�n����]<-�s���A�ϜY��F�j��(�R�q�!D�X~.��@�6q��>�{�Tg�i�M���f	�O+���h��w/�0G�6��_�볿Y��}bsbz����4#3�����h�v(�~���N/(��aL�h�""_mEm��:�.41�G�r�`ud�� 1zF�'?�f�A�=�2W��+���<���2�[:��;X����z;�����A9�:ù25�~���M-P����_q��"�wZ�C �0E" 9�Z����a̺�2�i�4Z�G5����~��ؠC�mo�����*�V!�/�<�-)��POO���r�2����ނ/���6?$��9���޴9O2�l�!�Ǖ�=	jѠY��٢��a:�@�%L7��H�ߏ+�.�}�ƺ����PK*�N��TJ��&R�f��)�����`�-����P��zS ���n���w�����C[X,�S�+*X��8#�S��1�+v�t|p�T�?
���B�A�|IRt�3�����Y�R�I#"�����ݭR�zB�?��Z∬5�j<	��--F=��XMz_����.7��LX1����b��<���}4�4�f�9ZB��e�딲1���Q׵7��e�I.��P����k����V{���%���v�_`�TG���4��R�,c���:![ g��aFl&�X���1m�B��;��g� .ͻ&�?&벧��wb�������	���e'�q�""� uRT^/������د�k@�c����O��#����Q��$3�;�ߔ�p#&�9Z�4��Agd<0@!I�
�"<'�o�Ղ����7�|��܀�����9#�E���4P�g�l��n{�a_��̷B�W���V�Hо�z~�z}Dq�*n�v2խ�@��C�D�7�r �0�npC64��r4��U�L3�$�?"�ǣ!��~�4��;T/ (��Kl��ۨ�EU`*U=qT⢢����9>�6w���B�����}��e��e�L׸[A���j�
$�
�k]C�@l����*�.��������[E�㌾��8�u{~���&q���E3b�����d�&��@sŇ����-���	��(%\���������E2�Q�?5>)
�.𹩻�{�Y6�9[X��?&���|���,��H�,�հGsz��z�h�'q��~��ԥ��ݟV7����r3;CҒ4&z�zb\�^$�)�U5?
�E/��'7�6�:q�Z�o���-���C2�йM8���/_�@�\�3����\k;�^P���4�Hn
�$��O$�yO��Z}$��/��wʰB�Q.��Z�C���F�7��8��u��ݧ�Ux��\���-8{x�f3�S�!�=�w�#)ٶf/j��_�#�a��V	��᲍�{f+�x�Q����	m�V�YUɋS����a\`N@Ԩ�3<YoARx���N�,:?�v�V�w�ۮ����+'al���\� c���M�6���T�4tp��C�f~5��`ͦB:&��"�[B�9|�nsw5e��������Gv4���sq�~wl�K'l\�ЊZB1�3��b�yƬ��N�9���j�uGmpo�/�Y�rWQt�K7�#pʳ���ͧMLd�c;AG� �y��H_�˾��JU�)�i�i�0��m~uK�n��C��S2��<iO��py����ZH��F�!�4:)�H	&ź�P���>��#��έ�)X�lo���]�PU��+�@�A�pF��5(������#e���i��ŀ��~ݲ�[����eI|���7�ƺe�RQ�� c����8(,A3�Jo����ᗳ6:��e��|b�M���2�B�=~H�W$\_�	^��VV�p������ש�M��hǞA������c��ϼz�A�R���c���Wqnl����sG�{����ߦ�Z��.ә�_��$�ӯ&pu�F�.�B˅g�X�G� ��NWG�?y�OI��TC#,ȑ2=N��'�l�2�B��,k^���h�����1���b�^��R���x~�"-#�,�.����u���[���f�T����|+�������B�IZف��l�]LE�|��+'�A������Hq�[7�ID�ٰ���X��~���}�4���,���U�O>�� S��j�8Z��}}�}5���?d������~W�h��a3�Nb��+k�n�J��+)I-8�di�0a�ҏ��%__ (��T��!͏��+ێ�J7�����<��	�!�9���ώ��x�H������[��f�b�X֜Ԙ�p���4�v��Z���0�����і����咷,�u�s��F�,��Jn��me
U���Ͱ����Ö�Gڎ�Dt	��A��s rW����<�i-�s�F������/4f��Xj�>�w,���|���)q��6�������2����֢���$bg�Vu�0�L�x���,M�F]v�>ӓ|`{2�[	J�f��ޙ��͋���{�I�ĝZ.�8��Z��\��}��DC)K1������g�u�����_BV�1���E`Yԇ��]������B��mV��k,}�X0*i�ÔԦI3n��u��sI\�������,U�1��A�!s�iЛ���u8dE�1�w��N��2.ʔ��L#a!4�pQ+5m�䕿F ��b����eLY�荞@%�c
T�x��.y6!�uk=V���%*|�<g�n~?9�[S�43XOŊl�e�L�m}��:c�3s�^�*�M8x]%U��7D����|�	@�ph�ۓi'oki�:��`�~�w�wY��(e��v�>�ބ-+?O�s��F+RD�pU�{Q�,lg����|��"]�]���-���p�nh��T2�\Q���i6_�	���>y�隰 ]L���$�BϸpJ�p�)l�D}}�@cs�'�V��kv7e��:��c���g��Q���d�AV~a�I0d�+��v�h����}ſ3��S����k8�!m�+�a�N�0!@���B��~|zcy��bO�g�j�R3kŚ����6�ڧ�ͧ<�*�z)"�ū�yQ���|#a<�o!.i�O ��6�6de@���oN�����.��9jLǛo��@fҎ�w���m{
�\�?�o�e������"�i�2���MG��f���)~3�QG�6�.Cbכ�6I$y���%�m.R�d��9o��]\�Vv���f��(NF7��;�1� �d�/�����r��hI�y��%deN�����UޛC����%������ג$0�9���l��0[�������H�	_��wLe�����B�)q�-	�墠Iյ�<:�Z�`jn�~��6���4� �O��o������e�� �н�8��� OFtVU��ɦ���,�2�h��+�	��X���ZS��Pe�z.GϓW�5*k���=��'���|��ڠ0��顱m2撋��=qT�Ț�W� ���)Y*c�>gIy��V��/�����Ӂ�3���/~"ax'��E�Tv�/jc���o��v�:"oe.Kw���/� ��@��O� ��)�ߪs�!�� ���3@U��>������^Z�z��#8[�̰�����ܘR�J�ћ������U���&ӻ�
{&��[
����*$Z�Þ#^ ᝉ�z�2�8�6��Q�y�:L���n�@U��b�^?��b����\x`��<�F����dv���5��qx[�U������ҁ��앤k����+��djȫ�o�dK�ED�([(��U"�����J�Wۥ)���gd�ZG�=��_R�Ё�5�UU��8ЀY�����/Lb`�I+|��
\�kc9t#��������%�3r�^fm���-��?���PT��w�!MH�4\�Ѿ�}�L#��:��&� ��%�O C^m���)�wד~�c'F��w���;�� i�X����^N.X��S�+[���{8Z��8��iZ�\�R�C��HvX�E���`���_�/����PG�S�:�GwtU�0���s�DFCFڦywD����sl�1G�Y&��)#����+��Ç��u0I�ew1nM�:j�K��_���t��<Ic�c<�̦��Z�^������&�ġd���Vs�dp��Wf��50hU���X����rꪊ��(����ʔ��P��2x�
ə�󡢎08��	��㊹L���@P��yKrTٕmz��Ġ��g-�#�l�Ͱ"�;8��
Z����`��P�J8hX!�U�}�@��$:Z�}d�1��WI�B�����'�t�{�	���$xX�x�*y7Y�\=F�CÝ��ý�����d�}�fq�v]�A4ՌB)?�"ͳ�����f����	��3N?n�D#^9�����_�[�_���I�#��.�ѓ��C��kM0{�l�!��A��dM�L �7�c��9�Q�#�
��4�>�B y�$d��ƻ�7E���f�V�1���}��j�Uq��N�X��AqW)j��2����U����0�5G��,`�ݟvv	�5eȽ��N���#�~?�gaP���n���g7U�:C�͛G2�ߌ�J��h���fp���1��%
�!�@ �Po׺3Z�Un�r��c]����D�|{�gͤ�y?U[^b_@s��۝S����F5w8�Q����t#C��%$�
�5��ມ�� �:��2|6!LL'���tW!!�{^׫��s��>2d�+�x'i3@��ݖ��<y�6�b�l�S3R�W�=����8:����VC!#ʲ��`<�͈T�L��}7�M	�@xJ�c㍢�^b8ј�ɪQ�Z��%u�tT�T�V�霝��~�)��R����S`��ƍ�|���|��t���	�1l� �u�QmZ����n���uC}ԓ֓�@��<��h�+&ȯ�N��,��ZS��l`¶�d۱����r1v��ۮ�tv���d��iTB�S�
^K�k'R�&���=����)��Jz���/�[ّzA҈�O\_�98����׉��5��BPȏbr�i������JQ|�������9��+�6�� ��S+^�A�����׃��>�4�1w/�(~堛Q$�ci�G,�m4d�7��L�V�vYa*�����|�OX��)�2�^�J�dȞ^;"��~�!;��8��Cev��e�ߩ����_�W${@p��.yKaCZ�I�=�8�x��Z��Я��6v?�<8t
,��j�~Y�ڟ8�#l�U�ٓVZ�f�#2˲=�����t{N��s}.L�,�|�L6�{Ik��C����d�%N�aj�����KV��9�ߜ��q�f��s]�k1�s�u���W���	<Ϗ5�YuD�_�|9���ȏ�#Py��S7?���g=u�V��R��_l�h=-�X��Oc���ʑ��Ep�q�ln~��ȿ��ˌ�C�D�l�ߦ	�	��s��~ 5��响�`r���J�M���$RK����}��� -�5�v� ��*wD��-PO�r�*eom[�`�e���)�e��#ُ����8Ӣ��M�ͩK~@��*X�E�#��f-9x�;$P.��y���o��0������W洮�ʌa&�8 �86�5ms��Y6���I��_)hS�K^��n�zKz��Q��Á�\�Y��;���/~`W��JV�¼)�(]Lm��YYV�����]B��h�R=|��G�'��.��ꄸ�b��N��M��@�ۣ4T�Bqk����r�us��V=�3~��pߩS��j:c剃Ģ���>bq³���������H%@��KM$�Ck@�O.� �[Ǫ�}�=G�*�����Dn�ɥ]���i������[�-�����m�C�y���OP�XuQՎ0�M�8�,8�7G�<�5.����d6��7_�W���#�1�VÚ�B��������B�i���� �>�4��T_�x=�
Y�k]�v����I�M��🎅_���]y9�L���.�K�{�]�W*�ǧd��A�Ky�褘ё����՛�7l�ӂ���X�j䱪�$6���O؉q���*��~^���w�?��M_�F�-E�Тƃ�n�ҺZx�'`p�je�# ���u�����8��*_��7t����S��!uб�3�5v=�C^gL��Wm���c��܆�Yi��<�2p�6�԰M��;�o8�4���t�Ń�m�)V��tA��#{�����(
;��SM�W6��TTv,�<h���Y.3[��<���9<sh�;I��#���[q�.&��[���o��@U�P��m$�1}�B��M��$�C'�zU�bЫ�Ӭ*�B��C��q�u@[?���z��[.���~�+&�]� �U�8�U5*�B��Q�k�D��ؙ>���������vР0 ��O
�2+hZ���nes/�����:��e���ၺ���1���fy+��<�3�c�#%�U�6�8�EN@�v�������o�=_��C*�b����Lq�!�И�آ�r�	�]/��&��[�"-�T�V�ڈ����gD�n�2�nN�(=S`R@0
�t��3ږ��b���]�h�%��!J;����D%^�\(��
2�Z_Rب{M|)b��\X�J�$���;<����������,+E�
ܮzSf�|*we���I.v���E��ZA5`��������T�o�o���3��J����/���,�Ȓ5���"�M$�CI_�A�op�C��c�6�>��t��R��9��P.���
W+�=ި�j-X_O�fѻ����B�2e��*P����/(����#Ŕu�Opy:���à ��s����� ���mHRpk���ƶY��%t��C�>�瘰�[p�%��\����XE� �bz����y�ݭu����pr�}F�4��� �3�ݰ�����v�Wя�^1�i�������LV���fڃ�� �9���Y�B��.*�TR�Ua�]�����.?J��(�yz̎HK��=@�[�/�U!��|n��D�' z��M���ۄv�Б.�/�R�R}��!Y8F�TKGaa�S�+hI��p��2;�Aw8���C)g�ޒQ���5���8�K��WtPdiʴ3�a4(�)Z�5�uݚ#�����W@���3�Xi��صW�����%YjF��Zv�)^{E�5���5`���,8�Y�G( �$��g"�ڮ����I2� ��+uMU34Y�Q�t�q��&��ru�ʾ�t�IRC-��}7!�W`Cγ���� c�MU�n�P4��l�U2 �XR��br9�αzL ���f|`���n�����{��A�u�`��ei�g3X��D�rjh��h��T�AK�ߌ~-�-3�X�X�G32\wJ��{�Q��Ot��?�~��ѹ����_I���x�L�aԫ=��E�p�c�xf*`z6�B������60�fY�3e��i�]�ðK�\�ӻ~	g���
*u�$l3Okۤ V��z齗����.��2�R(�K�t֞5�M�o�]���@��H��^0Z�(Ɲ��\��\�2��ѕb7�ڢ]G�V�P"�䇞Ϸ�K�A�R4[����������qX�������<��jl�w��k
y�Z����<�?����q�,��9>�W#{�d�أM1�+�h���UM
%/��b�D}+�A�t)��R�f�	�|�g�Xױ&�Y���{�!6��Ǆ;�#��2@I@��0Q�PS�~/X�>�r6S���H�V`�T|���5"a�����E��Ͳs�J?	$$ԯ�v#��q��Zn
í
�?�����H�dD�;�ut& eԛ2�ďmв[raUY���ӐC��U���f���҅��r���5� ��߻e�a ]��ŎyX?��W ��
!��:�v������W��[�4`ٱ��l)K�_�Uj�
���6�1���VXfe�c�EJv/�t��g9�:Ć~�2��0����FC��H@�?W�u4#ON�#$�����X�G3Pr���ME����~�(���V�)h�)x ߺd����8�������*��]�h�=��T��]�_uK�N��������	ϛ���*î��&�h@L�P}tC�x�<��ʇQ8��q$>ЇA�Zӌ���v����Fz�ޑ�᭧�4���N=D�=�P��80�.O�Bk��yk,���H	9K�9�4lT�c���|��*	o�I���YR�U�a��ѓŕ����Α��}��'+>R�ɇ�r�{��G���-�TC�W���Q���o>zxn[�F�$����Ӟ�QE�~�cx�� �ܩ����|3�KOݢz�-0i':(�iD�	�H�8�1��ua�D��u�+z"��9x؏Ѐ-�>
"�vg��#il���U#�s@�Z=���ة�L	�,9�fd!j�G4���R�pO_���ol����֛*��f��u�^L'�%���.��6Z�E9���\�nLk,\����b�I%�E�>pr̍~���k#�
VY ?hvg��O��"��y���&��mo�aϏH�e��cV0�Y�`�K�9���L��9WT� 8�5Ç�{[אQ��j)Oӎ�6{���1i��b=tY�%&�@obQ'�d��נ]��Y��xY�3��/[����uO�'�F�`DQ���7�xC`�h���/=z�R��o��8I���NY��1ܽ�6tam��b�y!��'���:|�Ω�\�eikh���6��lL�;;��z���aXɣ>�z���P槏J����%�$*���%�n/܍�8 ?�Ȗ��U�Vk�U$]�o�*���@�v���ly"=����P�#+lٜr�	άB�Z����̘�{]x��[���`�$�����% P�J�>m�߈�p{oҀ F`�#�=8�����{~΁��;�F�pEc�L���c�/��(��թTi�H9��J�>/�b²�]�;>�K`��	>Z���+{��d^��%r��X��7�!5�=ѧ��ì�V�n{q��C�pS�6Z���jR���bo:�).F0��N����Q��������{�9`|ַ��]w澦ι��$��$vt.?�S��7��fWom�eTvUkQ�r�2�}�:2y�߫�Ҕ�9�I���K��LS�~2����-Vu�4��2T-"���p!��y�:q��ZnK۾��-%o;��lu�G\���i��8���� sB���c���#:�1��Q�÷���8���%E�(5�H��� D�*��B<�:cc�I�ac��'�:���` �:H���i�*S(���5Ǝݸbt�O[5La6���sSU�%/e���%��ݢ��A^) q��U��Ȑ��Ym�%Q�FLR>#=!�=�{7�Y��"�@8KB��ً�s�i%ͧ �o|Q�R���|}
�}�l_io��#\_L-N�G}|벚�]��o��BU �����ώ7,�	�]��j��@1�?G߅��;i_��;�F��j�s���	�!�J]�A�Z�3��&���9$:�Í�����0?{�`�,�nj�׫{�p�E�����lY��.�O�������cSڠ0=���vꧼm熿�=@p\k�t���ߧf��S	���S�1ۈЖD���'�P�O�D�Q|q�߯.1��:��i��<!T��8��.ɵ_�t&㰲��7η�k��Ih� ���l��z�,�P�*�l	b��A�{gO���z�9*�3�d�(��Cgg8�,����[�Eׯ�'Jtn��P�o|v�u�����ć�3;��~�o~^Q2N�5�ʱ���be��!5�����U,^�3�6F+�GkA����5�ʨ���Zu�»Wpu�*�Ĉ1{��I�率wZGD�(7N�e���e��yX6
�q��vf�w��NQR}}�Di�����1#�n2��U��G&���$�s�����)���#���\;f��g�i|~�ރ��ji��H�{��[=8��oXމ�!�,)9�F�n��M�:�������|4�$���e�-�i{L+��v�]��G��tV�t�,�v�#Lw�+M�ډ�2�>]�\5^>��4\�w͖'h�٨��_Å��t`O[N����®t+�f}*�:�ͼ�d3��3�h�q#|L��R��*ȡ�E�+A �󍽯�BI�~�[\�Z�(y����7@�k�
.�6J�S�%�g�UJ%���%��]�p?L&��gE�h?G�Z��ڪ�B���yy�8�U��H |��S!�N�w�IU�F%,��>h,�2�Ѯ��S�A�V��LW� ̮a�	o/4�B�m�1��c9�V� du��Rв
���<¡�Fd\�a��.����l��Iq�9�gN�b5)��v�[�9�*(����1pu�z����X�d0�9P��Q5�W7ϰ8�� �ۢ��q���A���"�7�B���Ps�a����s#?��D�]�*�[�$�-O� �ݡ�F`��D�B��rw��NX�Q>%Z���	s�w�+U9�44٨�9?�f�qv�,�n�bwK��l��[��MP��3}9�R!�st�v�Ҏ ���L�<�V\��"�lT��kHf�V�>�R�+��kuTF%�&���/����~z����sh�Mr��/r�'��ܗ��
���D@����cYT.���o�u���^�6��x�LTy��1���@�/:��<`����^�e,�����V�q�Rj)���m�VW(5�/�GS�k���ƛ%����	�̀�Ք�а)�>]�BJ}�b٩>��74�����_�+q޵�CYR�ܶllz���|K�����5����Z��k�2
�U��A�m��U{	��}F���ٌ~4y�Ӽ��"}"�.ёFESS��kL�l�χ����y�P׺��^ga��ZI��:w���=�o�������WrY+�vE���R�&O�����U���봢��O0�� CV]�l��^&E4�Js7T�tzX�a��w{o����6�ϴ����� \�-z
�
��&����������I �q������No������W�TH_Oٖ	6�n�U'���[��H���[4�	��-gJJ*����0Z;6��������J�],�2��`z@,M�>B)�1}�h��}��05G�5�+R�3��]
n�N�3|r�"����qug�@�ɮ�>ک��2n�O8P��5�/��1j4Ye��;E�����T��s��iu�a����/L��G��e��Eܵs�k8���~U)��0��Aj>��J�Bk�V�������kK�>C���6�D�Lz�O�;�����H�\8&�{��TE��,'[�S p"�?�@J�t�쀯|t5��-X̶��3��fU�ٖm��.Q��q_e�ey�Սِl�ap�c��3�Q�R�1��a71��^�O����oe��'Ȣ�.��jCU<$Ɨ���X�^/ 9�\�����ʃg��!������X��*���A�:����\��w�������.��籦~X�&��f$n�w���U̧���x[.��w��"�{�y����j�����q� 0�jW��c4�a�,��"����v�X�zVR�����F��{���Q���ŷ��yj:M~�VF2�����SnBaU����wݯ��"�*�*���M]�G9�j����U%1y�=׬�>���D}i5�|�e�bP7Ғ�N����y��u@���b�vy�O�� �BOc�|,V[��mD+jSmUa�鼸��**�����@�k�4m���^��磤��=kb2�Z�ö��������R{V����~�ҫ3e:C3V�X8K����	L>�q�wKX��S�����T������T�du�A�ci�/�P5��q��gY%�K��x#␫�`�fr���y��z�bP�0���1� ��!c�^t�*	� �k����ݨ�o���3�ė}����ND�)�A�|\� �����-ﺸ�cR��=Dv����'ЊC��Qb�i�������eӆ��J]�da�ۅE/*2ԇ���񱽋1?f��~�z�y��E �\�\8ʭ��}M�/C��]C�9���{���a	M4���OE��}��q�*�.��a
��6rSd�O���;��~L0-y��]��ϼcȶ{7>6�4����,�QD�oV԰�Ԇ$�q�Ԅ����eIȆ)"$�ʢL�щi�:��I��A�h����m?L�=��苌�x	������Y/(N̰���]*=�Kc-,+P�pU��`�aj$|��%���t�,EM�R���>�f��N��^ME��b�D~P���\��$��y�jS�o���s��l�9-�\���W���g����Ϙr�߫�܀@��`��r��8��M��`]��I��v���v�H���>