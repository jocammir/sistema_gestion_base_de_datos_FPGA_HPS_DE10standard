��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��ᕫ��H��gq�f}���+����c��0�7�*�y�HXH�+��Y�Ar�#�<�k���bu�-��.���O�;����b���7pE+�������v@��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T幭xX��8�hG��kr��'�n�IK�v3�[B���fP�e�q���7V�&����J��v�(� ��n^�ӄ�`� S��JK��W�|�	�bL�Ԡu�%��x��@:՝v�����E�R+� ٖ�;�W�_��h>{�J{��O�xO�D���Ab���҉N��ʖ�MB����^�����y�'��b�|�����������V�V����/�"�b�m�sOf� t~ь�
��a�&�LԾ@�C4�6H\3�[?tctrs�9�|��;I3G��op/h���ؑ;�d0����4^����IV͘P�*
��G���%�:�*Ը.p� G�)#�7�Z����j���%�b��5?�
�QoX��ac�,��2������N�'�fDc_�PғJ���iP4����W���SA���q?!�oI��X����a��a.0%Gom������Ã(Q�^ �{S��>,�`!�@zQ���$b�Ǟ_s�����=��G�"ßW���.!���(4�M��Sǽ���6\o����>�:�Ҧ�(��4�J�!���&��a�^���m�������fS7"�pk-��s�
��v8��ѭ�6
h��]^�י*ȼ����KDMdJc:@�^��O|�����t%�v���u$�s-��>�#��O8'}�e-a٠Nt�� ��4l�� ��t&���@�6,���V�hS��7��2��	��:�J7�%X��r�B�c�]�P��H <�rM��
\�g>Rο�J̎����~c���U�MI�����{/L	�u|%�&�Sc�T{v��+�	Ɲ�>U��_�q{:G��C�J�|�������t�ʸ�$����;��˶�,���^��a7V�ܱK/I�e��ԆF�"�����$����ʹ���%���XA{Q~PMl�gv�$�b��4��H`���<��Q	�*I%�1	z)���N����T��_���{����B8-�r+p��륇_�B���	C�
�&�PR��x���'��1����9��C���x̻�Q�~��c����j"�m&��B�~i3�ѕV@O{ogQ͟�p&��]!A5���@31���3؎�X}B���9/�C�{"C[t³[�r����ӛcWWP8��C�c���.�/�����?K2����l��H?���.�|B��6����Ĕ5�;��J)����$��6�����6%�_#0E��i��~N�H�y��<+B�ja�{�H���������h��lW8ޛR�Yɣ5F���^�/&?�`{x>��z�ѭꙒ�իu��%fi���i�`��^%��TG��
��9:���N(��m�Y��[x�vb2��qӤ�R;6^3��M{�ה�1BRQvP�yI�7݈�Ȣ@sI��R_H����_Z�U��[9B�s���J������`|x;���%\!���뱦��6��v_�S���;A�L��K�y���	����+D��j�ҽ^%s����+:`(W1��sTy"�بxJ��E�yＨS�Y��������!?�%jJ��PS��-u�� ���u���6��qN)�t��a��:A�{�L�>��jk{Un�hWf����CE�jpR��e��
t.�ɶ�H��ؐD���&KR[P����CYQʂ�l'���I��JQ{G�j@0��"RPfuߤ�2rE�Nh�e��RSM�Hb��/H�J�<�Soڍv���a)x_9
b��싫Za��ԩ+eu��z�k�|�ѷ	@�{*�R����6fW_��I	���1��T�8�S6O��S``���X��B=5�{�OM잛�1���x� ��S����&O�qҊ��bpF���[��I)�%6�{�r�3��h5�<��n'�R{$q���%-Μ�ҳ�_Ӹp����Xv�i���Aw��&���{�*���9��Vɂ�>�1�g�T���;���2 .š�jr�����-�ԣx4�L�:��߳���.�L��zꩄ���G��$�8������K��l�ܔ$![+J���O掶_Q�L���X�rQ�.u��$��>e9
u5:䟌a(�ƾ�{eY헡?P�C��df��q�<�&���ҷN:'�l'�xX�!��;Ç��@��N��?Z�C��?��ٹ!8��*�~V)��y�ta�Ş��vT7�S��ZT��,>j򻾿��L�Z��؃/^c���K;�p%��Ho"w������DO�=d2�S���m��c�\"�a�l
\�^�Jn�k"�!�q����
�q�sb�Υg8M+�
A��$"����	w���jT���j3�d��8ñ��{�#��6�*n�n��2{� ��p�+�ةP�ܢ}�>�U��̰e�FD�;�����4��$]��1�#�Q�.8B���j�S��#��b2�\M�{Mɗk;�6:��H`�9�N����	"��cq��A��f�����0��#;ʪ&�tK5�Q���:�f+4Ť�#��?(Z�D��j,9�z���A-/zD� �y�e�lOx ��D@�p��>dl�c�JXp{><Mw��n_�|�3�}Ҽ �{2�BLDL^��|9���.}|�^x!�)5��0��Z�[�P��Bo�Y���ԾN�ű\�zP��1��Ԛ���s��������4�ꁟr����B�C>��N�.*b�X����R���E�����
�(����J��N���v���N� ���f[�m�e�m���.��]r��Z�릸/��g�NދXN ̀�I��N˵���[��3��R��:��`�6~`�k�j�Sm ��R���P̻w�0����*�M�F)4r̛
��E�����b$���Y���|���7Y.�ȝL.�WJ�����8��O�^�D1׺�:��ف���}��͡g��ƛv��/���@=��60s�N��b�;~��~�ӱ�@x,�rx�_�lG23 G���%ic���gi�8���r��Pqݳк�#*�!�1��2׸c8���F�&�g��w�KP%�mn�[Py�v��&Ghc��xV����gX����_Yc�MnJ��#+!���nG/^>Y�5�6��M��' :�H1���%�j��������1�eE��U7^�M�p.�_�q6~��쇦��*�}9�#�1���ǡe��Miv��8dJ�p�q�Pā�Yn�`}Z�ם9�s�;�U��
�!�V2�s�1�a?Qx��<�%Q�� ر�w����/�P<t��#�Nl3>S]�C��°��J�j���yqqP����!���:>zC)��D���~`n���w*Zq�Ō{v�Flmh䅋AN �q�1�F���5��n�xK6R��gEG\aV*���s!`�s"�]�Z
����`l�İ�/q����AGZI۷�dW��v�>i�8<d�u����ڢ�N��@�	�т����wa^g��o����h?+������Zx<.s�Q�ͩ�Y�q�
��]�EA���I	�������`0��lX�;�l���X���V��W[�A3"���/�g>�,[�gP�J�Gd��d@Y�"K4͍y[$U�g�G7@h)�IK%;*�)8�Bh��8m���gYq�=���DG-!~R8x�8�;��?��C����SPJ�Яc���(��Ӄ#x����MS�j7N"~6������oo�P�Z�!�n~LDv�Y�I����ԕu��z����%�7���@%�g��.��Wq�MQ��C�ײBߊ>*�+"A�A�
�F�ϊ�"���VVq�bNLX��{h �x�{_Ԅ�7s�/g�И��Ѹ�IE�9Oe�3o�I���H��ӮzmVl�nW�0Ijm%��P��6���ܙ�'�&�({Ygy����=2�Z4JJ1 �mle\O�&�"]�HA�5,��Ϝ�[�^�I��PL�[H;��q�>7�g>�)�,V	�i�ܣ�<��ma�7�]��$�b�S~.��
�L�?N�_���LE�T���0@�}�!M�]�V��^���,2�&�����!�J��,�(w��v�zj��VC������^<���� #�Lɒ�f�w�Wx��^�p����9�T�|����W�w�ˍ�n��tEnr��u1��]~c^w�ֳ6��u���ڲF�nW�n<�rh:�L��#1K��Z�%��s���LN�Z�[�[��"���iNK1G��5�pv�?�Z�-#�E�t�*�3�WN�u5ڃ�A�
jM�����3{{(��a۬�= �P��8;7�b)����03����M��;�V�K�B�o&M��&#���[kƻcׯI��m_.^u$ʈc��l�Sƕ�Xku��Gk�7o-13��� �)[�����H�KM������?�N,�d�����X�cBc�{���e.#t��ሇŢ�������!,���HTx墏h��'qS42?��*F���e��9�G�>Q;}�ON����� �2�叩��4s�y��k�t�S���F�Nɑ#��i4��j.����oJQ��U
u���B�H]Pq�[q�Aַ�0�`F����B�5J�D�JY񖡈�� ��aPj�K���v��\��X�İ!�F�̹&^�U���͘�Y\MN����W���+�BшyW]����Wk<Ja���f���}�R�L�l|��#�A�Xl5����o߮vN�.�[��M#�4$�G�1�s�(2קы56�}a�U����3$�ή�8@�~G+pƔe�M��O����z�
�,jeЛ�'9M9��5�)OA�w��r�/�ط@{l�?����=�� �N�5��C��9>r�~@������C|?��/?#ˋ��V>L�n<H����<�ų�Q����*���5�
;��*Fו �5��������7 ��Ώ�`ӿm��i-���sf�|�c?&������Vx9��r��I�'�����x6�C.*a�
�|���Ԩwˤ�kʀd��~�
!{��ﴵ���Il+%��þ���CO�����;�x�_���]���H5�nͮ2/ȑ��U@�m=7�(���)�[f.��(��%�{q��>*t�LD��ޒ.�&�pR����~݇���{�X��/2^��)���u�/F����A��
t;*"�
b͑4?O[���𛽿X��J<��Yt_�({��(�d�OL5K�{��h�!Y�J[=��@�VX�y��{�jT��`���f�=��!1�r8�I��W7AC'r���1��.;Ԝe
�b�z�+�)�q��$�n��"c돮��pۗ�0�%<k��[T~k����INŐJ�A�~�eI�����Gv�����Z���ȋ���D��Φfh_�ޓjؚ��x0c�6�5v��R\ W��P���z�i4��	�Up(ە���(�=	>œ
�m���@��{#�q�+�����v�4ą�3�N���;ڷ��#��f��G�@�)���B6�s[t��}�|���G$y���0�z�8���>��ڹzǐ���j���|h10�2�{��B~���TcB��w���t��BG�+�D���F�Ѓ�U���k�Ҵ�.WW��̴u�����;E1��~����xɏ�ɝ�W6:����Wt�aս*0gsD��ZB-�n��N��7U>��z!p=�R�?$�UK�q�h�RdB�ג�o�6Wb0:�\�������Y�q3!�eݮ��62xo:�ۥ泿3��)�ɳ���S~G]cJ���<���1������f��U��^3{ߡ<%[/�� ��UD��Oh.y�IO0����d!�H)�
�V7X=8�.������M��i~\��&��?i�q����._�ұ�7	^L����J� ��V���e������I��7��P�Ӄ�@z���[��(�]����R��ֲgM��Vb��
t6����]U�Y�Y?;,�fQ(/[IO���h��)��H�(�C,b��~����f˓*X�SP7�p����BCdşwj��:��B�@�K�b��~g�a+�R�;�)C������ܜ��*�эa��@�I�5�T� �K����	�\����4��
>
]��P�A�&�0��|�8��,R����@�##4`Wr�
T���g3�g���D���8�J�Fe��݅��"#D�f�"��` �7�/u�lT�Oh�?�c�ee�����G���L�!�_������ǅ�fW��}��$���c��_ohW�_DP|�����o���u����x��5�nM�+~��O땮�(:c��#q���[Ŗ����\��I,x���(�V-�*O�W�F/(R�_�Ӯ�K�<�4b��n�u�!�j���՝{�����2�\�RF(�OE�������,���2���_y��Ic2�^FۭVy��3��(wa68v\'�l����oR�8-Q����֑OD0�_�*���@'\��/>�j0O�\<t��T/��	�5���B�^Jw,��m�Y���7�Nꇁ�>�7��������,��#��c�MY6Fi�.�y�h;g@��ǝP���K���uZ�{�U*<��
ǵ�'�����BB�y׎�Y/������j���\p&��h�֙x�������U�ڦ�X��\���na�?���3;��HMQ��7��Y艸r���Ru=�6��d��|	��xȼ�I��Y�S����٘�ROf�&F.sN�)�JX		�=nOɡ{����`"��`\�YE�Ŝ��9��W�Y/��Ο��>�e�[#�ی��5�RW w5%^{��V��q���m��9�n�x*o�,��	�i*���b����l�8A{/	+�0~��L2>$�5�&�d4�MB4�W�=�����Ʈ�=F�
h^���o���"���f�WxP���t�m��=��"Ea�E�:�gg	G�i>�����lz�D��{�3:�b�v�:i�h�]`"a�C��;�f���b�&$�ʮ>��!'�5_���v�@�4�'�"��s�'AJzt@�N�U��خ�]G�T-�P����t�WVɢO��=�� ���-o#Q�w�N��O��`�3e��-R�Αy|Ȅ�L�M�v>7��K��2!~�yݟ�)U�ϩy�v�l!�/|�Ǿ�Ƈt��I��n��-���p<���%T�t8,�. Pt���,h=�Vk��2�ы�!A��ѧ���^�����@�����f���2})�qsl��0��0�бsT������+�e(�4��Mo�l5�/�G[l�I��*�
>ݡYNYN��̰�m����D�X��T�8��E�7����}rA�-�z$Y#���\`�Epv�Q��
�8���7y��rk������*�"S{(e�2`x9�*���aC@�	�c6�q��s�\�Y��7{����đA��Â��,����E탥q\P��T��A�F����H5�G������rH�[��w+ɷ�S�zjB\`[~�������к�i@��gneHٍr����%%��V�����ڶ����>�K�DV�z�C��s����$H�7��7����e��$�p�����.VJ��ً���C�x�'Wdx�B�R0�L�\�X�����O��	�j�X%�s �C�-lg|�h�c��~oY?���Ӷ����%)�h�����˯�,B�,�
����T��m4�����dR*���sxW �H{W>��qo�>��St�3�����^�C��CK2���D3<�@%�:��\*`�>�YJ}N�bI��IxO�_=Uc�Q(Lym���e�Hmpw�a1}��{�u��#:�]�7!�tr;s����1�{R�s�#���N��'}��H��n9�p��m	 �3��?';w�֟��	J�8�5ߙd\���r�R�Of!!��!���*[Tr��{D �`Ld�&V�/�5ou� ��/��퀀��G�#���w/�;����V��Wɉ��&��/��ρ�L�Lo3��[@�q����BRk)D!iT�)��1D�,�B5ô�Ns����Y�Z�x�f����G��St[�a�4⬜������ra�[�WE�Q2%��(�q��0�/��W��w��	ޚ|�7{�Ez7l����㱵�IYl�f
"� �A�a���������u���b�t��	�k�Þ�6t���|��C7TD���B6�����	��o��x����#��a���BU$�L����$r�/eB1��S�ieuf[�[7��՚�Q�@S/L�QPB�_�8���I�L)g6b�O�cj�޷[$lܶ��l��i�N=�6�$,��V^s�Xv�:u����[�f�&$���1�zi<$��J��d�=�Xl���2�tfݷj�����|C����R*�e�a����x�%�=H��܌GwI����~�*F>]��0��U��!����#<U��'�z����{���Н��Z�kpJ����Xw����P}�����ԙȮ�����ӈ�#�@G/�_w*.̊����2�k���R$���Nh+q?�ɜ�t�k�]1���ٳ�JT�J	u]����!Z)�-�#�cTP~V��[juw�y���֛|�s �Ā���ɤ)�{�^���V��%n�\O(PHz�K��%YH�!���<�ř���a��߀6���v��h��DU?��+�k���ו$�Wa����LA[!�U�H<w��zc�+@-�^����9�yqP-!��e1�@A��f�����c*-Q"*������k�=[�ې8+�0�Sq)� �����w�H*c����YU�Q�4��7W1��������/����M�ۓ�ξ\*OBz���>��9�x��_$z���j��fCg��2J
��y�2҃V-)|�뜰+~ɝu�ƨ(�i0k�g���y���U~�ƘIo�-��|�R�ɧ390����/
�$�K���K��%�9i`�/���%��>���WQ��G����<�����Vk�1P�%���,�@�0 EH�5yE�E��(���y��I'���Z5��RJq������}�m w*�È�oJ�����ƹ�0���&<�q����O�k�  �׊�?D؊Y�v�>Cߌ�:$j
n�?�j$��9A'�Ա���?�����>��d�|���V\Z�����A��ﺩ�o9Qʞ���z���k�jOw7��"������wB9�wi�����g·���3S�c�;|��-gc��+,Q�)���`.!f~��H���
1�H sn�~�����#[a�O;E�/b�>��B���5��9ҌT��ϙ,CTI*v4G+�`�Ӕ���)h�h�I�">�Ő��˅�J6�dˤ��4�{���4Q�|��?��E7+V�S䁝�jM+�2l� ���j�[5����{���c��D����P��2�+>Е,��O����\�� nyr�ŝf3˧NU@�w�A[��J���Fu�����܂0IR�"�����R^�V^y�q���[��c�����+I��hە �/}P���ǎd���4�*o�i�Vl����,^H��
�>��I;�}��m��]^3蓟4���g0��"Lq�{�9�tԀN��b���ѩ�̨�w��(�������4�q�����W�Z1:�z�6�r"©gOh�hm=ݔ_�u1��>n�;�a��ׯh�M
��@�騷��t[y0����F.�Q?��̝����F->Mt�ҭ��/���M�fn���%�^&a�F�v�]6�Y��./��ߓ�?�+2�©IJ��8/���N�B��h�<�h����+ߺ�����u�]P�H����ǣ���P`t���f_ؖ�{M���Z?�Ҩ�T�?Y)^ �}|Cm��*3+x�<k�X����/]
P���n�����g������`"�Q�M��L2����31Ɵ(o�!2aCq3,��Vg1�γ��(g�0Va���|{ Ħ�������@8]����z��)�=%�|I�w�4���\s֭��}�h牠�@/P���U�w�IU�$ �!{8�'Q�i�` *ٍ��GH@����1ڧ�½P�D��_)���&���6�r�����\���M�
2�e@d3��sH^%K%�@u&N�=Pe����ծ���ɖr���l��
tӋ��?�� U��_#y]E���e�|x��p~��xdмm��"�s������y��'���P�9-X@��\� �̫$�$�?��ٿ3>$���3�@���+�h?쒶����d�8�@,"�~�!V����e*�r����v�����oK*	}TBc�L �0#�2�%h�ac2����3���2���� �%3�Y}��l5���Ŷ��f�΅y�tA�@�T�V>�v�5x8�D��JJ��_��E"��Q�9�.y��"�8�x�V��Ǐ��4�b��S������Gmb�~�1�ve7�'/�54%��:if�m������3�F>!��'���Τ�7�r?���JƵ���0�1n�PÚ��L\�P�W���e�]��:�Rz�̯��U)if�/�}cE��#�3�t �1\"�v�ި������<3�1z�o��l*��I���a|�ft*�ZP\d��l��:0���3q�l��.@���Kr9�ս��>yb��	�.]8�\�ug��Y�ч�u<�	�����`v�q�M���EP�$�A_7L6ά�ԏ�4����̨/�S��pD�bѷX9���ㆣc��tO�b3l�F�7��G�jX(O)c�d�Ӳ�ҝA���Z,c�'�4�x��M�c����b��Q�Q�&C.��|WI�G\�X�e  N�w;�{@Pw��h`�lI�vR�9܎��t�o?h�mŎC9ϓ;�ł��B�g���#��J' �����F��O�J��6a��rt��S�Q���e}��b3X\Wf�VZ�ؑ�3��::Z