��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��ᕫ��H��gq�f}���+����c��0�7�*�y�HXH�+��Y�Ar�#�<�k���bu�-��.���O�;����b���7pE+�������v@��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T��F#YTĞ�ج�Vu��#/R,�DD\�o�+���6F����u7�7�JTY���!T�K��?��:ۣ�����y75$p53:n�<��|� a��筗��&oS�������"d�0w���9pݱ4��l]Lo}ڏGS�Z+.H�b�|`\��+V��~U!����c��b'I=o9��ýn��Q {\��0�W=��r���d��2�'ų	�u�<���3|@��e_�YC>��3�|��`r�1(`8��an�^��1��؅ˇ�h�0`F�:bn\��mp�<LA|Df���v}.��������%~��@��?{�s:���i���E����Ò�����<�fD99�,4O���||�~�J#���U<���ؑ,��4����1�j;Brf�~���^���"�%a
1	���c#m/ɓgn���n=�J����Ξ_�^�/H���>L8b]�9�w�)*%B�ȱ{<�y
t@/���A��c�@G�T�y��A6�0	���-T��6�KO�jFZF>���v�Ș%�H���N1%�۬��΋0��6w�Ic� �d�}��ڲOq��P��52�E�_d:�����ݴ�Ts&��ʰ��}�}Y�� B&�2y\��v��y�If��3y�9�� ��L)�M*r~��5����PT�^�ہǼDr��)�q_�0����M7�$R�Q�Ί[1��
����"�!�M��C̈D���n�hw
����^���L⟫�\\�2T�W�J��멯�6v8�������QB>���$�_�[f��6�հ�p�O���9����(���=+��������<���v����b���X��ȥ������Bם?�h2����#Ft�l��W�N��[�SM'6�a5g �= �῔Z�?�kZ�)��?��6]D�䘹Q�k܈�v�Y6�Aހ���-I��b2v0�Դ�f��!^���i��].��~������
|�$�!X���w��v��n-���Fe�6��%y�6�cx�Ɂ�y����Ě��9*}�|��g��������"��R!�	���C�3��Y��� �4���5�� \na=�nu8�����?E�ظi"����ue�T��í���<�Y��}$�5+l�3��r�[^�fz�Dy�RVg�j`EvUC�-�ʀА����\��N��q��oz�#�C�GM���e��И�A^^k��L��y����wa��J (�)�#���[-&��Zӄ)Y�$KԌL����7��@�k���u����\د��v7Ƈ�uۍ �PdM�c�T��L������GGz��w�@/~1���I���Q�'&q���l�֩�Xu�,��EHrt|�u���_���}����EN�H�N��Ыo�a��֔�t�U)nV�zd�KĒ��(��ˡ���9�"kX�b<�r[������ْ͑5���A��M���q�b�c��C��#�� �&��?�	c|j����T���ɺT��Iy �ߝ���#J���B�%��Up�܈O����w� ���O�<MY���*v0��3Ԝ³����Ͽ��!>Y�M���f���y��"�m��[�N�1��)����DK*vx�9���-Ȥ'Q�p�E�����B�Z�aS�jK��h�0&��˽mo�-��(�n���mL�^K5��{�:^���3�c�g&;�*Z���4��M�M����X�����d	�@���I�un�!yvˮ{U9�E�x�As2�0#w������ˢ�T\^��ܺ�Ru�@��À��g�����{a��k�[3鳍���t�qu��C�E��wKy�ySu`�1hf�i襘�S�	Z�&�9}g��L��.���&�
�JP�Z�i��A�{ʎ:V^����t���MdX��$6�CZ$�<���5vjqK`3��ؙ	c�(=�š�&���q�j��Wfh��&���[e3gZ3(��m�S���it�f�fu�w�+a=U����Ӗ$�)��5�Ug�4�8VrNjZ����1�t��u�`���j�����v:'�����
�a�_C�UUhEhF�V���P���I��tc���ܺ.�o;�}����CVM q��.H�%��f^y����#T`c6����r��F��Ə�v)|�{xZ˴�i��k����=�dl�Գ�/�gdiR�7{��ʒ��1�����f��G�霪��g9�}�����0wC����Q��PT�i񪯄^��p�7-�D��Sw7^N5�����-��I�e�3��*��JA��5.��p.��.���I�]��a7K�H�$�m%%7�;DU�U�@U�(�����W���K�=��a��A�<|W�33�B��tWMV��P]\��Oc�^wںV�0�Y�Iq�`w�8┡("���\z�ܪ��c��Pc</Uu�8��Y��j.�j�L!��z_�}s�2�e���e�KKz�t�XL�{!��H'�dߤ��7o�d]��e��^�Y��ѥĀw>�ۢ�qj	��(�ߐ�PJ�b�~��,��D�� ���<��ΡO.@U����?��n���ZO���0�R���+�V��3��1;�Lz�����EG˼/+� p�x|` 1t��m�P�LN_ �+a)�q����w�gj�{*@�pO�[}o�eF��%���mN�m��n��2�&�.�<Y���G�:�.l���D���^A��jcU
KGE�)\F^Fj:��<���Q�ڵ���R��#��}�a,�0�qh=��}�c��;��B���>�W��|��n�Z'��v�R ��|���< ��G֦*}I�'%u��t�$� ���xA�&��K�N�I�0��j�������x�^�ǔN�\ϻ�(�
����s�\?����Yu����a�%رĊ� �`�X]x�gUl��P����W e�	�OƄţC6��ȣjڅn[����_����b}l0��z�Lk�jwS���I*��|nX�[O*�p��@�p&]AM/�ȧKD�9p���U2\85��!�w��}�׈���;í��a�rΤ�׿>��L�7 'ǻ���CEK:.S���W�@�r�����Z�	�7͞.�|�	��oj���*����2�1ˍ|_����u�P	�5-�ڦk+{��B�w2�2G�-�N�H�/4���϶LH�=ɮ��t�~�Լ�§�*��z�G�'�v����oc��Y��6��J�	2/G�,ȇ���^[Υ�]���:�*'U�L��^��⹄�w�3��JP��%�|}%����W<�V�� �B�^�m�Y��Pz2Z����j��<Z�K1Zۃ(�{4ڽLB��{����p
ax�@C�k��"CL�L� �D���")F#�.(��B�P�]��%�[W�֏h!׳_�J���?�Q��&���6��A�a��|���$cu��%��'�GI�a�P�!t����Q�0F*s'��#�ɕ�Ӹۺu����vb�b��p �*�"yb�ڈ�/���XP�H�aj�~��0 WD扒�#���;��4�R`:�9HPm��ԁ���)�jZ?�Tc�����p�'y���Rl�㐡��\G&�cۗֆ� K'�
�L�I#d��i��A�� X)L��,:�9�6.��uQ������p�t�ۊ��8����ͩ@#�J[Ys� ��GR�$�Fq#S�'Egg�z��Eh�b��0�[̰K��G�i�/>A�0j2!��@�l�]�'=�N%�S���$S>,��SC�)��.3�5W��-���^���ڰ�����!���t���#��io1��ia[���Dt�w�c.Ё�4�9f�ٰ��GCy�ȹs4�g�W/�p�	F-ʱ�IF���6�v�5�2!KG�_ZQR�zƁ�I�3�f��]�F�ђ��}>��lδ4ٺ��}�q��oW�
�ہ�Y9��\�f4��|����}�֪�r��;�/��FR���؄�%X{��g�����	4!E��ɒ]U7�zP�,��x�@q�#�sl�S�w-�"L�����h��!��ڐ|K����������]RL)��4��zq��@c���C�����#^"��:L�*�6���u.  �3�^��ቿ`��n�S�Gtz+�Q2r�r���X�{�4|��t��� ��gÛ�qr��EMj)���b�s{�;?�l�A*�
x��&O�����(I�����q܍�n>��bHMh�ңBިV.�[��
#P;�y�5]�xo�7�������>�c�ڤjZ��@�k���p�]6��4 -��ҽ'灉�v&f#���(��!�>����TBdO�_w��S�-;h2D?��vrb�n�"+2M��Y�[,��=�\_��S�?`O��K(E��̖����mYn�\��=?��X��b7�X6�i�n ���,�k�J���&�[��6$�MY�_�8�8�S�` ��P�.��g�|>���Lq���=;�{�H�(�)��d�L�ҨRAH-�_*L86p��������cU�KG�:�]���
�"Ū�}�I�=�I+�B�M~�*��{�%�j���-	P:^wI(�|�DCrc�:�������z�z��1������N���T-\a�>'��'ˁH�:�ωH;a3��8$_�Okl<y5!n]�i�`هe�\rp����A�"�~��. �;���F�0'�N2��\���<�U!1ϽE_B���Ɂ��T�X� Q|�1�L:�����6j�D?��Lѫ��*H��x���L��j6D���{ϾBK��c)eej�g{�lr����r����á��x �ˋ�zWYL
�����JF�t|���p�c�Tr��n�৊�)"�"�����������`brT1��f��j�%����9@��m\��O<NauZ��x�(��Qy���]��J3�R�d�bJ��S;��X����%n6N��P����)��x_8Υ�����U�\ց��C��0u������-�+����8� ��.5�]Ļ�'͖��}<��8�_	�穈�#:�\��f�w�b���?{�k����j*��aL�#�T-�-h���W�����������ȒCq]O?����^��!���4�nO�3 ��Ja���v��G�)/.�rtO���ġ�2�{���9G?�"��0l��h���H�HV3�7���D�,PV�ir5;{��x����ܦ���b�1ђ�K�1˟�#^G�m�;���Af㍧gY&'�H"<���Ķ�1"��:�L*ɘ�4GcT��̄��@��jQ�)�[F�@�U�?HΒ��,I�[�Yr '-;O&\~P/�Ѿ&��^*cNN��]�2~q��X��/�w�毄��W�MY�����a�F�����\��+���T����u�YM˯�"�I��Jf�_{e�q�.��fC���t%�+{�8��Ɨ�m�Ֆ��� Y�羽���3cɊ�x����q	�zk[��������5��6�P����t5�u�V��T2h�J{��[cԩ�����7*]{���EG�ش�¹�z�y�=���`�b)��(�$�j�����@Xi��O�uK7�ɲ{��^��U����ׯ��E�D<��y���i^�K�ن��S���נ����B*Tۯ��[R��oBn���a=b���c�v��/�u�I�s�ũ:�
�8�Ҳ;�-]Ȧ�CA�!e ���K���$d�Q���&|��<��>���0f`��tuР���A"b�NX�����5.��x���
�/�ʳ�8���o�?uͳ����Ѐ.�K���),Q���$4e�o�,��^*M�<�؝���I���M�븡����@����~bJ���ѓ�p��	�M0j.��I4���a���T�rM`��46i�C|�%چ��S�`gx��3�f��ı�����"ۉ;��Ĉ LF�g�K�S�v�L�n!�ɓDfET�V>Ն���%�#����2�����d����r���1i�b#�[#���_�Τ`IX$Ӱ���#����l�K��Ѿ&��}�\��R쀻z�����LS6�[�[tʷz����ݮ-��'�\���&�A�T�2����qK�-*K�k@N��E�nP�a��<LP�˂b��Y� p(ڌ�lV#�(w63�/����g���0��`##3�+U�E㣇>0B�����Z���kj�[T�ͳ�bR���M�)+�"�c��]��]���9�P�F�����b(�n��k��� P�do�P����Q�l���w~ؑ!�ŝ�����^�F.�s��~�X���F/��� e� "I��h�׎�i1���i���2�� �DW�<��2{1�����&�}�c�U�3
�Ǻo8*u� m��6��C����U�Zd6��P�«:#h�DY�:�02�L3Pn�����J��$5Jq�Ǹ��qbϦ;�q��"�?<�rk�K5�J�'L�t��S�&,�ǌbiA�Wx��4��d:1�_�|@�-����E�yNT�~���!�D���>U��a6!��
����m�Xr�)?�X��J�-(b��5�a�A�MB�����
:�^������?���)��eQ�c��i���"+��%��
Kr���-3�=�WF��y_3HCN��.��iZ��UC`�:��0��~��|��2���SXB��Ca�y)� �Y����e���'	�ذ9���SJ1H���r_J�Ȇk�����i�emK7��yb �M6Y�~0������/��*�)ں��pq��L��3���Z��y
by��rt:���8�W+(��u���T�l�n]<"��7�j�'Qw���L'_Ύ*c"�2&$kcMs��E�D�k!�Z,���sث�g�:r\G�d�}�
^a{���T<����b@Q��kX{��I*��d\:��.>5��O��/��9 ��`PV�j��} s.�\�l_�����)u��e@��DJC@���Jl��_�#���Z^Rc�(�Z���Ϥ����*�K_pi-�As���1p͚����h���]FثN��>�S�
O{t�yxV��R��eq�C�	X[���F�-y�V&�`���n��O1��0��zE%�dY>� =3͹S-l��w�*�jeI6_�%�i�%�^��/+�O��IDkx��&
VT�-�]�sI���<�1�<e�4���"�����y��A����)�wk������5l���ߓ���c��;���F�]7C�p����������T��q��".9O�ĺ��n���Ps�+*�V%��/��Y>YĬ�T��ZcO�)/���i��6�,�V7
?2�"����7��V&��U_sd�y@]�
��Bu���Ҙ�K�7����<�GCb�Z3y���@��w��c7�mJ�Y�s�z��[m�|�����Rtν��"��\x�UQq�Y� F��z�����䙭���φ�(�c���'*��ƔV�xW'W}��P�"���,�j��h��$?bB��� 
��i��k�]���A��s�\2�5��[v�'���"��X���owtIe�/~��ʙi)pl5�0���ll�Y�g��܍�u ��-�ԣ8Lmh[��m���	�L|�62����q�Z�1.��ar��
��.�����l��`:�w�;	aa7�FM��A�{?Zg^��wyrFK�e3�u^[��P��<$)Xe�|w��9�,R[T�^9Q9J���4�u��m��hf�	+d�U�d�ԧ����2 �S�������ٰ��H��*��_���Jȟ�N}�Bn>=�T�B(]`_R�Ѭ1�&��ey	E��Z��Q��qp[����	���%O*��Ռ7^P��5���߄y��yl�t$vM��d�s!��!/ข����-���?-}?۝`��#���}� |"`�c��~�n5�M����RΞ����o��-K���
��_6� U�=E[[���c��|�h�Mx����W��ZT��Y����B�i���4~Zl���'Ä5���.�7��ؤ�#��J^���s��6U�#*#���gg/�u�P��eb��u$0
�=[t���m������^၀�����뒒��c4�\��S@{��In*c}Q�,��Is(_rb7��0���ڶ�Myd��"O��d�5g��my-���Q̡�c�1�< ��>��և���]0"U�9�D!*O0����[/\!:)��"�	1����m�GZ7�YU{(���AŮ�s�dt�" U(���R����~x�q��̢��w~m���x���		��m¥�
�->;A@��e�]���ű�zz����Hf���tM����ĥ�ˈ�HF��g�:`A�
cl��A-���9�1���oP�,�c�QP+�):vL�&D�O�%z�o�ق|����}|��js��|���#���g�\e���ט�fG��^D=���<���m���
���fy�Q[Z&}�Ph�^��)��8��)����� �Bg�^�w������Koq����=��x��@���<��,�E�1?L��z����P��]���[r��λ(��v;�xM���%n:���H���9�,�L����(�>VI��zƻD��7}ߟA�t������e��py�\�E�I�M��'�LV��L���S�3j[vj�A��t��BD
{��;�Z7��6%��KX�}�f43���p���?��t+��d��:o�ͫ\���W$m26��L��o�*L����	�WF�J`��	V�@��9�Miw��V >����	�����<Y��F q+��:�ֱ� �xr��Y��K��`�;k�#3��L�e�htc�E�c��y���h�\,�]��f���93i�ZHAi�5^_D��O�V���̭a���OY\���t�f}�{o��lb�e	(�Z�"<��'gB,�$�Kg��҄<y�ρO�z��$����=��8����~��A3z�*����R��8ksn~n�] /*��>��p�/3��	N�F���%@ք�� �.��&cb�:3s��+*W��H�G�`G�:��N����R����f_x6>w���ǅʃգA���͛ �	y�pr#(-Y��ۈK׷mkI@D*N)�yꯖ�٘�I���/j��O���T��=#�.?�2����"�"Fv'~n�x���3 �kzK�Pl�H��(�ޘ��,q樺"2)	8�P��pmr۾�(v�N���sȧ�A>�ԥP�-�e/��BY��~k���V�F5!H(�!���P\J~�n��~�� ,��uw�%�N�|���:���zoV ��'��z�����T�*r"+�<���ފ�RW7G��)e��4����I�JJ�������AP�$�z���;�ԬW��r�
���:����x���_�I���~�������9����k\����\\R'�y��?��������ٝ� ��9�*1��2���ĳ�F���_��������Ϥ>�Z��8�sZ�P�6庶���wl=��C�"�Y&�$��b�{{�>u}Z���Jv�qo������b���:Q�hK�k�f�D�}��p� ���%�k�0���}���+�*A�zӁ�؊���,�[�0A�o�K����ce��5?��)��5�ƾE�:;h5����b�9�pB�� /�qIt��ҋ���`;���VH�)M���ض�!�4q�-'6~�ʬِ6���KԲ����e�����;�.�J$��O���`�qO�#�S���b��r�<i�ISQon]�*5�%�N����`�.��׾/��
�G	l����Yrr�4���kA�Z�j�f5.(D�a(̉Rw�Ux�3������w2�-n��> �.�P�͊��;2��b4ĝ��Tϫ�N@?~��A N��d���'��N���kCU���i����z�'ژ��~؇�d�a��`�6Oy��7�$P�R�Au������d�|Ʌ�hq�!?/ĉ,F�t�%������@	e�,�s��o�lӭ,��Vg��I
BDo-��Ue��`h``ȊS'�k����ْ�D�o��}*y��=�=���!��n�f����{pk�ӿ�|�p����e���AB/Cq|������:�樆�E�bH����+$N����8�`l�6��O�O^{���q�����]xL�(C1�>������3��+�Jɐ��9)0^+���Ͻ@H����`4E-݁!��hB�}�-b���b����c��mz�%�Z1i��um�c�w�Gh��g�X�i�3��G�A�.����x�ì���-��B�逅�@��{Ĺpbs�z�8��-	#r���#ߚ=�sMh����f��k��a ² ��]J^�Q���O�4Ꝯ��;I�'�����9ŕ��ݬ5�Է4+U'/a7���f�Ȱ��/�6D��ŉ�u��rO=�ݓӺ�����E��H���q���R�C���#w���4�g�<�'[�'A���Z4W%N�$hO~O<��q ��U������D����U���z����O˘��_�F���ud�A������O�o�:���9N�bH�἖ ���p*�͒B������x�]�i��p�W3�4�f#Y�ZA8ݰKAߕn�%U��_�;py��_N�=i�j�{N����I���+��إ	;���k�Hv��9!W�j�޻m�]����`E���%c5��=T]
��Jf(�$#8� ��Z5%�C�%&���5��QY��;D���3�;����Qg(�����<�mj�{1w���N��ð��d(�I�����M��#+��ȗ̖�.�3e3g��c�x�(wfYuX`y�`���}$�=�F��ԅ������Q���C���%�7˅?�r��2Kd���>��%��u�;:׼�ˋ���+��#ԥae�������Ű���^��)���E�����f�۸U7�Ah�o�mDM��㢴utt�EV���qթ�[����$.ҵ�z��$����sU�f��$�Ƚ��2����-���Xb:!ϳX,#�<�!�@��aW<����V�lH�Qz�HER��G{��\�!�ww)�d+3�M�%���Aˏ�kx5���7Q���/
$���B#�P�x�(	��2$��(^O���~G�Ҁ@\�1�����mk {/`�g�$��y6���7���d=l��8ɺ���a�O��DRC:�>�b�p�����k��y/ȼa���QG��,G*T�H.�/����v^�U��K���=ae� ��F{й,�?Z�Y���+�u��3/	�fꈠd�tw�[	mFi�s0��k�h�7�4	�P��R�8��wu��s�hte��看|e�߶^cQ��mvR��`_S��>��}aKru�d���>��0��#�K�k�I�l Od�h,�&-)�~���6_���8���^��:bC&7��1xM� �o��~��ծ&�~+��ؿ ���Z��s�a�]����&�)T�2���H�0�������wI�-���ٮA�G��傚������9��/������븋Γvn�9���x��c�zIG�9�8Hkݯ71|�����3*�V�"���z`Y��J��%-o�X!�	����#��?�Iַ���Ss�����O�e���;�4Q2��AB$s8��S�N�}��]����	s��A�"W��%�����A�ʎ8�ި��\0�v�v���&��Ý}d�$��+�ԨB������{���E�A7�|VJ�E;��D�cE����t���vB�����&j��|�XXܸ�]��6��_v������ZƗg"��v��2
&�u�'��Zb����r�ώ���K��>��tw�Ȉ/�(�;�6e%��I!K*r���_��Cuy�k܁����@����půS�mpH9>�_-Z�>F�eΖ���X\���s�����٩����B�5E��C�y�
���&<x&�f��Uv��C�r[�ضDL���Y�}�J_r�y���ż㟔g��@����.a�shS��@)�#��l�b8�,_����<:t�U`�@�x���!� ���k��r%m?ky��*NE�(R18ӕw�u�A'�R��G����Q'�8��nMLÄ��t�t+�*��;�Bӥ��9������]�=9��6���o?R>��Bӥ�곣��0b4���>7���6�����)n/��w�~��)8z8�Ա�ʹ��r��pF�t�tt:@[����&-;*�6D�f�"I���U]�.3O���mE��Vu�󲫞���8�%@�����-j{���v����a�/a%��HN �:�t��߮���Q&��S��le!�=�"���6�;��f.�8\���2��  ����s�pЋk�i�}M�b�PHϩ�yK��f�n��6�=Xd{a���#v�up>(J�Hbk����������Jop�*�XX�Q.����;6=�ϣ���M�D�l��|��l�������䭈�/�"�"�U�ȓ K�i���8��@�T���7d����a��>���G����F�Q�(��`�w��1�MS��]��m��?���D�����O�MDJϒ�F�Ȝ»�t��U��[���L@�♎'oC	�xܡ�l�	�|����`��A zmM&7Y�LG�(��a~�����z ɤ���2�C�h���C<]��ɪs]��|�W�Bnޫ� g�;;���9�T݃�����|��vj�i?F]#�UH�K�9�u?��o](�i�W��o��k�ҧ�'@��������<՛[SYH�N�-�[�!s�=�#��{[b�>�/�7��([Qߜ��-*�m.��s<����k���m���g!�Ej�*��?��������� �X�ؙmD&)91��ެh��ϲ(�7���_C��Ί��B!F+��зF�X�gC:�GҰV�6�O;�#$�#g*����cc]�1`��p}&&�(9/HJ�{�`:�w���Pw��46 jO�4�o��-��~":��%����z�e���~ �^�c��.BRs[R�O�i\���=�IN�������w~�T������, #đ�2m��/V���+J�0	�(�&'ɼ�~49i}�"G��@B�O>;�D24lų�I$�9�u��y���I�^l�l�J���.9B���
P�6��æ������	��Zw[�{���!��Ü��J��>9,�ƇN��y�I���w��ƍ�Z���ȏ�'�q��]�'3�2{y>���Ud�-ΣOm�^�!zj�wE��-����gF���z��D������~�{e~��$��<��uq ac�O�X@>A��y�M�?��2����tk>-	�]��5*��4}��kV�EZ�܌���eD��9Y�վ�x�ǿ"��c�QAK�@��c-�����j."�`��@L�:"�u�L��\XnVc{12x���#h#y�C������ʑu'
AF���@@�Xl���ɡnR�hd� �� �5|䞇S�Z��IvX�<$!+�Q��h�������]W���1��9��e�^S��w��kWB�ɍz"bK�����9��*M�� "��ò�1��y��8>�_��$-��0g2VP<�ڶ��w�=WY+EK���T��$�˭��/E�b�����ܖzvB�cܜ�d~�v�J�d�q���b�{/;�^����(I���P �����i��Gs��vRv أ�����8b���F^��V1�	cCCKҶtm�����WkFὛ}������a��� =���Ƭ��%]3G>ܪA��و��VJ3�μ�Ԇ 	lq���Slb"��GP���S� d�;�����׫�K���0xѮ�婒�O�W=-�����%�2���nT�Zq7�-6w�{�{t!�����U�R�7�{#3�17ۗ�*�����G��& �X���ӟ1H ��=+�}��i�X�mB��͙���>��rFU��^F���TL/�/R�bU~g�T���/<(��?��L�ӈm>a8G�A������f���T/��^���c��_�<����V�.�	�L�=z�W�ag4�b��_ �s��8ʺ���c��3�MU��%���@�|$:YK�'�I�-�,4���±�h�{�5��y-Û~V��O`�I�����风����J;0���ެ�9i�;t�E$O��De"J �V/�(���ߥ\�G�
�(�O�H�׆���B�V�����&��{�z�
f�Y	�ѿ�SC�8cyI�PO�W �g���o�B'�'�oso$l4�L*�#/)��z�������a�),�j!|��gA�\�u���j�"J�����l��=��?.�5gP��\͗�ЧkY����J���5[1� ),�hQ).����P��}v��Acr~	H��I����R[-8��u0�c`v�����^������;�#%��s$yG�	�d7��3	��^i�zM@��q�C����e�2xW��0�8 1VK��͉u�dq,W�8��|-�����J���pX�AoW��hQ3����1�Lo��eYܙ�����ʄ.�� �U#y��������k��Ǧ����zl���

Wk칆��F�����������Z��y(F4�����2M���3�Y'mgIC�d8�m[��������^���e����%#�t9� s��4�Ld@���;zz�e�{4���h�R��LՉ?�A2���Q�_"��'�c;]�(}G���� A�*K�T�s�,�T|��'n?�ep?���?���x�r���F KC�qi' �d���Nb�c'��j�Vh^���:0d)�c��En�	�����8�[xR3���"y�ƌFxj/\��^R΃���s��zRɱ�ى���Q��%c���k���y�� ��iH0�/E^������8�S*D[&���+���|y���n*f;��</�n�]Q�G��Y��F�t}�[~���1�z�|��~��T��]*E��m��+���Y;�M�C���T��Ɉ.S�m:W$�����9���!�=Z��(�G嬱L���.��׆�@N�J���Lf"O����܋� z�9��$!R��~k��/��{�
�اz�<Ъk��b����T�v���w�\\�>7���oE=�]�Ŏv�����z�f�a���=4��5tJM�< �y�_[5�ǆ#��Z,��7<1����%��g#|x�%\{o,$,-�薺��\mS�z�ZGw1����R>ŉ����E6�">�m�e����Y%��9��p5Oҳ�%�K��l g8ʉ�ZOmC�mp�J�.ݴ����*��N�*��s$��!w�~�E��?����C�5k&�,�/�ld�pZc� �ǌ)��d�Vnr�HZ��O5 ���=x�,��,����L�B���{.�_�{1�i�	�ֲ@'
8���� <���;�n�6:p㜗�Ez���)��y���'��k���w�OZVA�s����`!�tx29ؒ�Z	7��Ug�`��Z'auKL�TQ�.�Z�E���y u����ƶ���*c�:wE��V~=�2-��UM��7��5����c�וd]��,w�Nf�z���^z�y�����y����۱Yz۫����Q��^�|�-X�f�$oA�h���SZX�M���[�%�9�p��ȯ �j�QԀ�xe*'ّh��Z�I���l8���u�#pMnѲ\o�I��@7>�����̩��ġ��� ������!?��F�|Es��F]c�S�{d���X7y`��� ���ߘ�@���M�t<[jŴ���{[*���;�b�Рp���C���*����
$f��X��;iv��)�������0M2@��g�`۸zybh��Ӊ����ʞؕ�a�w��W��M>�(�`Ip�Ey�>g����/ΜX�	7��z$��˔y����40�#h"Tb������<�"��\ރ���K{=�7���U��@������<�**
��g��!�7��q�fp�/p��+��l0EDf�u[c��ȁ+#�޷{ה%7jQ���N6	�O)���Τj�/>�i�h��tYx���\�b%��5Lu7��ѳl;�b.���Q�;�m�g8	ݟ׿�K'�R�[�0.�K-0����NO<1���{�R��'�#fH06��phV����M�*�O#�v�"�g��Ρ��7�L
)fX�e����F��(Q�8��O)���e��[�	�sw���<�jq��j�|�9�.�M�K5�������z���3��Z����fO�A��焫
Җ/k��6���`���F��tĤԁ�!_I&�g��D�q뙺�Z��?�9,w ��I=8X��ڕ��t�v�OYrU�\`U�� > 7�`�@7�N3W3E��7�Iy���>�D�]���ˉ�v۫��?`�$lޅ�1���&i+����؄�����"�a>�����t<�$��W��m�+���]?�I����6�����N�|z��-6!�O4.�n��p��d���p��QN����[���:tf���`���祡��5���whҩ�~)A�������e������i�'�{��-��X�F�0�O���p��{)2Vc���"˄ۀ|�Pl�Y�(���,쑸����� �?��R��Ci�Fd%��$����_�[��@�m'C�Qu��F��*�^EiX�P���Đ��dU��J��|7~���EQ�^M��h�t� �j'@�+�6�篊3�)�h���5��LW�Ƣ�I�J�ryJ�^w �㡰�0���
���Q�\��bx�l6�7р6D��Ck�o�;J������.t�ʑ��KJ�F�
v)�Z�3��`�Vpb���nIhO�	���\V�g�|����@פ$�}{�"�M-�+5�܎Yh��"c�����Nد�XX���O{�D@�o�FY3˟K�D@u������m�F���;�0����X|�5+#If~>��5����\,}��d���]�DD@�����w����3��6�����R����� Q�<KdO�����)]������'_C�wN`y8���?��2"&��f>�J/�̶����KThD������:f����S��( ?�ô֪ҋ�&�����F����a�X�o[�L�iXK����S}p3�`� �"�;�V'>jo�� :�]z*o�m _�/e����<x�j�Y�`�`����*I�pb��;��Nh�Q<1�;ХL��c�v�=M�)]��.D�	��cuH��>__��`g
���z�3������d�E�U[��#���yʊ�N�����"҄�_�q��&��Ӣ�X�c��v��V�u~�sv4�Dm�`��2�d���9�VV�G��l�����F?fTĽ��]���-A�|��[y?�-C��h?��F�[M� :wݒ��x>���7\���G�}m�b$B�!�ѤHZ(�&��ϼ�hCҝmu!G���3:|�]y�7��x���n�8�����)&�����%�
l$���ǜRy���] �
��l��9��S�%�K�6��7�~�;�`=����5�i��i���Հ�x�k���J��̓<U�Ryܰ�m�>N�׏��)��?qu��MS���=��)�:��/���X\Q�W�>���wo�ts006Z.02N��E����2OY����BJkv��R��,��;m�᤻�oJu:�0�}3���]:Ϻ���];uf�߁2���8�K-�4�)ZA����M@#_��*���Lu�����-��8�hC>b�/`".���z��RH|!Y�ua���s�����Z��1�6���>�X��}KI�[�`�5�TC���~	�ȸ�\u?»��F[���˂����5oIw@�fg�-O�T�SC������N�H��'9C�}`�9�)BJ ����9)�o�:'���~c](�Sz����ɕ~c8��
p,��l����^]�)�
'��$ H�F-K��A93�(�v�_�P�Z0��5�:�9Q�2���^�+�������<=4ɀ3n	n��_P|��������kƽj-�98Oyâ�^*oқ�*�&)��i�$W�@�]2�g����]�J�gS,ӛ����XC̩�ʪQM��E����]A�=���<��%���{9;Z��[�7�\F�\�Q�d��m|��8�0����% �q�*�4�1xPly3�3G��Ӻ���Q���"�*�-�j��>���>���
�����17�HXPjr�ٮ\2N3{tKhكh�et{�� ��LD�3v2I+��N���g�'�Ɇ�,�DN%�.��	�yl�n�ۈ�+x�ګS���.3^%!���ۋ��
��_�_@���%�w���raqYV�"2p��d�=p���\\K���RxDk��'Rw{>����X!{�'i�_E��͞+�2+0H(Q����*�l���_�U��%��!�����b1���:��P�C>ub�pP>8U�P��ʑ����=��ѩB�G����ZV$�8�3�I��W²#���1�n	�suq�j*~���%/�q�"��G�k.���Ս�+�N���9{��[KNo�Oc��2}�	N�M{TF����Z�+$�B~R���/��<���2gIf������2v�J�MN��SZFEp�8O��2dI��`�	��M+��H|p���4��8	��� ���=�O��6�� \nV��* ϒ�G�EESڮ_�^���gݪD �����cJ����c��92�`']�a~�è�*2��䄰]?e���g��n��2�]�N�D��M��O��í������l�G��� ��Zic��:���u��A}'+5n1�����ig�� _���������@p���w`���:c��3�/�A�47�g��C^D���J��v5��eء"���P�_�;զ��uR��Sy���@q���j�&���: �`)��x�mX;�BQ�o�s).?pq�WO��6�����OnY�ΕUNh�y-��1a@�L�����5 ��%>H��e͜f*v��㹣G�$��k	�,p��
-��;��-��[dԄ
I,��f�C"��a��j�}��iO�\0��y�}�͑dfE� �H��Q����WrG�{�'�(�ͩ�S��QI��.tZ�4V���2ry�qq0�PNC����y�.�l/x��!����}��J�/g�%Vg�C4����z-�)@�Ҁc��A��tO/�Q���Яy�O,�?RQC��қ��L������Ȱ����՞X���[We6�N���&�Z�34f�>�!6�x���j�!~��߫{���폯S̶>t�we�Ґ�^kM8����|��o@�WJ��Ȉ.�\�!�q��%W��]*nܥ�6�����U6;I	,��ѡ��`p&L�z,0]xK �V@�(i��� �1��3R�mY�E�*��(Ǚޘ�Ca�H̤�U�6��@ex"N�K�R �?�8$�L��iO���5�����!��t�{��� H��R���w�.���|�XL�}x]�XZ��/������\(ge�Q�e�-��P�J؞DN|���m��;������|�����0q�Ktq�����M���Ϸ�w�q ����ڤ��vB�^;ݷ}z��d)N��UG|�r�=�0�N���/X�R�诓]m*,{��ti	���;R=b_~xT��Հ���w���G����Ұ[MW�g�:�i����\�z�X�M�?���4Hv�������\��Z��ľ�R ��_j���؅�%~���t�.��	;�L�3M�Z��n��z:smAyA��M}�_��#��Rb�˛y0�Υ�Ē�!mo(���^ۖ�`�[X��џ��{8�E��~�w5l"����Y���@�C������� � 7h�h�t��4&c��a��fQ�I�r�b��%5U����V좺�����\���qM���$�8aT�lv9�*!Ϊ�:��}c#���$�sa�3�3�+�9�+imo��|F�[��p��eyE���e;�6�UV��Ua5v�F6��;�_��e��7��T�F�cNL�����|����Tv|C��)o������,����P��s�I4e?f�Nb,r�B
��t��nM@ӹֵ�t���&S��h�q!���3����d{���e�hT���l�ޑ�	����n�m쬭�D�T�����z��JwK�����ȼ�U�$-�A�i���	�`Tѭ���l����#�aaT|��Rm=���Π�Vb$;�f �c�tD�N�"�G��I8I����җF{ul��>��Y��*��^8�!{�\���U�ů\�-d滊ba���h�Q8�)v\��BF��7O�H��&��HzX�A �_7��/7���D���Z�������C�b�������އع��q�,[[A���S���T'��X뫲�&�!4���BL^����`���Q����_���`��~H@Av=�>C�KX�*wڞ'������i�sز�ɸ$�7�n��(6%�$�3ݰ6�:�B'� hW����	)=��[�n(�f�.��t"��#�HT|�5A��2#�Gz��Y@�;�N�E�sQv;`p(��K ���耣��D�o��k�r�p��� M0����k�r))�ܯ�<o�R��~!����ۮ~�*�j)�r�H�������@=�v�\��ҵP
�୸>��K�vX��i�}���&`�b�U��w�h�##
-T:c��
�{��%�J-�y������B���\T�Tݿi����"�{�rc��2M�|� �"��.�'��4��=)�"�[S�y˦^�lp5|�yd��x�͵n�*�mU�C�=��:�9M��*����H�X�4����h�܄Z�oC�Pv��@�1U*<ޗϼ;v��P��$�i5� v7��o����2�s�^�b�[��D/FJ')�{��2|���#?-�u�;�`N8ѐG���re���0��},�+@ 49��á��@��A���_�7w`����W���v ���L���֤�i�"�o;���2nc�ݦ�)�;ӚM^,z>�`v�/v ��\w��z�Mz�A��Y�O:���q'If���ɬ�ߙ�����C?p����g�,Z2·%$[&��Uf���r�b煣<e+�����̤d�j>�c#�(j5]7�����)}���D��ґX�U�Ѡ`�XN��f��H��a�6V�oȞ�Qtk��V��z0��#k���R��K2NO���h�����+��2���+�_�E�j��4md`(�rX�x��t׌3|Sr� g��Q-�AH�mSZ�x�=�[��T��C&yipy�wy�����O
Z��p�/󔖆���Ҿ�D�@���Q���,�j�{r���C#���N�b���R��$�'6>�� )Z6���b4�ܞ��e>�3��7Tog�fI1�lK���ڇ;/�Y30�pf�n�N\�B�pq�Nq��k�#�7�����[1�a&�Q�!���׹->)�6�O(��-��د�A��q���:�b�4���_۲��k��β�"���TE`���rIq���CRg#X�������F��͢�k�d6dX\W�����)D2_�%<��F���N��I�J�bͪD�Zv�u59;ܗ�6ΥA�?&\� g���7��kg�bPqj{�p~�#v�Գ�a�� a�0 ��r��\c`XX�F	�*�U/��8XQ ��e�g����OZڶ9iC������(���ޣOS����43�����F�H��}RW#����׽�;=~��$p�����d���
�� ��K
_�zi��kg1��g7�M���-2@��Q:hU_��0Ϊ�v���XpD���A;v^���[s6 �>��>�g4�6�Ё�D�+Sz#me(7"1�?T���ҳAȭY$������nu��y-Mh��3����3XPQZKֳN����%+3q��m	�js�wL�J���>N�̔\��v"�񐇱C�~)V!}�����qv�y�%��	5���~n��o���ACo�7�@{C�`��'�S�Mb,%�iW9��l���?qr��Y�lQ���٢����s���v�J���Sw	�[k�UП��I}�:�t%�e|al}o�Ef/�X��<�_1S�D,5�������1����K:,h�����4p~��V}��R��oOw`{��y�W��>2C��Y�iGa�1i�Y.>���?�3;���Ǣ�*�ϴ�dt����������\�̴蛮�����S�=�h��$4M3�\����3��d�:VZ;6�o�wދ���hS:���E�_˃LR/c�E	��@�L^���Р�	�`���;]z�x�f�X��9������Y�`�3�KbJX��y�1�������jJ���N*��_Ks���d��S���.&��0XͧրΕ��ʹ8��>D�<�
�.�ESi?�����]Ø�Х��V�"�������aF��쀌t$�#�xx}�QE�n���io�gI2n���Vsb{��d�*�f�q�O�W�CB����P2d��U��k�ݔ^>>Sti������V����X�����u��u�Dx�C~V���U(qQ��=)�&�V �Tb���#"?���¹
�g�-�l8�����lA/9.p,6`����P���p�-	I���� tY�դ%#kЁQ�s����X��L5�:'���猬?�>DV��/@� m�2b	�IH����FR�\wYJ���䥫�d,գ����1&�K����6�=U��Yq�7M��%�!�X:0l''8%^sZ��숵�H���,@��5<e���7^��4��wZR�EK�*�qH,v&�xV��p �"C�ls����p|�����;�w��'r㯛=B�G!��Fw��'����9�X\.�]�Yܱ�N���S�X�:�����I�!��>1�¶"~�e����#�=�?r��ZI�ŏ�6��dԅ�����/�k���Z�*���F'�� ���19I�/�U��ZM�w`Ν�!�}H�+s�>V��DoZ��)�uX=z�}�g|�	�JI2u�kY�kwcz��v�'��[qDON��DgU.��Ǘ�Ւ�3�.G��N��󎬌���Y8OK��R��p���N��#�{�%�g�Ϻ��#�
��i��ŵ�$���rp�=����馶�ϩ���}��\��/��B��Q`��k�b��3�i��.�j�I�G?Cn�W���;Fˡ�8!5 I���wk��C�)w���̏+Ʒ���/ʫ8�E��$���Y-�����s:�����$�_3z+��e���ˈ�8Jb�y|���?�N��eE!������.*c9���h����o��P��~�J`=λ�h3�`�������hƳ�@3�&x�<f��A�[1g�ګaY9d����� O7�?tt��Yi0Z�V12�Fy.�Ng ]��@�5`��:�cKS�����pc[���i�j޽[ʻ o^��	��	��0�܃u1�P��gR���@57�YT�R�F<k��"e*�ݝ��Q���Cտ]�h�
��ٙj9��ਵ~H��u��� �j��뜒β�X�q�AlK���(,�w�L/ �	a����际Z�5��+���,S61��;5����{O�.G3aZ�~c���p���r>,�1��L��|�ZG��OᄄF��,�����b�h�;,о��-���	�F�s��a��x��v�%,ruI��i�����9va�(����H�z)�4���5jճ����H�DR6p��H7ը��i5����C4jh����N�P��ŋv����ڎ��S�R�h�EǪxk�baϺ�${�K�/k�]��H7W�o���;��k,G�������R��N�U_��F�Sm�`�]��7��[v�T!7������L݃V�#b-�J��ɍF
�!�g8�~�.�!��|%3/�;�;ZK��c����\��i��l54~=��a�_����{m��|��H��5���9'B�WTQ/���3ş3"[V�4����B��GS=�/��miܬ;3����� ��p�S���.����Ht��@G
�X����m�����D>���a�=���1���a���}k��a�8�pf��-��sR���ƹ�-)JQ�߿/�St����W��9Õ��fi1y�3di�
��!uD�D���Kg��y8Յ�X������Ѣ�Y�d�.����K҇T�]��<��T�{���I��@��5WU8@���z��[��6�{��p �,|MK��������|�*�?m��N;�O�H4��a�5���̩�i����E�H^�E	�_#வ ;�O��9n}ٍ��0����%p�
���zh�k�m��mk�������;��S��6��#��]Oz]H�s@��zU�2k^�
�!�?��;�(ׂ\���I^$��WއAݾ�̶�]��������A�7�U��o�|�]QC�G���#3�(�j����ΰ�2��l�V���q�lC2�|`���F}�\���L���(y���yH:���k�6�7�IWAHxhU������ �1$�E��rDH�=*���Nݐ�x�<A@-t0�6؈�g�HIWO�sxg��Q,_Zƴ��T�J튉����:�fQ�8�8����k٘�P��]ͭF����J(���`�c@|B��[�vo���yRU`���>�S��l�0��
a��t5�+xf{��ױ$��\���]���̓�fCm`��]67��XZ��H���^{��fU?����O��㮩B�.��$z�<!��B��(M�܊�dO@�#1O� Tf�*��6����&�wg'���+���a���緲���}J�����t��1��fN��}�k0[�o皌`A���r�C�/��̯��Vw���K$� �ɶ&ow/?|����s%p�k�PS-9y�$��Y��v!ϷLc�34������k	*�_�Qx�!oȏ�6�:\�������Xy��WlM�����Ń͘�:{ �{L��O�k��5&ojd�F�[��ʋ^��h�ya*��H��F|aV��18�R���ܫ��XXeh
����}���l�iE%��DxSĺ�j�#�UM���\x����+��V�DSbև���+F���>6�0�9��i��Q�V[���و�6H?��;_]0 ZP�݁D��= f��.�,�{SҨ���C%Xcn���J��MB��xi*]�5�|0�ǔ"$fG�?ٮ�����a�|κ��Я�7���ob�leY�qϜ����V<A�,iX���<+������P���*�����-��2����x�Qp(Ξ�$}5���z=�_W69�T������ ����M��i��j�q�M� ~��i�{p\�yS6�������m��Z�1�!ɋ��lw�@I�����L ��9��tosp)����Hɔi$�v�#�h{�{�2�$���5CDǙܜ��q�]*�c�_��y�8�e#�[�ᾟ�����o|����7o01>?Q������@ӷ�p��לX6kf�]�>�^���,}�� a��g��4k��U�^��ܫ�̮	_c�h8l힧�ۭ��Mܸ��vRR�� Y���p��O����B�?�'\�?nwj�Йu��Ԕ���nO<�0��`�܉�c4������ �)��
+G��%��c�+�4ɸ6�0�|��b2�d���r�E�(&6qAC䀦$��:�6�wf֙����2yc����h�e2Bƒ����6���c$�b3{M���GV̳���?-3�𵇖ś�t�7T+�ƨ,�b[��l�O佧�x�����h͘�Z5����1n\���Α+YbWMU�\x^�&&t��l��(H`r��(E:�U9�ɿ�q�}<�Cf@�=X��9�����~Q�F���k����ރd^t``��QZuj�{߷%̢�iS�Ap�V�*��'KtV��B`����)���Ty~ޡ�ͩ�#J��Y˴恎"�^��f_��7��ZS������"�%疞�	f�w6�?����)�\���k�s�@❦�\�U��f�,���흋.� n��|nN"����sS�gEh���^SmOԁS9��l 5}�3���u�Ou��v�U��eW��?��RA��aJ������aU����r^=t�Z�B-��{�]S
�!LT�[U0tz��:_�\�@�VpR��+knp��k��m��Nk��U:%��A��D���r�u^H����/_NIH�$ũ�K�N�@�Y�,���vgIb�W�8�������+��mQF�r��@C�}$��e)�ٽ5I�)Ywѻ�zyc���%qS-
5z+�C"�����eU��]�6LY-4��)�鐭$I`�a�)��|$! ��������w����[�� �J�х��S��]��#�ٺ�����É��b��H�]�� �<��U��xEک��^�j�v�}����huF(yw�0Y����:�� ��5qȺ���}סF�^<�;�7Ow�*X3�ڈl6 O�>My�*ݫ ��7b!�m��{Q�@���9��0��=U��a�8p�	�F�+��T����(��M�q6e|�e�
3�AU���y�Nw3W��h�֬c�H���#�q��+�m>K�E7�k�4�x�L`h�'�k����:���څ�̕Y�Rʉ��j��I�%>c�a�I�4)���+aSCb���S0C1V�@�)�\�䊻��o��=b�}�4��˘_�[�����f����p~��A�B=s�=k3�V����� �3C��R�p���-���1?m�O�g�ܘA����$���' _E�Q
x��Oqk6�)<��m6��fv���B�<�_5l���-g
�2z��w�Ad��ыyO
�"~�a���2������� 2Ef'f@�$�%L".�|%�;�d i4ฮ�!�|�U�l��aѫ]�l6g�t���l.�/R�� [��}�:(��3���[@˾�3�^�dCe�H,�	��@.�{ն�n, �Wyߨ��PuuTN ^�'�������+A��L��/P�D��;_t�9?ô�!�WRHpu����S�$����.V� cFwX�p����d�D�CV�8���%Z4�Pe���ǟ�:
�{��#��W�h��RH��w9�e(	�(69\i�_�cq�`XR}N��~�r��Da�|A��1�M�g�.nՉ߆x *w~�!���g���������W�g��8.-p������|��e��V�/�B���ɢ��ր9���6�G�d&j����J��$T$��-H@�M��kD3��;�D7.}�e|����W�R��8���#51gR���Wڣ	�`2a��f1U��!����aQ<�:q����.3�=����@�y��N��c�Y�V.��L����Rh����}���h�S����ۄ3����uB;GJ��K}A�m�xf ��*6�IW M5�.�� Ư�"E�ho�;^,T27�Ѹ��q�v�����"�0W"\�)�aC���&�D�)*�VPS�2D�y0���-i1x!qm09�J�e�0\X�RB�ϯ0u<��^laK�\�;\Fn����b)ľ�O8!�h|� 29�:��zf����ϼJ�	,t�8���)-��{�ha˭�2)���tS�4e愺PCa-:�m�1^����<���X��P��+�tm a�
4|��}�X��cG|��]�Q	s8�/��7���u�k0��5��Qx���1���kl��gt�FC'���<�a�r7B�Ep�I1��-��1��a!��CrO_�V���ʶȜ9�o�+M�፼�h��*��gT�,ĞȘ5ң��R�Dw�<.�S��+��(N�_TEds�6c۱�,5e���ޥb-թ��z�Q��j
����&1��AB���;�m��P;Drj�L����'���%��&�Y�o���_�>���?Fn��O	l�K�` O��A�Y.^�Jp �O���iҁa9�~.��:�'���PnInbm�� 떮�N���;�C�2Ç������6?��O��=�� $3o�K�:f�R��������`�=�B�p�D~�$���r9aP��^�^2qu (��@�є��/G�)�uW��	�K�$�� ��".+|s��>�Ϫz�V2��`��0X2U�f��I\Dꪜ���	�$zP��Tp;f8H:���P�l��O uF��ɵw�xu~�ډ��0���<�l�q�{�˰07T�[ӚvC�C��L����y��י~��f��~2�3�����!>�S�Vŕ�u���`����񘉀UC=9M�?�2쌻�0vgr�|�2�6q|��h#�h\����mM�ZGU��B��_SA<s�7�]�C��sӽi]�w���ezV��_4E�I;͢�� \���c!����N41�Om他�ʨ\�K�!�y���j��a��������0��	nhV7:�%�y�w;X����ғw�P�M��W9ʍ�v�����5�;?V�G�moL�y�c����0�)|���%N-LQ� �Ğ�*G��g�l�*����h1~V�a��� ��pܡ/��v0�8+�ʹ���Vbg��78�N��u�)��S��9�;��[�iBP��0�ZK<M^F�ᕅ��L��ؾ���8E�u{L8�R��:���-F��}�ay7�>��n9���?��B�/�u~�M�㝬aYN��T,x�\�f5��E��H�����)B)�M}:�R�y?=e�T�S0��X��x�5ڝ�}�����W7�'z�|k��B�}{!��a	��2A��(NP�	I���?�e�(u����[����f�V���*��5�y���]����_��ic��vi@�YG)�Qg�*�H�V>�X��P�{���C������,�(� _���I�9���b�~��� _���IG��u�[��"M�{�
�  [y-
��zlJ���詾����H�%mC��O�ΎkԨ�r_}%K5�fG[��{ګ��K���ѹXh\��~��<�J�������Rjl�2�� h���75Nޮ"B�J��^�#�K3&r�͑J�r��z�Kx6&�о�/�����4Ăq��H	��.g �F�B�z�����Ýqґg��@��s�^�a��6}�#(�&��>�a�_�\j���w6��eC���nh0e�����0��[�20������͚�L�(Nn��Ò{oV����c�y��&�I䘕��w<�[���}O?�V*&� 5k�L����a��N�𸤂;t�`�_x��҅��o]�巋)����_���`	.�i���(�tçhS��G�E:v�`�(�y4��*�mE4��%w�͌�O�j:L��V��@,���;��b�h�6T(��=/���|�=��+��rtD>���:����j|0��+w���I�@�탛}~���m�)]K� �	�]b�,띥�N�������ն�aJ��!KoؙL3^S�r%����v�O���:_�t5^��-�V�֬��{���W��U�jfT����"g��H��X&��źf�ꏓ�&vm��?�����H���v@9#F؂j�6���v���'/5y��b�t���<hXUrrLDz�I�?�xW��>�vO���CNDopqg�$���{�W�A.������[#v�4���ARC����8eR�7���E��O�n������.խ��(.7����Y˘�Z]��u�0�m�4�*��u	zG�؂3���Y���+�Ju�U���9E�^��������{UL������6>Fj��}�>��^t�Y������U���)��J�|*�"Hn���~�a4k��~6ak������O�86�����O�Ǽ5n�+�3�6���7p�QP�3�����|s�>7�j�)^�� Y�<��l)��J�2���x x� �L��A��𝝻����0	��}?���TZgTesh���=1��G��]ihڱ����������&i(�St�&D�3���Sq���p��0D���ѪǤ �zm15/��k峟�D�������j� 7A���= (���l�{u!��	�l�Ʋ�o��>���y��r��2	@��h]��GeqE��V^�m�d�|�r�H�]� -���ۃU����o��'�N�4��j�Ps��텝V5�c�`Yf�
�Y�6�x4�L�Ձ..���bQ�������A��pB��S$��N��/�1{K��(4i�D���W�𒶘��
,����]�&��q�Ll�G�03�JS��v?��8�S�k�ķ�Jc=�_׏�T�-�|?���������3��N�Q��#O�?l6�]�~k"e��)u��v���G�%,��l_=��|8O�=:C�܅�F��4�dk��}k$����?��U�����yq�aIøW=A��dԼf���޵��~��e�D�n���[D0,�G���M�s��`��˚\��?4�!�`g/�YS1M�-�u� 7f�̹�A��­��8�ʟ����%M!M��ޣ�����,껱=ƴ�gw$���b�hk�	�]>cRE�{�;�l���#�ڳ?=���~E'9��(ʭ��yx�@�Q��Uƌ����5�Nt٣N:zר��s��,�;M�q�?��9�s�@	�M_�u�x?�
�H�Kz�!0���f+)-z�qbq��+v�G���j���!�|�|�iW=U*2�ø��ON2lc̑��h쉼`���҅���2gW��?�9'�m����G�
�C>�'�fp��A<Y�K��^c=���4���n�:��ݯ�̢a��U�L�Q���l�oح�Y�l�@�V�;p^�ex�\���1�����j'����_�M2;{ۑ�t	5�Gq:��.��:+��'�[�������3Li�;Mt/��Ks�Ý2H��rH��1�%�?#��!�Ӗ�&8� lʂ�h��R����g@s!��	s�@��7��>�gD}���R�<��uF<�ZkҔZ�Һ�~��6�#�����5U�1��a�uEw��-n5+��Xc�d7���T�ţy�3�QAc6Tڄ�C�6�Ti��?	Lu�m�E��rJ��e�l�9����V[��|�Z�eo�p���	6��؞6р�pa��!#x���ڶ�g�������:��D[�Jn?�f&:����󱍀��:N�0o��9B4 �{J:�"#���Q|{./v{���^��}��'ᤎﯖ�,ko�œ�7���[S>-9�,g�_���%}:f3Лi$��'~2�6F���Ҫ�2�����d�V�}n�or��8�����zQ/�b%�j��aᦚ�� 8�� TAFBk��>����T��cW��1b�7�K_W��h)7�)�YDǨ.p�2���A�b��2�4H�TMs1\�٪�� �a�q{1Ĺ�KW��;�9<���,Y*��D��{h�'�(�����q�������,�J�kt�э�W��8��c���]1C%��JBJ_L� a�@o��$ �1��xHfa_ez �&�@�: �t�`��P�Ù���BC7�A�lܣۗ!�C�&�"OQN�\&X箖>���/��$Q��n�|�Ҥ�r�!��ۚ�/0v��g��v+��:�Z\M��$��b���	M�Ё6[�a��������/re��%��M�Q�#�t&�]
��k�Ȗ���������A>����WTs|ݴ�t��b�����ʣ��u5�gX?�_4ڱ�nvSh�X���ʹ��hi1������A!ۂvD�X�97M�`���E�h$CR�����X����_�݂�U+��8�|������~ʯ�\ο����nbi$ Z���.�u#�*:��',�ej\�ѹ��"����ɪ:ʫ%0'I���p��s���k�$(�����d�Gh�*ݶ�6Ҡ��gr��������jѾ+�;����J���^:L`ޓ�R2���fH��np�OWB�S�>-մA�,�""R� ۲���?a�9�"%�f^�>B_G�/����&;��C���T�PHN}��xR'��m~e����G���!�X't(O�X�jN��\�]�~��3�c#6�u�`V�?��Ƴ�4.�W�"��x5�S�i'�Ѹ�g^~��	�mLE�҂H����l�G��9�C�5��T��	6/���6�1/h7c�[��"�pDڲm��s��<���0�]�W�6$GC��{���T�Ϊ�^�:/���	����g���"B�$�	����-�a�X�h^U�@�e6A��||QJe���4�<ls[{JNݱ�:��US^A�����2��d��{�?N���;�y�j[e���4_D^�}���oȾ#,։���(Ze "bi�˒�6 �Y��[33Ph$��򆠎��z	>U��e�Dj�agY��Tus�6P�Fa�o��C�V�YZ�6�2�/�u��;�'K@}�-G�Q��%g(�Ӧ�뜇Pg;�Tي=t��j�%`�������L��!�-���'M�{Z��SB{Ϲ���[�������=���Q��=z���[׳@[Z88��������0��'�q�{(GީX��`�d��#'�1*�����i5<-!�W�ԡ�����TWa��q�s���aZ�&��K������xn�}M|���?&��ˋ�\�W�HT�� ���\E�;������D����Pk��?2M�4��_�ϡb�L��P��(�8��):'������A��nW���Ac�`Wv�X�:w�����O��D�o�ll|�UR?�RR���j>��z
���� e��YT�E��:��2w3g~�8eؖ!!�����琘����lh��t���	��5��#gP	(�~g���x�)@��t�L͈5}��jj ��|��d��Vhq*�S��*�o���z/�T�6�VG��o��2J�k��ع�͜�;��g^'�0d�x.�� 0n+�+XA�S�x�Ud����ϣ�jÎ�6π��������:�|jrH��h��桱���DD<T7�=K��$}���	޽|p�DD��LZ�o� !ú�`E�X�0�w�j���E�]U���ӫ��Mppl�@_�H�9"��|�y�3��I��HEX�*�h�����)̘y����ðgEl����z�U��U�Fy��4��i�2m�hl�#C��j��r�^h�W�@/�L���9!c��2\4�D3�$�y=���p;�����FC����/{tO����`j�����]��V�RzBt�l��X#*P��Ҍ���Ե,R�ݿ@'M*ˢ��E�����ju��O��t5t��ai�����+��/rab�T*��6)F[���� ���g3��� i1��-�H��Qm�!vF
��K�W��9�'t�N�FZE�k�S�[r���O~���m�#ao�b�'�[���nȎ?t�Ŗ�`���uk��ծ c}�tnt��\�(�r��e���L��O)���9��XY/�s���I��C0Y���PC�@YF�_^o���1����I�t�\�6� � :*��խ�!�u�; [x�����5�k[�Â���G՚b�[��7����'��� �_�(U�Y�5�?6N<*:�/P�����H���2x�e�6
�T��$LiJb�	��ܹGm�U�:��C\Dַ��\�l2�k�:}d?�U��W.K۷�n�H孌�d�ř�,X7j�i�Z��X�tJ��A�Bz}HS_�j����L�H������[(zI`4�'�)"d8[U�5/����?��6�٩R�l�}�O�X�Qg���p���:A�,n�u�~1g�w�`���W4�m!8�� ��x�Cx7*��Q�t��Y'�̣���kb�	cf�!|G�	��.����/4?�:�M��b���o���U[CӻL�
l�w`2@��J�v�9�8/za�nDv�P�Kw �:-��V=N�P^ۢ�R�Ҫ���g����z�vpaå/m�I;D��g����
9�{b~�f!I9��NO�	`��c�zZIe=�s\)'�91�W=㢏�R	���T��5P��%w1Ȳ7�~�V�!�H��U�ȩ|�L��I����ɝ��e�)��C(��n��f�1��<�Hnc��[��L�3���#���1���^�/*/��{%��[nշ���7$Q̌@��HY��u4���ʽa�P�+k��NL1ۿY�ý²��9���ʙ��]*䘁�$���j��qB�*7=�De�ͮ��~|ot�F�#���}1�Y���U(�㾳H�1�B\���W�Ħe�Xs�<�R���� `����q�Mc�UO�N]�/J�c���m$;A���7�������:3��S�ݤ������XuI"��{[=Z�8=,�]��	/5�)��%�['���u�A����0
k������p,6�0Y�����w�P|�,�.��e䘎?,��O4"H �q�N*-&@�GT�ls�v�����Ӛ=��[� G&y9�?h���p��` J�-DY���d�+�)&�1�x�07g�L�+�P'!�l�ڎp`����V��$䃖@���_��Λ�x��/�>U�i:����})9�k+�/ٴ�ds��#(�
�7��P�!�~a��=�Y�	` ��1�-#��a�N�l@Z��\d�z[<��D$�^�~�w�d�D՚2�����b�P�!�Ct�������oS�lx��XY��Xcn���������#�cN�^#c_�~�V#�gY	[�s������g���Ҵ�q�X�;h����-�Re��^y 
R�p���y/�P��A���:ZR�w���!�ёOV���{�?1bi���b��#5P{-��	쟖���SD��u@@�05aF(%1 ����:��1xF؈�rܩQl��;Qm��8\���}_�޽8Xz��{%�0󖥳P5�t�H���v�Lz��x�l�ڥw�L�n2�~b�c��	���q��IF���kl���a|����]2��k��6� �[�cI1Ӓ(#L
���յ �nh�F�Ŵп�j��ږ>XT�_�7_~�����,�: �W�/�Y2���;*��u7���d�K�k�{������.X�����[8�L�O�s#@��90�o�.��Z,��T{�\�P�u�4�c(�о��J�2����?wM^2�cX|+�=�y����D��QZS�e�')QH��lqXN�G 7W�!�����@�������ӵ�5N��z�.��1�X#k���6]�#8-�EY�XC�>dB\9��/ɫ�GCv��6_g�hW�	-�)�V�;���V�a�ۛ쒯x�Am��ăm���Şf�R��@O��w���%����r�Dc�D�CZ��'R�	��/��O�8 (؟^Pci�}�q���Dy�V82�oy�4.���(�t�K��N@���͠�ǆ��F����O��n6x����f� ��8qa�CzSa-�Ou��u�
��U�c��E�Ͼ_)(J���e~A?p���R��LQ�aA@�/ �Zt�&��M������J;]0A*om�VcP�k*���Y,O��ۑ���ܴ�+0�����Eh�d��X^�[�*c�b#/�M�i1ɼ�Te��U�������LXD��NH}��)�<�݀f�ej��F��&#8��=����1�[���pt�� QA�(�r�H�����ؒ8�k)�G$R���b�1�)#/�@��
�M �A�y�2���,$^ɑ�}�!J�m���������s-|�;j��>��%��Z�}��,g{��nR>!�1���Fe�B��-���!��ʪ���2����5,�Л�d��+������(�T�O[���&%���}W��s#]�x�5����7׭|<�2��>������7�eBETu��Gԩ�A�;�FZ��[��؊���>����u��j�����a�A�m�IO�����)�L%��]��
jM�M��ok�r��{:�Sn��ҷ��*aX����_'-D��[��������{��_Ih@�K�<� |��xI�d�g���.�|�¿�4;L'�@Z�����H[D�_��^A�o���q����t#�`���CF�d��(�����+���_��h��N�� �9W�i�'�wX������R}��c-�����:!�����y�
G���W�(�Z��|��eE��o�w۷jp�u��rC�dB�^wM�aڄ]��@[�oR��yq@̎�������A��
K�L�֖���E<if@tӡTݣ�M��3
���Xt3����ץۏ��F3��-U�BT"L
���U3oWc�#k�,�����շ�4��.��°!�8��a_���m�OW31K�E%�D�B'�H�NN�+��{F=�45N]���{�dT�rq[����j.��lwl��|��&�N��C����p�2�|��Ϊ�wu��z��[Z�gJ%�<����g����GB�І�uX���K��"�d%������k�����O	.��;��o�u�Vz�`�x��h�M�!��4�E�<א,ir��*� �]��#Z����L�����9�~�����c�;���lad����z�`��r��
5s�,ψ[t��z*����}۞e	�+�e苤�F'C���?�D[ײpi����g\������=$RX'��UW�A ����Ĩ�|�:�$��3�/�j��kc9U��f���g����S�L�ӂe�:4�`�˂g10��k>����P��S�S�OZ����\�1���0/��	\�������}�0�ƾ�9$���ʪp7����mRlY����E��bG�M���Y�p���=&Y�b�7��gbC������$��܎}��\�F)5�]z���N8N
����OW�����B%�GƥR�q=�1�Q��j+��aE��$<`)������I���_�vSJw��4-80��q�����[S����~Fr�8֢�!�q5D��ZC�~W��^�.�Ӂ��p���4H�e�5V������Z�/j��q�^Bb$��\n�O�~Y������C�GN�E���3c�|j葄�,�	� �#�h���xj�0y�!�	�c�� :<�����d@3�O�Cר���$��uI���9���J�T���<�޹i~��=��q�+ת���&�x^����;q1�;=��Ⱙ&�����L�ffk��������}&�땆#���s�����Jŝ�aF�詞�v7�77��'�~?���#/.Ս�j�Je(��J4R�e���m؆� ��"�)VB�|��:Ɔ&:�""7��H:k�p�8��މ:ċ�4�8���u�z�[5���5�&Q���`�C��>-�4p���&�<+R�]:]��g�SP�����Z�aΚ��Rl��8��(��� j�n���_�Ax[1�s,�CUa[��W�߼�pǟ>0�9�`	���r���S�졷Q8AI0Nc�����]����V�� ::q�m9rhm�{X�S/���9��>M��d�sHU�1(gH�^�v��Y��|��<RkI���LVEæ�hW2/#��V>ǧ����KEu���\ӧD~��<�C��X�up���$��"�'N���L��_�2�h�
�{u�~�\��Ю_�ӷ���CUa�q��>`r�*r�05�&L�X~e������A4	�{�f�����׳#��e�9�Qϒ��m��>��ˈ��q�ŋ:�W�g��TQˊ���c��1��!�hQ<�aѷ�l�8�]E�m����,�]+���~A�G��v�FD+�QJ�~6q�D�!�];�a�����S�갪N.~�1���"!� ����?���s(��RY�Y�����߮n~	�{�8�����}�!��:���Q�ܑ{INHpVC$Z]�`������l��L���aK��q6:�P�T������CV��8�(U5��'��\�~�A�m�uϛ��Uju���dG�m�a3�OՂe��	ڻ�x��?�������>s�x��mA��y˘�j�
��]N&Jv�� ���4��d"ag
��{���!Q��$���P[�F��Mk��8�yAD -�];�H֧����4U'8�,��\��M]c��2���d�_>��$L]b;9������b牻Q�\P^��N�߸A8{�x'@���_9�a[�!�3��Iޕ�mD딇�/7���G�|�Ή�if.�D��=��2x"���q���u�qJw'�B�ǩ���T�34i�����͢?��`ؐ�3��e>���1lT�����l+�T-�䍬�a�g!q�L&�B�wf@/L`��J���c�����{����A�"�0_a�`�Bk���o.��Z�-�0�`Č��NZD��R��H�/��ϫ����Q�I�3�,v��� �r|z�ͦ�0�簹�Z���i_a�G�e8���k���hq ���ϖ(mp������(b�u��%��
����"DJ���F� ���<}Sz�h�~i*m����-N�~�W��v3+o�6�w�E���	5�I��[�g�	�� �����[����yY{�����@���-�u�Rd�3��g�����]�Ɖ������gM�S�w5��J�e �������ou�b#��Qo�O����!�a4���q!Z°�V���|庳o/6���0��j⺽(+�Ւ�|>G�zbm'��'tTUĈK�Nn���a��0���:�;A+
�� ���;C/���tՂ�q�Ci7ʨZHM?ƹ�� �����`Q.�3-��v Z{nJJ�ik���%ή�\�Z3�8��� ���x�e��L���8t�A��ә�ߛ��;.�����xVr��WMs�ȝ�0 �~􌭿��I���<�ĈQv�����}��<�r@x�����ʎX��L(A8\P�L�4~x����a���h��=3g��3���!�E����n���9��5��w/K��J��\�9��uk�?�4ȦdkW��>�L"\�j2Sk �� t�^@w	;�=����)�ˇ��Í��:�>j���չ��ԁ��	���1��yw�м*��17�O�Z�oLFڥ���&�����������������yqR�C}��+��Y=k{�������� `���q�L���8O*��f'�\ݵQݰ5��ߧ{*.m;�B\��E��I�[��7v�.��k��qe��Q���NW=�Iu��i&��e��lw)��/������dt�dJE�D�l�Ѹ�gn/��?p�Q5�0g9�-SHYZX�����.KJ���g���1�H��Q<�����/��)��œ.��&��R�B��vV\M�ֿ>d6X�?�4�-A����A'�䄀�L���p�����9�������tv9�ѐ,m��n��Nݯ ��%�9F$8�x)��EC�h�VX7V�<��.��r��
,N��&Zj�ͧ��2Ѿn�Ȝ��Jϓ]�lqF�iMw���� �#O�ؖ����b����Rx�+��,�Wٔ��^�c	��P�oE?d)��m���LO�G�$�.�'*�u�b�� G�m}5RSDp�"G�OB�R�4l�R�4X���\H�E	�33N��5b���� >i�N������&x߯�W
o�p}�Q[���y/]�����F>y[������"y���O%Lo�=�Ɩ-�т2+�x-��vU������_E*5��������i�F����X�ç�R���wߢ,<���K����W"U�@��X�:T��
�[�v�W����\=�T��Lݚ+���6@�ħ튭p��R8�����]u�z�DP3�(��w�_bpE'�hWOk'�w�>��?tT^�iO�܁�9�Ht��ߜAtCBM�Vb���#/����Sd�ddܬ Ɓ�RʈKe.$� �'}ր��VM�f�Cx���m��6�RY�E����o],첽�{�-���=���
b�\n\Q��B��60���Z��ɽ�H�37��ِ)U��\^�y9�q��Y�撦Ay�n)3���t-�`��B�0���ݞK���>%�$�l�&�LW�(��?s�o��*-m�H�eM<�]Z0�f<�B��A_b���q�冊�Md�⠶��_ū*���H�Mu�s�(w� =��TD�`츭g,�_1�X^=�˫°����rM��#'��6F�t��)j�9X+8ᙚ�敢��*��!r�uP��b��8.q�}�m|]������h��ғ��K���8�:��	{�h`.� �Mr���(P��-�ni��Q��Ü#�cCd���^HL�`��K��T^{�Ob4]��f�����R��.M��J)"�mQs�S�� HF<�֍L��k�Փ#�_bm{0(�H|H�!�D��L�A�k��;v�7����6�"��~�#�A�a��Et�� ���rp帙�(� Ql\�j[�Kh)��Z����a�9�F, r�w^��"�Ψ`�˅��o󮠯Y�2�U&:�4�jKj����XsOC�����mo���6%Tb�R����8�4��hL;�n5��f�:����3�[�YKk��z�������w!h%�Ó�?|��$��&������dt�;9+�"��S^13=%�޿�R赎1�������/���} ��$�q�c�HC����P���U��f�:`��a�zmA�d?{t�y:2+��qj����7��D��c-ǘ���x|� �N�ߚ~&�*��	�J]7�w�z0�7YP�� �Jx��$Oҟ��y�oO �>	�t4�sg��u�.�ڍ^(�[�p��թ��ԯ=����<����.�!�k������!��!}��y��Ԟ^?>��"t���!3���$�j�ߚȘr���JUb�W�b�v�|�s��|�탇<yT ��pطi[ǜ���웧�g��N �;��W~A#f�_��,*t�mh�lCh�5Dp�k��DޱF���(܄�2�R������B��A��w�]���k�.)����fb~A04�lOIߍGAE	���Pr�o�7��s���y�Η���s6�)1�z��@��(w=�JDq���~8J�DV�H�BŖ�2^�A���-DB���R�lJh2E"�E�Y*�������Y9�o弧F2���m�a�M�b̜Z��u�.����*���5U�c�/Էz���h�¾��k���<���c���"$�f@y>Z��r�.cI�2*���=��Y�u�>��m�]��'�,\�!^���?n��q!�Ϸ
[�$Ԩ��|U�@؈��,ڑ�C%d{Ĩ���A������]!�x�3��L\��򌝵C�^v�ρ�(��ZPS��\�%���Sd�?����j1H�p&�1�hb��yi�$���F 9�}�V�F!B|���t\p�MHd�X�jQ0��q����6�t%�d��/y��'����n�IfL��/Ƿ�m���6�w�?D�cHd����2��c��U���q;(��$c���oz�4�yɠ�$Z C��XCa;�J��������G�B#W��Z���N�sc�2�]!v�i��#1�,�E��1���^�d$ƁKv�˔F����`��J�v��L�! �C�:dHtseA�%��\6��I�r��R�l�B�_��y�����h�.��3��'Jf;:S��x��'k3h�-���g.�uT�����1�"$��N1�G���o���xO��K/��]5����MGY] �{��=�IUZW�h�J٬}�Eza1�ʥ63B�V��V���Υɗ�ѰNn�d,CE9ч�z�}��*�"Ve�
��Q13��$fô�=v}B �Fw���!e_��Z�$Fc3)��ԧ�:�� �y�k�{Q�b� �86O��3!B�`߀�x��|����d۞xg���R����b|=�@-*pF�����3$_�mp_�
��jb�n�~`hKe�6!�-~�8��P-�W����]{>���Aq��)	���	dF�ߓw��T�g�N5����Z�JEu� fF���Z����1?����ٯ0�P�B�%
X��{���h�Y�(J%�!�N����3$ܵ�w�$��r1^&�(<��$��J��k;gd6O�3�����,�F�'��_w�<j�\��U���w��E��,f��3�.t@%�����?^��G��㦻\��C!@�;.d֑3{'	��C�!G�	�kc��&m��V��9����D�FߒK�/�����J1�g��f�gq���` �u�+�"��>Y�1RRM�{�bl��+���K��k���׆��O�H.��c��!A��ב����W���Xm���I�!�����@zJ�_ö��{&U�' {��~�^2�Uȷ62�W'|H8BV>�H�Y;C ����xC��������	џ`��[�&S��q��2>�3�U_N~!�H�Ra�E�;B78[�H �%��t�|� ���RKF�C�p}Io�#����ޞ]o�t��k�#V>��3aeV�l�IJ%O�����%L<�D�Vs�(,���u|Tg����7�xr
�,5�����{Y�۾?P���C��	�D����&��kG����¤�BAxs��Ћ��h���}]��k(��{fy?,Q�;v|9F����W��m@�lY��oQCL���-�0��dۘYs��p1�1Ǩsj�E��d����+y,�w:�p9�)q0B��`�J�Ца��3�So����� ��$>v�y_���������ϓ����/EA�h�/���}+��p��#��Dk��1c���e1?(�yr�u[��=���\J��s���M'VSD�GgM����,�R���>E����u8}P���=�ɟ��tio��YN��@��h�e���^�ں�"KiOPs���R��U$�z�dBzJ��b�2)o[N6�Q�%^�`X.�CX_�3�Ĥ�c���G�jC,�4�J�	J����w�bZ����juu��CVl�'-�7q��*A�S;�>���Ot5/��7�[�"��{^��P�!�I6�[�>F4% `������>�i&}��`_�L��6��i��V�yR����=�ħ�oHȡ�ڒHu����l��T�6*�g5
r�&�iN�n�� �u7�ș�҇� Y������EB�n��%��w*o��������t����1:�0gj�Ԥ,��Y������gI�|�u
�T~��^ߴ�PwKʖL�C�}B�d�a`c��y<���HæLա�/Cˇ"&0�Y����ǲ����ؘI	^�������qf��z͈ǈ��0�F�y�̃���F�ǎ}���ǣ���s}��� ���q��{˰��K��6l��cH'倨�h.Ⱥ��$X��S�˨fW.���4�w̝e§�LT�6��_��O�9��D��w��P=��S�d���ɬ�>�}FL:l�x&\u"[�Cc�Tp�o�-���;��ɻ G�6�X4N��
V?�Y�u�����<W�ꔷJ�/�wY���y��I��9��'�bM2�P��JՒ���&#e���L�O�������ߦ�i#PVE��^=!d�q��B{@iR>ۤJ�����g��E�	㇣Ę��mH`2���	�I���_�~�X�&nr�Hq����ʌ�PS����{ꞑ��<.I�����٢*���-	��uͩ�]�R��y��pvg���+��+�(y[��nj�<׌���,$�82/���󦥙�ֱ���{͞����[﯋��׌B*�`�q��K��\�x��|�lwBl�3�D ���ݿ�2�=�B��R�s5E�q�^Yl��z�~��Q��)�u�ٰ=]�a ~���pb�U������)�_8�@y�4&��^�+'�\�h#
�A]��z��*W8���{���}���[����ck�C�$V����t;ya)�>Y�03#��N7cL@���%�q��0.ND���������e����3_iCF5� B�v�fD~�}u�K}(�T�Q�%)��s���`��rZ����Nڣ�@�����N�&���hΞ[��
[�n�*��RXt�;Ȳ[��Z�<�3�#4S�CY����c���<��;=KviْB(|�&3!|�yV���)�qvS��:�w?[�����0��K/����3Lymk>qw钵t���I5�Z�̂WW�ҀY\��� ��NB�P������5x��f��=��2\pO�A�s�Q��-���t~|��y�!�q��Q���v��Re�]��2t��+�3�f��7R�s�S��b
�Y4$.��9������޷2�e�8�O�!��?& 	���˻$�˱p���;��<�2���*"��.��]������X��'��F��.�� �ID-f��B�
+�Cs�{�w٧�0ա��37�V�6���x:��VSYգ�#�z~���O�_[�6�t[�8�$y��Yp�J��?������1���I�#�J=;KZD	�Pn>Ƨ�mX�ψlcGê�8`6n�!����8��%��Fێ�6��v;CK�-(A���(g��,aXJs�`g�L9��5ʞ����(�p6 =�pw�>ܶIē�22  ��g�&��ˆ>�n��_�eZ��,i#����飓4�[�
Q�qKqw���FA��k�lmF�4D��"��\� �>�	�L��;��������ι��fƠU��yx�cѪ^�s#? $<�&����I���[).u�B�~�C�����]W�
;��f����\��L��["1����ŗ�������@x3G���i�)}l|��K���w-8C�2�e��;X��;#��(���}�`Cg7�z�WTwh����!�Q �BJ]5j�I��J���������mP�0s������F�-M��FZ\0�������-�����y+C�!����pix/��-𨪣�P-�#x"�j'I����_���:����|=���^;�虆������jǃ�G��d��Iw��T�y��ٙ5&�<��3ӽU&���jR��'f�H��9LCo��w�����-:�LT�Ԍ5@�L��齪����ϝ÷�P��!0:�
��"�j�i��d$�[Z���� M��5���l�%�R_S��Э��c�BM�$��c:�hN�����ū¯�Cn_�Eن��:���
Y�Dysˡ��p����]�%�����8/��T;�"�� �c?�˶�_2pǑb̕�~߽� ���5�0�C�R'�Z��oФE�� ]S�K�i��G3�3�U�g�m����;�G�)k'�����]������z���^��L�<#%�uUQ���#.a�
�S��CW��X3&+�����$��S���#[%#�a�r�j� ��8Åڥ�����gn܁a	�B��8/�7��^#S�𴈬���F�TG��L��KR�A�"���>�W^Xކ[�I/�G������r�I���=��aOcܸ�w�2U3H��d���{�F�Z� Q������4���qb8����<�h9Xt�܏��=᱀qn�St�z����H���]�U3�T��zRQ��0��)��'�/&�-"�T�(-C�~���}od��(���k*�a+N���;H�n�1C�l��K���3���T�d�E��ǚv!A��`��6�j���q����`�3�B5L��}�J�A��嬸�<�r.a��	��&�X��H����ƈx�yˌ�tDް�Ԕ��P�z�99��w�fd���%�@�9��0��)��Iw�8{�kd�p˓��(A�d}�����^6���2����Ymr�G �0�R/\5�H��V�,a��^�b����/U����7���	��|�k�$#T����x6�	p�N��e��_2��N(^�2�����0�� �}c޿v��]���-}	�����*�K�[� �M�����fIw�f�2��c��s�N�#>)���S�h��|�6�I�|���.LG�-j'��g��z�?ֺ��a��7���@��> �b#B��%	�Y7'_�
�w��\е����{w�1;���'֟~�Tg��f64���_+��Ώ^�&�ꖚ�J����q3�����m�(�`�C��~��eݽG�9�'9��i�`F4��;�>V�d/S��Z)X��C_�15y�,�j�6����Cʶ�� \��O0U�Y��^p����1r6&�	��B`��h�:G5
)��,�[���"�P�U��n,��H�|���Iw�VY/sB�ezj�hwl���O�͸O�%W�5+
E!�(���R]-ߖ��h��=j�ւ���V �_�v�䈯|��Z�]�I�5���^)G\v�����"��g�����~#���W�]�*I��m�'z�Q�����䴥q2�1�AZ׶.$�p�]��Į��۪�x�|s�fs�i�{j���!�T�}׷�[3#"�Uj�	���fu��+'���*�f�T�Y���ধ��K��yu��?J!(M��V�-�4�\�h����+��#uW�UۆY/��:V�܎�"F��7(@K0	"s�)*Zg��ѳ��Š����>�ku�f����C�26g�19̜��Q
�i��R���\���X�z�s�{�RN�܉�jL�j���2�sa�N`_C;�	ȑ�<�a��O�jL%+c:�b�O���W����`�g�@|}����]B��J��f���Ib���t8͘|�N��P��^W�?{X�[0e�<���<A�cWc�	˃���4���f����D�5ߔ��x*M�ѿ/`}�0Ca\x�SS9�t>A� ��EL\�&'W���`�;QVq� �zQ�`�:�`=B�V�q|���p�9�pK��Y��^�����"�m�)i~�'0��q�m���.������\mǳ�ń��dK�M��0>;����:BtaJ䕟�}O|�,���{�.1�r_�cz��R'��ْ��ӭ�@�d��ET?7��n�9��
L�i��:�^�g��i�/�S�bY ����ݰ�!wR��,�7��+��K�B��R�k��=��9�3ŋ���*�V���$�s1��8	F�>a͝��I�:�����w��k�q?p��<�x�{�$��E�y�6�I�C�G��5�lf�j;�v&��𶌴k���FQ�{��!��Һ����9�aص�^��I��Ml�=(�x�	x��8�3�3�a��"��4��k��%�J*jtIq]�-êGp�
&����kCj�{��c"ׁN���i��c��Z��wǌ]I�P�#�����J�&�2�/�V9Q9�9��)̅�$5#���K��"�w*1�Vm̢ p�lΌ��=�C��_���y��5:a�F"w;�w]]lufB��m;��C�#U�߫U"���}��JO�����`���<P��w���>�� ��QR#�P@���F��`�}p�tu��	1��G�	Xs,=8 �-�5@��ʉ��BZ��1�]��[�Qi�>�m�e�SKAWuJoU���B͢��i�!�R�9;a�C��B���DKQXOC�3*$,�ơ�wm}U$�"�=18�X�)W�$(A�'�����WKq�C����<-����AZv�� )�ã��pT��mT��xg�PϺj���OTz"��ڝJ���}5m��l������d����)	ɽ��T���~D)���	1V�AJ���Ji};���y+�g�5�\.���$&��r%�pŖ;l�����n�K���6<�>���{)7|��H�ׯ�v�(9��̈́Iv�K@��˶�c�g��s`�s�%pSp�4}Q��.!�yB��Ȕ� + �Ism��ؒ�niZ��'���`�&Z��lߡ���(�u�@џ�w�BcO��L���x��t*�F�e�)~Ke*+j��;Og�Qf�M�0��"b�D�,e)��u�%�u��RR���D̄�^> ��Ͱ�fͬܨ�6���	�x��	Xg����{2�g�ݗ��3=zuo��8���wnAP���VP}(��l�v�;�������.u� ���8?�)���wfs1��q(�>�`�TCgS� .���fd��a�� �N���m�c�u�m2���|���w���oj�����G��E͋}p/��a$�^;W���P�B;c*�#���.�V���o��;y�������(�?�ñU���MWPQ��Gvし���1ɕ^��E��C�E����n��UWM�=��Rp��ea��,��)���E�- k���7�>��EXǞ\%�ژl��ZW��A��y�`��n}a��,���	���C]k��\!-ZC���3�V-)ȩ��?r��v�~q���f�QM�cA�M?y���������X#����A�xK)jtZ*>��o U.��$F-����4��a�cҲ��w��lUd�	�"��6��2k!R|>g=���c�������%����������B�P`˶s��1m闹��KNцc���n\��Q&���\Y�����\lY_���'9q($�L'���.N�g��~���Ǒ�nJ�/��չ�La5���D�;=�6��o�Q�_ 85��ǩ�rt6�X��}�+�2� ��'�O�x��'�@�C��J֊�ʦ�p{��CD�VV���������໵4|Z���&�袁ج��qhZ�8��Y�3�V���uz�v��� �IO�N��q�����m��Յ<ڛη�[7V�)��'c�+v.����q�k?��Vo��#�s6�����RX*:Y�iR�K�:r�a*gT4�W�GA����� �sB�7o���h%3~O��:�̯P2����iH�|��b���w�x8�z�Y���]w�Eu���zV+iLR��pU�a��l�A[X$`u��K������)X��Dթ�5p1��wt��6�{�u	��%#�!���R$��0%�PR�Z^&��U-��q�T|z���c���G}ȃ�y>ʘ��58��oS'$�C���~�6�vL���n�5��͠�����[�DC5�ۺ���8�t��M>����!0~L��S�|W�*��V������������)�g�z��8'$(Q�ǅC�3����ګ�	b��J�U|"Q�m��Y��a)�ƻ�9��cA-Ъ�(J��r"�@H��(jR.�
�j�4���%�#-���^�ۤ�PC�a���'�SWZ�? &�r�4�FU�眼1[�Y|[,%P��P}ێp �&Ⱦ9s��lx�o]�8�t�d�#�b�� ���("������p˰A�����ðI���Ԣ�d�FJ��U��}j��}��T�9�\��s��73��c��bL[x3M�yj��,��Ո�C����"$e_�)�p�Ϳ8�ԓ�2�C�&�����]Y���Ay'�w搒���֒/�����puv�\'QT Ԁ�_�З���Gu~���f-��-V"���.ào�8яU9���u�Q�X�)�׭&�J�-�~R��C�I�O���M]ì]�,�?,E|mݦ��C`t ��[�[m�v�f�{�!���v >p��.���(�K-�G��(MR�dtE��w��� �	��m���D.��sygS���[��#�wt��nV���Rx{��rv�&[$��U;Q��^mt ��!�V���j��Dk�<�=�λ���_��^�}�^o�?�n`.�Q�mMM��bT�Zxi�`��W��[B��TZ�����c�_z����S���輼ֳ�����^�g��T>>���L~���6/F�&�$r�D49ŭz��yn�\�����!TX�,X�1(��mg~-�Ń�7KM_��!aN�*<���S�b�ki�L��E���n���9mS��ק����������Σ���	���2AT|����qq)p0=�X���]e�s����>b�Ji����X��$����$�=Lv��l�,����9!E�����%���m@�mK��Б�6�f4F=��\X���̙�'�x�ћ��%Z��|���Pl��C:�22��;D0��rP��� ��S��ЩiC�C��W|"�$�Uz�,�l�Yε":��-H��I��z�����#���?�"U@.*?F�x��������@=�[rx3��6��{���?�n��V]�R�DW,�x0�'��_��A���ҍ���֒Qd|c�w~AH�y�TR��B�F��4�O�d�ω>���Vh3z�O��~w(�G�$�7�N��>G]��7��9^W�X���+^Z�m�oAr�B$����%��2���0ņ(�sZ��\-W'�����3� ��N?��g�)1%��2Б����)uZ�l�l�Ŋ?z��72Y0w*U��/��ma����l/��A{��v��CbQy�0.�Uy�!�$?'�~��s�&BMs8"����a'�"K�G���a��S���ƹ�z<�Q�ځ���m�;���,�[������A��_�V=���'G�z�F���ME7F�#�BY3j�G��1'0��vj��-C:i��n�� �0��FIp��{a�6t�*������n����3m�rhG��L��G�0��w�����2���j�2j0������O���T�ܽT/�%!}��v��~��y���it��˶��<����aJ�,-s�����l0+ƀ�^�u��r�AzV�b榆��ôzHS�_o��!uD�9�+1|�6�Zbɧf���ŵ�8�*��s,4��uA�΃��$Mc�bX7�@��op7)��.�@Ӈ��D;�*`�N���{ߜ�|:�]b�v������:� ����>������3�:Lڜ�\&(�}r��u��M-���y��C>���[�z���#3��M��"�V����B�T��ltV?W���q@Ue��������L%���/V�'p�]����=u�NK�yk�&<���D����'�e�/\��$s=@-����t��r9j�<˳���1)��"��� j9N�"f���y4D7~�Zqz�'b{S�$W ��P)XN!6�u��n�]ktQ]��� ���Ka�k�b�_�9M�f#.�D��yO�+"�t��j�|;���L�\�#���K�� [l�!̃@���K�Է�ĕN�G�s�tzkqK�!��m��C�t�X�������:�!�,J�j|�nJ0G�Nd�	U)����+��|�!���I���.�J����`��6�*hY�P�םq�de�NsK� ,�i�mB�ľ��+��Jպ[G�s�n�&���@���K������$n��C��i�v%�	�`~s���:�����2�ZO:�q���c�5���c��U����C?0"s�\����ҷ�[���;����BG�a�:�)yQk��^dvS)0c.rb�Ʃ��u?�$MU\x��dTBP��Q���_v�Ղ�L>J�@�\ϕ�����T>���@.��B��x9LK�!�Y>�?�ܿs�;�)�*���S�嚸ob�jC'\1��j��>�����`���	EmDCh��d����mh�n	��4��b����&�goq��g��!X��XW,O�,ɝO.���6��5�n���5������}k���8�%K=c"�p��B	��3���H��0�f�2��u=c��>��>�<bA4��j���GU.�pT�<`!]���&�d��݀o�SG�$l)�A�\C�ʸ�F�W���A���wc�yѿ�٦Q���0d9�6pU��$�����A���E
gաP�.���o��7k�ش���R	���kՙ�r��}Q�(׌H�����s˦�:ȷ@�|��@��.$���5`ǈ;R��첮~����UI��4���^'H�m�9�g-��y���!:�U&�]~Y%k}k�PKu���@�'a}jPHn����r��ݚe�����ի�G؛�^���1;�^s\�x���@��dw��i���web���F:ڈĄv'bUL��sM僤6��"��M��F^�eo=oW�En�2�YP�5{��@2T)��#Y�A-����^i�Gk���b����u3��3��&�i���;�"���(��(-�Ma3�g��c��=��v#�`��Xp�OT<uȻz��U���}����A�d?�:Y�$s�!��~r�F��_2��(�l��Mفt��Y�l�Nߧ$}�v�%-ʾ2˝G�2l�Ҿ�Пf�#e��r��ƋU0�Ҷ�q�&��%��;����e;��:(R��@��R�����~�p#ю�'���]z�{�j⢚5��r�3Y�7�ʇ��i���I���\�
�k���4=�(�gcd���i���ejÄ6��Q���z��v��]h��YE(Z�8aX�S(�g�%s%�]��}(v�-{�P��&������wOf��qݸyL�5~k���Z�:hH�P*��.���7 �?4�G"�O3eE��$�t�%frų��wiK77��.�x�^����ɴ{g���Sy ?A���$޶p$��0�8r,�l�]xj��ۯ3C����Xj�}�$1�Y�̆�ozZ�	T�������� N�̷� ��u<̅�Rb4~��������Z=@e}T^�7@d�=.�����9�^�OX	�̡L�O�ʙ�ٚ�3˗��,7V)���H5m�y�fW9��-T?��l�g��_��8�NH��:`H�����w�sD�֌vmH_	�Μ�d���5���Lϴ��;
����]�kᴠ�W&V����|��)�Kt���j���14�??�5d�$R�������޹��C�Wm��L����f�%a� �=���?p,���D��m�?�T�'#H.�� �S�AIJ�9��fTK��7�Sb�W��
�R���㧀
��'A�����G�$����(n�U�̭uwg3���f?��Z��� Qɐs����� ���B-��q$��y�Cx��vI�[D ������|�����׳oOQB��G��l�?�i���ݗ{P<*�ȍ:��ᄱR���� ��y~��Q�AC��]���#e>�.=�����<l����|W�s�V���S��onW/��q�W+!�@�TB�>D���,-:�簡d=��.<4ΡcZHOJaXs��2�][�l�3�+�]�ʩ�초�ˁ���H�	����ҿl��sgF��Q�����P�d��J�\K�j@]bꇚ���ML!<�3ؒ#k�o�:���Y��-�<��0�nHf��j ���g��0 ����
�Z�/2ץ�8������81g� ���۔��2�t��X<��1�S��fv�- C��B�,?L�W�w��ZR��H#u,d�u���VL��0��Ƞ��R�WZ������T�>�)B��
�!�p���� U����A"���0��JX�\b�W�Z�O��P��-2�S0��8���k�O�/(�1~���R�l��~��"�����lH��T��܆�<����2?Eo�37ܐ�OiĽ�>&��U{?���7�3'c���a���|�lC`e�X�E��*s���ɿ�;��K����	Qސ��t��]f�D��<�_:_h Qs ��Ԏ]�M�qN`qਨ�YFܒG:'j���T�ay�[�����BΗ�H�GZ%!1ND�C�õ�u{�6![�@�dY$+G�S��	�u���<3(�l��7���ݵ^5r�K遜���6��.
��/ �$E���ݱ�q׌IOK�A,�|������`�R�F07шǎE��v�է��#La1}ֵ�@��D+qd�u����O�X�16*�z�e�H�����x�ח�p�]M[�V���ҬZ�m�#4�Ċ X��5ɷ�-�����8ߢ��G!zg� h�F��B�j���)�]iKޣ�Lk�(���5}�z�����R,7j;���nt��ڬ�:'M��{̡�2߆�p�j��,�9b��r�ΞӬ<$L����~�w�&�Q��ˌn�k�!k�o�Ib��zcۚ	�x8�����S����0V*=���]A�y��6*���I��k7����Z���#����F魵��Z�Y�G[��w9��
��Y����lY@�k�^�����Aø�p��[O��1V���BQi�������-/�W2�MM��C�M�d�4�����j���5b�	˝o$�2\q��ڱ����F6+���v�P�V��	�G�.�s3ܛ��̅U8����F�̀���m;�R1kc6��X�yn��9V�G���l!�P�����{	��8�5s�����i9gv<��Ӛ����Nx�\��A�SV�Ni�9y���#���o�(
�!Q��![�f�hO)�j��V�H_�v�jvZn�:c�-԰5�ֺv��<��ȹ �|j(��e����5����,X�jp>1�s;�}���"k�!����Y,s	ja�D4
����}�y Nz�$�؎��������͆�h�j��pG/	��u���2�����7>�&R�G"8������\�Mk�m��0:�X��b�I�;�T�X<�HX�┞��#jMw	a�C���,��Xh���[��ӵo[N/��K7���zC|�f ��3%N�Ӏ��} ~y+��NT�/W��έ���Fج�d�z���	h�R U��D~]�S�,4�@�G�=�i���5 �?��IY��y%��j3#p5�M����2W;JШ�,A:�G<�!IO'��c7ߍ�Q[��K�H$x��ZP�]��;ڃb�l�\q S���h���Ŭ��Xڸ��ڏ�$������s�V�%t��$�|��x�|�$v���,H@	�V�W���V���{�_����t�*�8C�|�#>z�M`�&�������ڻh��$��Q�7
0%�$# Ny�43q<�����7�W4y䕷s%�9��԰��IuMt�xV?�tC�Ԯ`�*CZI�H��waz��"�#�N߀B
�,c�z`�o!���~N�8i�~�%C�����*I�n
K������>)g �ڦ5HfD��~- @FX����W�)�j�I�U�"�pn�Z��)�b��Z�I4VnN'1����ȿ<�8���8�ͪ�����kA-A$[S_�'u��፜⭹��S�!t{jo��\�
�禐1���l'RCEAQ���d;��> e���Hb��/*Vã���;�WZ�������^�x�,�Tyњ�_4�K��Y�9qP�D`y�Vj>��=�1�P����ܘ�t���=瘊@{7�7l�Wn��+�J'`w�@�8���k�D��(���E�je�Rl/�ZS�(8q�i+��qt��S��ϝne3������q_,�s��͋�T�h�t�}]����\t%y��Z��Ȝܞ�����)-����T��Tj�����C�Y����G��I����k�*lK��H�	����c���ՠƎt�	��3����K&>��{���O|�ʳ�I�"�e�'��DM���e.+]�(A��i��-�q�~(~!� )�����Gl�^5���̯/9�$�5d�)�;b�uA]��jS)�Ů��"\B�o��;IL�װ�5�fsz�p�t�s����;Q-
����,`d��P�k��a����B�|2e�!m�s)>��аt�M�ÿmrz���6�%�gf��J����xB L�y_Wt��E�1tm[���S#�F�'��u�6��E�P�\�h%aw&'a2�T%Q�j�(OG\(5DNϛ�ё�� o�R�8���:��A�`��i�h*���;��6ț�	N��Z�e[�����Y����#��_��3����
���uB�ԫmd���Jl�?��?�A��� V?���>)�ӯ��?1��D3�Uc�^�<8��J}�"{%|VFw歯�+�>�r���`����n>""L~�H�e��24��l5K�����yI"*���m��:��b@;�9S�>�p�[�]�L�c�����Wd�����kQ�� :]������%Ȳ
�ǽ���4����O+��,t� �ј\\ub%��'\�_^�e��.��x��j݊��w~�s�J�օj�W!'*%H���ɶ�E	��V�%UqI��(I�|�l�r�����Č�WQ�d5�u�8��^@x�;GB�v���%#DNXv6#>V���u��O���O����d��\]�`~����X�G���X*�1�}�X��M|�
۰�╕'e��e'��K����f"5��m��{C[�I�z_��>/N��Mق]#��3'�O�� ��(���v%�����=����[������metyPS�6|�Pt�&��.�#�m�),��tw8eN��5�}��Eb�憃��h+�q!u�)����eL�	v+`�^�MPp����9΃6�%g#XtSe 7�=�`Ԯ�\�G��#̴s%��(]J��`�@<}��M��6��Wa�lȦ���	>�7V�6yp���R1�^�a��=��ЀaAt�S^�BY�_j+	�0 ;ű�®,a�	�,�
C�2�II����4DG@֨���'�-��ݻw��n�˚����(����s�2*\a9��H�iM��I�8�}���/"�s�D��]�����(W�"m@�h>B����aX#���-H^;3�:vwo}1l��oE�29hݰ����3v�V7ks;��lnε�d��JKA*��׏=�����y�gSpcn�$v�4m{M�O�B���ؔ������3�X݉�ᡰ�$eٗ��&(����к�BX@��@zi�9��9/��1<��&n�l���x	�M���dM�OƐHP�5�g�;����6���������!�ߣ������\��A,!����-Qy�y��>��v&6�~_��ML�"{bv�E����ϣ�}�3A8pk�<�"1��t|�Mɇ�S��Q8�f粧��DH�d)����2�<P��^�O[�p������wN���n�:�vT�KgښM��x����ZB.�#׍�h,�;�V@�����-Ǭ����K�	P� X��~�g5��J� �+EJ*���ȅ�C sQ�MO�
W�K��f��Vvl��רvm[ˮոMd��C
(� ?�:(��^�T؈N�碑��S�KFQp�N�%��!�
0=��}��ܚ����J����LR&
r�����9��R 1L�(��'�z 5��W�b�<��qq[U��H��F��N�&��ŸbdʷmT4�
*�xt$���P��-_�͖���~B��3�b6c�SnM�D��!�o�,��
�4���P�̪��{<�$��6�,�%HF��
���P�IrP+3U؃w�0��n�nK�:�z"��nL�5�d��$�/��3d�=n_�k=��xRQ ��Et�d
�7):�C����"ݡ��CKI��6�4��4 �\��/מ�(���#�㗣�?N/��iLp��ga��SK _L���h��Ө��\���=�	Tة���j@<*L��Y<f`�������,�Fo4d���&2Q��/��9��E�tV�'X�ܑ�ta�� e#}:j��GOw6uuo�s�������nӻG0��Z����F�8�Li��S/啼���l+�]�b���b�A����5{,qM7�C1�ݙ�vɹ�!��/���}���&s�(5�ѭp���V�&�)c߱�l��r.o�JF�oV��ί >8Nq�盗�]S�Z��:ǃ��L�Y{�F_�$6�!����V��n��z��p����������!t�0�C�o.�P'�d^CDT��N��׶rJ{�V����-?�� �8�F֒wh3�o梱�i�p��}z��2����R�&5�h���\B-×����	6�
pؖ愈���j����J��LI�+�T�iW����m�-�'&(m�K�)bS���4�AjF X�]��
�8�`�p�eW.a�C�(��U�&�{\m��Zן��ʆZ�n����#��]/=�ji�h}{L�����Q�5�!����R�?����={5����j@�iٴ5<��uGy�����L��E�AHB8��+n8���Li��G�cF�3��jS~�
�*5�s�����t��N���D��ک�zL�X��R�bc4
���5�ݮ�b4DO�>1n�����o1MRD$&�0��\�q��h�5'@6�gzn��"�g'�w� aZڥBI�F���� �/�1�K��4�5G���x�8[��_�S�����"y�"r�Z{ao�E��L��,��r3l�D!��6@Q�'�s�v~ϕ�<�4�<�J*YPӞ��VAu��'q�v�Bd�428�Ѕ1Qr��hf����o	Q^ �\�x��?Qo��U_b�S���
���4���g����L(4Y䎋J�.Us�?B `՘m�"�Q���,���R�{"���:j7W��pe�_X}�bHG:-�ׁWO���s����rU�sȖ_��Q���a;��*�7�U�OFj��bYZ�c<����QN~,C��θN|���!�b|e`�6P2��"!CH舍��,[�Lέ�<��ݴo��l�hB�+n���3)+�0�b:`�]��{M��
����M�+�##|�S��x��!���1�\�P�m�g���Ǻ�ʷ`�͟�]��s [�+���#��.��M"���5-:�\��	����I��:�T9j���Z�r�m�Z���Ώ�?Y}&Ó\������m%��OV�\�%PML�{aBӫW����$L^t2x`�YA�8p�Hv��k��6}�Ox?�o��E�v�Ϡ����$�n��$H�S�n��q� �&�6���q8����H�	���o��83����b@�n��bg��^�ul���~����/o�����J �\�bNb�N 
��n��D�4����s?��|���|XM�Í�a������e�fg@[h����:�i`��5���q�L�`��?Ck�G���r��lB~l�[��֋���<I?x�;y��?�'�*y(�h��a㴪9����`�2�pa�*P�����F�����`���Nld���л�.���ˈBH�a%,$a��R�lƱ�]g��B�Z���őҢ!���洓8����6z ;`��jZ.�G��,��v��۵�m�,���A���#kZ����!U�� �0� ������Sb4/-�3�7�S�*8�����I�~ezna��O�s��͏cq\`�pgj��;�����A /q���\�9e�~��x���33�6���2ǿw�
8��հ�윆UM��dEg����ߠLw" g�
�Z��,w.�g~�WQ[:�S�Zm�}��/�g���y�_�p�<7�k�ܕ�O��Z��s��c���>��<�Т�
E��
�͐�Æ��2;7�H�dl�c����!��_I}���z� gV�r���ty�up+ĳ��#����_��|�~vr�����pq�#,Ic�o�߸���%o�s�c;nC�J Ӥ�H�K~J_(\l����Ӽ�}��Zkg@#n�~�G��-/h̡0��<~K���L��D�<_3Ί�%�5�O�?:������2$���(ud�@s�n|+���r�����G#Wi��`�殮S�|A�!�wiL�����O�ut~z�]�`��s>/Ĩ�@D�U#�Pv*rG�?��(U�Zj�VҼ�;:UMh �
<��@�E���ޣ�y�:��ey�^];-,��n��WW�Q�3�Q4E(��ZKy��ݦ��D=~�L��Z>�/��i���G��wF��q��%f�V�E��&
����H�>8�zA�"��c��t�y
���J�.k��J}���v4���5��P^���-!��ܿ������<N�ciVw�5�ؘDϹq8cg#fPm��9�(��Φ (����y������Ӝ�T;b7��f#�'���1��J��8w�΀ҩVO���F� ䷎%��Fm�l������&#9s~��E(���[
EP���c�n7yY�M���8��y� ����1��4�zq|϶��9@�d8�=�g��C��t_Vzlɺ�5�Ǝ&�/�T���a��Fa�K�I��(���Yh�`P�&��č��	 D�Q�����,�"7� �u�4�-֝S�@5���.]�_�E��q:E2Ss���}6��k��%§(M�n�{{3�o�G
m�|o�0h�)�7Q��3�m"�������@��:����A��_ɴĞ�ajZ��Vir���/!���9�����""�Z!�?��A��՟S����
��U�����_UF����H�qtr�K.�w	��6��j��m��қ-���|�\���r7?�[bc��_�!���>>'z�N'4G�$�NQt����$I�V�Ў�u�)�o��'e=+��zV3��	M1TL.nͳ�ߵ*/?�R��:�B%�Jk���N����^���v`���+����������c+����ˠ���q7s�&���a3�\ps�|7����2��:�Y�-�[�]�k)+.)F<��li7�$�UR���7��Am�<��!���:y����m�����/_���'����K���~���U1����cu�,�[Lm��e�ګ�Y��X���=q����j��:c�k�S���)� I���7����'�aG($+��]Q^�����:/��b�T.p�W��e��$�<U�ǣq����>+c�L�#A�L��`�(1�� i�5���|H8P�JQ�x��*�RQ��:�]DҰ�����ϋ䜨q볈S&�SB`��ih��Ǟ��Z���:��ߜ�Ì�>HY�#�F�fY*� @&C�?��& `��J�
ϕ���0W3�5P�W��U��Q�d�=̛����'�]�R���$�n��Q �>� LJ� 3���\���
h��&0A��rЂ�����Ŭ)���%�1͖���~J�!��Q�Օ��C�I��Ogqe�dI�*B隣V�	�u�_�g��q�W!2��}2Gw�#�:���U���[f�������8��W�t��,���W�p�h!�`H�����J������8�.L�!̪? Z���nV+T���u�M��;X�5g�t`��R����&>t��쩬Qs���z�s�e�fQB�df�;�S䤷'�U.�m�b���}ZN��ޡ�Жҡ��Ie�ԥ��[?P\a�#����	�f��0Y���A�OΌ�O���W�]7k]�9���+��5�=�)x�q�e4�@��D#X�����'�d?�K��#Y�>��\
t#�"!B�X���c2�X�fJ�'p6��x/"�0N~��&��r�k�N�
�R<��^�cw�����.yw�%�<9Va���<2X�3W��}+�ޟ{��L��o����S��f�¦���'94[\ʔ���<���N�Q����;�m$n��)�t��Bp�`�Lc����3�R�\���,"�K��PV���f����,C�:�4�|Bpn�:��q������#�+X�e~��v9�B_� ��z�kR0���x���%��ͫRw�M]����q����� �l�P�Ei#���^睱3�h�3(�F'�����l��)�@
0k����zj�!�p/"wR11����(X
e�I�w���v(~s�b��4?n"���𧻓{]񭎢��|>�=Z�Je�=�E��`��;�12�إ��.!Xp6�LII�@��/�}`����۝0p��&��Ў	���`��x2b�i�"�'���O��˒�s6$_X�P���<P�q@_d,��O����3��ʲ$_m0�~E�-��1v+�FW��� 2���VZ��DI�EF�n���7:���p'���/�g�ֱ`ӈyR��);�NJ��Ѻ$���]��$#�ʘ���\��9��Vpa��~�z�;�<i�h���T_�0��}j eOK2���U���0sP'�Eu�y�KC�BJ�ӿ�v� ����y�����AH/��P�b�������kt.ֹM��T���ޚʬ�����ϝ�d��,��Y�﯐S)��|В��9 �D�lTf93r���E(�]?�7�ƵX����$��!����_>c�:�f��:�Ff��3�>L�Ĕ��vl�	dL�T�U��>�l,]-�������\���/��U�e&�̩�i.�?�� �l�t!�?���-���X�?VR9�]~�h���YsJ۹Uݣ�-�`*��XVK4���q�C�������$$%�c�[&�H⮸"��|r4�?�J����Z~�L_�(���	�)٫Bqf!gѳ��oul��{vvރ�������;���l���Q|A*�C�ld#P���ͫeܽ0��@������OT(���X��x�H���[�H�����l�.}����*q5�1�p�c�g{q��K�1)9�j�ZcC9	I�\���l��k���}�s. /�kJ�-��8��1h�҆S'g����:^�e��{r��z��+��L�����F$�x~�{��]qkcQYm��r��Y��[��Э,~�=�ycn'Dj":����iLYBN�a�}��IS��x��8�%}�=�:�>�����y��������YkpB�cd��;���W�J&�/�c���4���g'	��?��>-|�Gk��1���ǎ^�2�g�(�i�\�.@ÿf%���tf�p2��D�@�����^�J��7�|{=�U1�WA����~�X�t紺��5�k<�sh�y
�)�W�D��)�<��;��m�H�\E�M�+2��%z{�:�����2�Eh���C[z�&-i��'/5�����{.��vd-�^���Ó -᭍�IQ^�p�,��}��V��<c��m��JU׺���绷 T��K/�������0H�΂�ڛZy;̞�DHbZ���:d�b����H��ӂ�-���'`�¦D�8��������,��Vo�o8v������=7r��T$���lC�����gD+���5,Ya@m��ҽ��ͫp��[�1r�-�:|��%M�iEC5�i8���6+�¡�Y��h�"���D8c��������ɼ����~]E�8 a��h~��6cf�o�Z����\F%��Ah��r�Hx_='��wА��i	W�z+E�p��7�����O<M��!�����'$_���]�l�d��W��/!#��A�M	'�$5��7[�M���F��2��6N��2B������w����)	�.���@�c����ڟ+�ɸ81r�􊏢��0���Q_7���q,܄\:��)3i\� ���	�#	sLK0�}\ �c�or�Q��F��nID��ޭ����y�Ld������w����R��P��S����\��|e�xu�/HxC&�>��*����|@� `�H�gQr�l����	p�<0^((iU�&
�ǫ^��M	��/VAi��`74�Tm	/�n�OL��7Q��k�
 ��ȯ��,�������e�Hk�P]Ip�������NH����;�&�C73a�H�O�|^O�.y�0L��E21Z��&ύ�a͵��.���o��dG���T�B�P��maQ��q?U��oԵ��u�x�J�o�I��7��c��Bh��ǖݿ�^G7��YW|�\�rM~�*��aa�f�FT��Ȋ�Ӝ+T�ʘ��̆�7���[��)'H.��!o��T�43z���1!�N=>�9��J;�zb4/��$�޺3��2l���	����q15f�X\��i)�܀�|�$/�I*o[� �(�W̜a�K'�z�f��_���M�Y��{yU'�P�:\1'�ąf��4�2�F��gXMv���NX=�A7[�j5�T��uOS�_�x=C�og���V{S�2ۉLg�z���</oP?<�ė'���\��.{�ʃ�V+`Q��EW�[|�uܧ-jٖ4N�S��z_���s4�O1~u�Vpc�n�������l"p�m,�B�+Ф�����{�L~�}Y��G��!]�K�f�Hu59k2/��P�З@DF4��/�t�1���?6=�2��I\��ˣӗB�12'Q�c�nP)��'P-�v��`Y��_���s�μT��P>��p�U�������M���/ڒ@�j��4D�G��*+���T�(yM�"*�'��d�(B"�n �2C]c�Z�zSDB���ҧ6��<+�|�U���8uf��j�
aD���h	隔	r���ke��J��[�h�mT%�F���Fc�ҩ��O7d$�4Ee���i�r�#�a���}N�i-� ^��˒�7J���bSbr\�������
Ik�Э�^����hƯ�ԽD�P�c�Iw�,�����-��S��$8.���w_�t�_ːb�؏ے��E�rC��kuN�W��/[{�9�q,g���Ԁ�)���(X���ys0��iqq�1�ȕI�^$ȴK�.�fr��;�	٣�҄)��א	���wM��|T¤bR�U��:������&�����\=�e�@ϫ7�6kW���xh,@hq��ø2Ä�{���I�]�]Ǽ�S-��!��;v��&|����m��X�hL�c|��E*�,#h>��xh: �����,���z�/e�,AF��s�G�����ީ��-0�E��,h3��P޼
.^����ß�'��}�q�'7��d:O$�Op2O�&�b+.'C59���f�*����?�t�u
Șf����5tR��#�Q�!'��H�&ycR���X�}1>QeS�Z�~���P��I�? ����d�'�'�B�m�V�$�@$��p��FKQ����}_Z��Ņ�\�nH�/�!�u�Q`h(Yٜ�.��k��㡯����E��7�{�Y~����K.�\�<&M����8Y�ٗ>��*�x����gE����9��~���K��Fj�uKb�8�������D����IU��^�����5#��$�㓘�T��E&��^[A��Vbd3��u��?c�e =�A�с��8"�m$�Ծ����O!����I���iٲ�_zT�:� Ig+ӥl��s�Ƥmo1axһ#H���K�I�%kjl�p�)���)���C���qC�D�c�C^e��%Sr����[�B*���ml���d����%TL!���H������T���:��j`Ru�q;m�X���|@m���'(6+Ar����њ�[�Y!²�CQ!#^LXYxU5^����V���&9�����C1�$3�Elc��ި�Z}t�z��*�$��:�W1$����������d�>�5�Oւ��h���)K$Y���2Ĥ=�3�p����_[0˭Ԃ���ڶ��6߆��E�z.��Β/�f��j"�!�Ox~~_��s�]�M^�w ����o�>Җ1�wF���a�$&t��x��+�8�x�İ������@j�X]�O�����t��0�^2���s���INv1M
�+I�����p$�Pus�BJ�l容W���	a�T�i��Jݬ�d�|�ϕ.w8���'�x��Uǉ{៰�8Z�����ˇ��������aҔ��$�9|��Ô/�����Z��z@}MK3g��r�G�*Z���p3�.+��"We�q��}�*���Ѭ&�My��=&�J�O��)��|�3��.�߁�j!�t:
�>�H���L*��v�䲘~���i@P��6ZT^%ջq'�`NI��,3�F֨�]��.�A"U[zr����je��*��\��9�*U�7�tc�B����2
އ��x+�R�R;(jB��ST_S:��U�"'�B�][d�?��Z��U�W>�7=
���XO��9����"��m��'�}� ��k�;�{>���;x�4���T�/C�-�G�7d�'�����.��o2\2��l�ԟ��ҽ'5 �%�s`Ȍ�����h�$�����;��L��=��G8�&ˏ�BF�T��%�p�
$?�vR�K��U: �b�a��vQ�[Ʋ3���%{������^���#����^Y�G����ꐛ��k1*o.��oWȈ�����35��C�/��_�N��o�D�Y����!��S�'挕5�a+l�.;�շ \R?��|	��8���y��u�y�D����b*��~lzb�Sͳ����W�g#�D�-㻒�1��Ty{Q�,< ,C�ݠ�N[嶄v�I�q��\���;����QũÁ3�����R�����mюfZ��G�)u�Զ�u�
\'S�׍"�������?���:u�wqB��S�]���$4)g�(��r�E���{�U��'�0��:� �]����HMr�U0�'�����a��	GgȲ!���ơ�CL���ћ�f��e�L���Vc	�Q�^�"�p:�![��h�"�}�� t���s�ڷ����K3���-�HO��Xe�>{����a"�	��Y$*����n��S��|wi�+�*�)�Wk���rI�xVaTX;���λ7}��?jȚ����૮�ܠ���}#3$�r�{+_�O�ڧ��)�ɖZ�\"%�m���3�Sv��N��� J���Zx�&ļ�}�+s���M�{�|糑;��_/�����ࣛ+E�lO���
�P�?"�?I��J�+���*}��q�/�	`��uCM|m���d��%�˪\,�vS�q�4��_��n��˓	�F�'���OM��UF��а�~����<GF�Jr��K������|��=[u_=bl���(jF��D�����p�����K���=z���?���	ȯM+��2J �cH;r(���0@��QA��Y��Z\wF�Z)�bf��m����.�����"���w�A�wՌ�j����1�+E����H4S�C?�Z��r��ì�I��v$�Zf��c�V�9^k"����l���azHb��Z���m/���/�
��5�jx#�[��?ok,m�]�A����ס��W�!��3��N3���J9�
^��|�Y\EB���s���'~�Ѱ��X�p~�a¯�;inei9�/ˮ��$���{ƺ��v����nk�K �z'v�-�nъ&�ۜ�p^���U�V\茬���L2޼��l(�`��7l`��-%�)1�m�Sak���;�)#=ڐ��3/�L��4��@�?���
��,�!��Զ�;��ۥa���\g��}��.�s� K����:�e�~�Ca?[]�����06�5g�d���8)���RY�ؙ N�K����7U_I�������V�"v�'�!˃<���`\u�?�'c|�u��&����*�X�X�f�Z�5Q�L(]�4��P�!C��v�t��68&���~��z�Y9���A|�2Mij�:i�<	4��CF唭���[�ly�6qxV�͉��3��
���������E��P���r옎؎ g�fN�C�y g����{��@֒ܲ'����%|2�SE)M�t--��a&@��X��������eN�d|h�Dp��>�U��V����f�*�� �2���SM��a��=�ؑ �1�n,^�	��2���&"����V�}�Đy�CPBULO�	㫰P#J�ѤW��F�(yx�I6q�i}���"�bHC���a3)C���9^~.�&��2oI�[�=�?�[9|���3�S��_��>di��C�'�z�u��ka���H9֞\�\΂��Aƴ�.�Q��z��"N�5JQ��}�Qi��Sb�,*���b�}R�A��D,	����EfbS��J��)=����dU|���
O����\a�.C�i����� ]9	,}��Ui��ܞ�A�9�Y�F�g��x(�498�Ҫ�J��_���ᢡ\3Ӽ�%�I ݞ0�cᖿ(}�� ��Z��� ��[�����G���1l@8��)3�k�戧#���V���i��FZR���D�m��C�����-ٌ�'::��>fP�isM$� �)��4��LF+q���^X���U��2�K�1ֈ7;vn9��%��=�oP%��3�]���Ș�P��#�6���_s�=~�,F{?b�3�Q�LH�N<�̉e�_�i
���~@��t�vB+��J�[�b��oI��3����GF�3P�x��OX�7�C�X��C6��;�!����R�ń��"���+�]����u)�P-�͋HwrR	���uf��Ť�.A]�=�5��|�g4Vۣ%	��-�����uy˝*�c' �if�oZqqs�R��P����Z��s��̖3��oi��d�?�F�
XG����J��~զ�g�Qe<~ڙ���}��J ����w���֚�ק	���S�F��KW�矏��yRB�|���/J,�Mrb\���Ē�
�Ȇ7A���r;�`���u�3��jd�{�kZ-�c���]�?yGE��4��C�>�������=_�R~w���K��D3xғ���8w�`���Iup,��<+!.�H�\$#&�v�����a<��{�pY�z�����3܎+�6�B�+b�uϮn�;��s�5������z���=�3�l��Fj��<�uK�t�Du���G<�0c��Ւyy6�S;�U��*3�p �EBL��
�F� �[ @���tf�T�+4m��W�M ��ֺ�Wݩ�D���>?�?pzp'�P{_����<�P���)��ZM]S�p»d *}kѧ�Toւ�b+�z��f6�[v/�/wAn�j �'�������{c�?ӂu!;Z-&_+�h� 
�LVQ���-�������؁l�j"R�j���	#6�qȦ��om
��=�`_�G=�x�H�|3��"j�N��d���/��T��HVѢ
B��Ce\:J�`1�P�a|���lc��M��um\�� pT��fdC{1W�ZІP�2�Λ�1��*������±U���1�|`S��l��Jl�7�9�冾����pQ���&�iΩr���'����nr��.�t�ЅYf�S�N��^�[�G֙�q����p$0�xɓ�h��V����o3Ot��S�|�pA��jjFEJ��<���Q��^�]ʤP<rw�VK���!��T��iÏa̻�P6��eQ������T�3�6C@���X%��+^=����{��n���>Ϩ(+��3@�w9D�9Q@���K��e�N���69�]��P�����_��t,ML��D���ػ�I�Q���1{���]}d���׫z*Y�E�0��p�5 9�v�בV�h�1��[�3nƍܴ7���<kg��g�D(�MO�2��k���~:�R���a�:z���D�1����0������$N�ޝ!��D�C&���S����%������Y��=G��i.�۩J�y�����EC�(:��~�|}��Y��Ɇw�0�Js�h����9
,�I��b�޺ �Q�G����E��ո?�o�7����1�,�+D��D( ��B:]�����8��ҍ��J��M�{�
R��g*�Nk 2�S�S&�d	G �'p��2a	BQD�R�P���1q�G�~0+~凶��^T oi�O�oW�C	���/��YR��j	|����S6�j���m�g
$"�6䩧p�m�o(�cC:X�t��7���1d�������7�Uʽ��J��8k���E7�6��ܮ|��/�(n��e8-�y�.��x���Ҡ��x"�d�層r<�o3
ͻ(�B;'��$�nB�y������ ύ.��{�y����U���o�eUOy,Y���x9+j��1�M�0 �[�NFf�,Ǐ�����=��K?�6�I�)���
�P��.E�نB�f��7H�blY��pЗZ�;�	�#+��n/�-�?��#�,)��k��-� ����k��ܠH�&����a��X2��0��ebR5�k�LV����BYP �:qn�B��,��sã�/��#���l'ij���ψ�X=���O����e)������9s[c�i�:w��Gr�et�-v<��tm����B�:����|���}������ݩ��,X�"t#ظ��W��0�)���i64{:�kĸ�8M�����?p�r��5�K���ɓ=�fݏ��@�,�H	5�g&~P���38F�Pmկ}
���͉�źs�`I��Qc����zp;�����y$�20�0�8����5���Ȏc_
��d񟇕���P=�wZ%�ig����`P"R+c96t���ۧ��Ho����L�+� ӆ�^������]��u����Zgn���\���HmL=����V���ㄉ��؇!�FqQK7��_4��-�
�����V׭�����i�Ҷ!�du�H�'6���1c��<b��j|�l�74�\?-�<ic^y�GZǤqY��(��]������	��~���r�ߏfӊ��e`]�Z�@T�l�'�Ξ�o��R�_�x����jajήC/�O��sDd����9��\�d��O(�q9h��N/s������_n9@wT�<(��ۢ�r�L ����A�h���Q�[��&b.\��Ԍ?-��>$�1D��w��+�Q@V��~d��<�K{eB�ƙ0���M�8�"��)3^z�?���cE9~���Ɨ�d�`�$�L�ctѧ�Ev)U����8!�$�)�4~��|~��
OЋ���r�;C�ٷ#�ت��u��$������{�&�Q�{����D�|F�?gL��Z{!_�%�&^��l��\˴Ō���d*�����o�g�l"b-[������ro1'T�I�-8(�>j��z)'�E�V���������#"'�C<@5S���-%`S�:JBl�MGT��p��ya�6�t�뜭dE�w�%*NK84�<�T~�)�G�ͬ�Pٵ���8�DB]��ț���#	5�F�a��Gʤ�z�q�Iqֵ������|��ec3��tқ��&����{u�����Xj�mtqz2�_|�ڗ����`Q��]|4�!�oGiNj� �M'��\�ו�i���c�A����qp��6��:�P``S�{����|8G_�E�⨣�Չ�>m-;CQ�ʄ�ɻ����L\�8��g�Jm/��w��ZA����"�r:�ZA���6�?��h�1���a�	���zO�ka>R�Ć��3Y��th�V�E���:�قC��j���d��y	ଂ��j�1*z�8�js������xg�6i=��k��7��z�kCd5������Å��t[����y59z$β����z&!�I����lu�ە+⡉�,;i��7�Y���K�Xd#�!Аq�ZSy]%0�p$G�(����5���3	Q['D�C-��,�:���UZu}LD��I�������v_Tdi6Q�I�FFn�#x�-Ñť^%�˴�}�lm1f�iԼN���I�?w5��#Y��o@<�����8a�XB8���=i��c|�>�0�pJI��@<��X���5�kl�-HʎK���l�+��?��TT<�L�Z���i��{������\�����l��.z��W����
�ǌ���ѿNw�m�� q�΍�����Nd���eY�-��Y)ʒe�}�7iOT�)���VEj���}�N��6 ��T�� � ��M�"$� w���=Ƽ�KqZ��`���{*m�醈�5��ǿ]h���gI���6QD�6H�o�)�8�'~���}m:�ɑ�Z�L�#/˿�kR�B>:��h���c�?h�|�V�,���I���ȃ�o g�+'R{�!c1&=O��5V'dQˈ�����h��7 F!���^��3��h�9��912셝{�X>O*k� �2͸���X<:����ۭ�Zc��Z݆���vܬl!�� ��M�%$:�"?s�R2ƍ� �O'���J0^{���E[� k�T��D /�U��)-�O���@wY��k~��q���t"��,�j�`���M�WK�'�Z���5G�<��z��6���Z��C�V�>����~���&�9��G��9�S�����ĂQI.��	���l�g딪�Q�۩LCf�~�-{)3	�ն�s��Ws,5�G�Z�����P��`P�~+E��F��:OG!/F��+C:eua^��'�g�0#��4H���ɌH}o��Ã�]�}{*7�p�b��@glt��U��z�X0�èL���'�i�y(_��� !�Éꤱ�d-vIa�	'Ғ�a��ǉ�&Q�wɏ�@����ڸ�	RqP�:�.��K:#�S��3��C��O��ຠÁnT��<�l��f}��;th3���;w�Y���$���k[�s"�����~���Nd3*�P�L�0�,|e1� �Y@<}�4��)������G�D (�`bֳ{b"�s9�9�����I�����+�Z@�٠�
$@ -�NZ(JTN� ����+���
��N>�!� �@*��W%E�%V�00ў�r��;i�X�aY�_pU~���AC>F��݀���e`������c���{c`C��\�N{�z3KN%=�ձ+ҿS{2��)��3��E�0E�����������z�\H���"g�xq�Fk�WE�Lǌ��k6�8�����Vy	�=pO���P^E���j�sH 'EP�bF�Nl��>Yc�WF�,��G�K�Iy��r��y��r��F����e;ä8W�B(@��P��ur~��PY��a��7���b�f֪m��C�d�̊�Ʒ<3���V[�ak�*�a�6K�r��p(��r�i�P�p��	���
iYe�.��B��<���*]��DY���sܿ��7O����,I �Xz��چS,�R���p�օ��k�[FA��m�mU���D�Jv�b��83|�#&��0�u*�2*E��E��])��[b�E�pH��y-�k�����dwl��,+O��Ś�تP�0���,�[�Q`��жl*+y/�yw�`�	����L�!]�2vy�r*���=��{GC���5m?��N	�q�&3R�f3d!ժ�(�M�W$�sx��b>�Mf̖ß*�z���F�8K��㻕D0HpsR��R�
����H�Sol�"�̕����V9$ⶓ�W���h��r#���G�gF�J�2U�.�����H�`�P�\�أ��L�l�<c&1V p��*�S
=d�4E�kψJ?��@u��"㸔���������ݺ����ks�������jm��x�-Na= �'�yXgb�g�(iiV�8�.���9�14�����S�ȗڃ{��ߵ�`͑�u���-w�:D��Tls(��1?<@�2�j����h����x����G�ȭ&�o����,z���a�*7�h�E�%=}A���߳Kb�JOeI�����-\.݂̦cE3Q�I5�X%G^����V�eaS�E{��X��Y;�_�vRy�ݿU��ݻ^����Fl���=0w����C��[x�O�����P����>�c���.{?�R!z�����M`@�N�,�Oc�=ch!f���Wܦ�	'���u&�E>�l�7�V����|�g��#�54#���8B
�]���{���+K�r6N�S���"�94�`[��������`h��
�O��e9�ڂ�O �s͎�1�����Dk��YE���G,��I����U�-jli�;&3EF�*�|	���B�� �z�fN$��-t�
�I�f���OC�{���]8n	_tt�hiG��y|�ߔЛM�v��A�Z�SU5ގ��UC��ձ\!�_��h	��7��[`���
>����k[G�]���T���qN�H�@�Ԙܷ�d=]�[F��I1	�*��q��L</��z� [������)g�B
5����Ix���?/=�J˟g�A�����dK����� 뚞)L5�zj`ԃnv�E)�����Bjvt��IA
`�<#��l���a��/�9�����
�I�͍��A��'�F�(^��\��I�Qa�T���ꗋ�.���Co��o"�P��(� �E�~�����{l@��]�g��}x''�D�zB������%���c�m)�B��ZS8��b���1Ȝ����D��)6��@�7�[w�r�19B ]����pG���f~Q&D�d�/�S0���j�*q��uP���-,�`�����;�[��c�$��ZQ�W���g/U{4���r�#2 �~��N���ҹ��!�F���<zZ�O{H>���W��k�O6�x-�	��s[��&!��F\*0�uث���ta�����规���9���VCy�f�� �q����`��I�=�~*L��(!�����ߌ=�G2(Y���$��~�5���wl@�tT<!��<`���-'ŀc�U��ޔҷ��d�"h~���t�aB{5��N��A�Q��*�8N"�N����rA%i�D;��Ѵ����2���VoK���m������Ff�֎V��h��B[ۀ�>�Gz#7ȝŔB%��|} e�"2;G�M� �x�����fيN�[�5��;s�
��F�ݸ�����{�(���� @��2�l+�ß�u�x�,	䤳��)2����I����s_��&+|��9Qшh)Z����ͣ�����ܧpG֝����P�e����n堣���i�SA�i]�G�L�jU*bX�oI��S �et�dg1�(J�ڧBP���.��Ǿ�}��F��h�،�LC(9@	��U(�f�>�L�������\
�%���Q$���p������M�b"U�nQq�O�1�����c��XY��Lv��2��cx�!*�?)<�=�5���4K�E��RN�ղ��(��L�<�~����?��/SFZ�V�Ӓ7v.a�ж3�<�ع2#A6�欓����S�-K��&%#0"ѯ��<nz���=h�9[��i������5lУ6���&\[�P9�fz�˙����\�!� ��jl�0�"�"Ѓ�wZ����5�;�Ì��7��9��M��ֺ�u>�0��m�
�"�F�un�EEۯߤ,�j`����JQ <�rJ�}��'�Ȭ_��bVh2U�0=�p����9ߏA���Z��Ϩw����F)d���cV\2��
:�����/����K=^*�I�NM�|唵���m�>��߇�G	��46��sp7,B��z���0[Wa�I�s^N~B�j�1��5���dE�����O�_e�$�l��;�챃_��Dy�x|�_{���rI�gE��^�,p�;��Ss�=���r���j�s\�}?j��� Ԣ0B�$2�!I	+�*@�#��<ﲾʡj|��yvd�y[SC�J5h6���'�U�2����m��2�+N�����7shs���E���	,������_�oh�l���H��}T�K:��X�@?��T̠=��W7�R^���D��[�so �UrtZ����bá �%�#�7�0��J/y��L"n��*���"'��~Ϊ�p�h[t�Y���[c�6��q��7�/��� �]�i�����S*syx����v#���%cf�<�j�}'ߌINd*t4�CT������#�d��%�r�� Hp�����$m͡>����7�����޽���k'��VqXQ˻�zj0޵�֢�h��ߟA�%����B��t�SPFu��[��.=��a��΄;Y��8]������?u ٙ�ٱ��7�!��iಟ�1� d�8q�Ͼ���τ.�+�"l��TnP2/�w�QuW��ǉC�+2B���+���&m����l*��|^
t<��<?�o*}_�O�}�S�i�!���u�~�j�\�v�8�4���Z�b�����a��	���5Ncf|���� נ{G�:�m`�^��-L��|H��	Z�@{B߶8���)f@�v�9�O��Z��gZOaR[�tvL�/L���'a��,�D� Įy�@sT�qd�+��������(a���������9Θ]�0�C�=7���9�SU �T
�I�C�61d+� cl?��fx�k��f��]eɞT�J�P1f�:���|��f���Sf&1XB��N	�]���[~�����Fa��|� ��!g����il�'A)E��y!#0.x�ݒ"���m#���s�����2>�p�қ�5,�P1��"�rD{�7�_4����V��?Yc?�M�R� 4ti��"� ʷ�;d���zѾp�v�E$�FO��[��@MbC����Sb����N�쉉V�%�.rO/Ͽ�0�BMa����L>sy�e�p�p���2�B��� }FPW]i��5	��_ח�E����*o��ü��y't2[M���?ؽ4ġ��P@�]8�-m�e�}4�E��Nh�Z&��w ��yǽI�H���q:-w�W��j�w_�D�y,��!wq���[�xF���ggM�J�i�y$���M{����	�un�
vc��׬C}�|p���xP粺��8@�R�z9�H�̃l�[��Z�Gt���\�6c	�]�Sn+94	+����$Z���bi}'X|d�3�x���Þ�tr
�{�F�C����)�4@���hƛ)�@�<�r0���d�뜉��L���1"@r�����:�>ی�z��|���̛��c�VuA���������)+�\�����%��O4@Z8P9��Yts����lÏ=���U�p��F,>)�Z�9�毟	O�P����y���a�E<К؊�q�Իb'��7�ǕuO�6gD����w����wؖ�Oj�U�������ӹ��?؟�Bq"�]��!5�4�d�:�N!�}8���/Q$AW.�5�z�7Ɛ=����� '���s^�d�QZ�e�m��[.6f����M�����q�����q����נ<�~��QYܨudp{�!|B��
ۃ8Y/���75Q��-3G�v�|�a��� Vr� 3�jֻ����Ȭ�9�x�8�NP�O�����ﲷ��8�4��<��v�����Da� O.ZP���E�m�T(�-��4�
H,Й��"�(���A{��.��;I)�4��ؠ�������06<��3�ȍ0N�.>l����d}n�R�Y�M=�}�y̩iQ���V�I���m�`�e�b�RG����Y"���F�L+��h9�r��ntKOk�[���vE/Ͽ�~Cdp�T�hW,��t|�0*m@M��7!�������'����#48��G�텝->v4���\0�V舛�a��d>sV|��M���آ��{VG�����=����~o�n��� ��
�8NA{�
Os�贯�c�m�u��bUMx�0�m�Qj��g蝄�h�^�[�"ޔP������?�lMxIV�p�+���XB�����H)،R
�w<�Kj=t.s��B�@�4�;m$
^<�u���'2-�CU��>���E�\:${n-��[R��Ln�âoLJe�$-8YR>O�^HX����߀:��@͸����*�R�Wo��"qĤxt�|�k5�-��&���"�a�n:ԏ��V(��X����f�f�VZ�n��5�
ff�)Z���B�J"�O��yl�:���Z[������\E��w�{"�o������>^��(zf��@�_�OA^��9�L�� ��2��{ߏk����V�4+���L��p�9Z��"9����h�O$o6cu�*�q��{k�$�He�Evd��EY1k�?&���
�~QБ��e�,i��s��E/���Q��PtM� S�R��y�?�:�	�0�V�W�Τ���D��Ѭ������g�F?#����rkB'r�a{�D//۾��r\M�z<��35V����v�X&e�L8M��B�b�/�m��D}��ZR$w4�&��{�]��}F^ ��Uj|���h{C�Eb:i��Ձ7/��.|bߩ�hܕd����ma�3�7%��'��9�&�i6�'��8`6�Gu@5��}� ����L����A�7}l�$���6dX���x�r�E�X5g`�0�R�lD�鍡C�Ź!��uaL�p}0s���/�S./6ag��M�)�8��U�n|�9��oj���g���8V�$�w�K��M�J��`���:~�U+���~���;��V7{�`��XW��I���Ƣ�̨�zoޞW�@5~|vL���:�4wg&yVM�B<�%���ۢ$c�D���A�&�.{�7��`�Xh�d��Y�U��\B޼�a@5�
`���VC[u��6��mU�$���:H���8Z3��"�=��$N��"E ~���C�pHb��l{�Ƌz��av�V_-��T��a2��,�D����}z!���_�!ԉCH͆u߁^șL5 9!��XT������'*�Y��~��m�[�`��m���*���!p�O�6>M�U��K����;���<n�\�IV�V���|�?oޯ*�w��U)Cҙ�cQL	_��`��/���i0�:��<���&ţ��0p�m�\�u�2�1�4��`5�[<	�ܯB�w����aB�6�)����!'"��i�R:wX��� �Y^��I.��K�$6�%�ܭQ'��{d"T����c�`EÓ��n1'�;�l(MY66!��\�V�2d-�t>�t�����I&��h�;p�ռ�H;���h9��B'�!�>{��(1r #tc1-�h2�:�[��>�}Y���NV���8�U*����ta�����y�"W��d�ŰFH1<�c�m?WX��]���p�q���	�l/�a�E<��8=:Em d8ݐb;L��`T��L���䆋��ebA��4L�ƅ���sc��uK9t,������r�>(�v��#��ӗa)*b��L�e �@��u/��N�t����[�7���J��Q%�'cvAߪ�'��OͺE�S%�iX��s���<R�k
��#������hyB������AOD�m@nK|�0��hS���.n�M�J�g��u-O�\�iYfݮG�D��Ȕ�l�e�y�Ѝ�ERy9)"D�ZӖ;��s��<^��gzwyQ%U@���a~��7������a�+n��嬶�x�<�PKP��t��:q{�M��/�:s�������ч"��c�[�L��˘����OK��
�}�85	*v� �?�)�7ـ�����J�@�א,���T+j�4��+CQӘ�#�'� vq���f!-�1j4pIGCb�:��8�k���'o��8G�%	�fXop���8��~�'"�}��Z��	?�o���Kh�0P�-/,��ib��=��$�>���F'Ї��|G�\�QSd����#��w��g��ߕe�]z`K�~��Q���@���E�}Ԁַ�Z{��v�no^�������	C�NἯ�
;k��3��O9�d�g͒}I���1����	��ZRm�ǥ��&m
���a�$�Vù�k�v�����YM��ٙ7J���Rt�������}�?�S�)�@y���cbI��5�����Y|��=�SM�o����s.��ڟu�Q��A��Pj��H� ��4=ժ�6h��NZ��*��g��e�U�Y6O�����s�u8��"kl_^r�E�@�����z����,m�C�]�L�G��5C~��Bx.�F��>� �Cl�P7�s.��ڹ�13���|u�u���
�M�$�H|���(������+�h�a�Dj���\­0�����;/�gT�n-2�m�z&�N�f���	3+��K?����T�Y�4$�6�8,#:���-��!M�z�-�l %��r�4*[���	����HE��X֞�Zt۰R*҅�2������:� ���'f�;ӏ�IYd���4�{䟼 � ��q�pv�mF�$EB��O�MhE�a�-&_�h}L '��6��.�nM�q�!�X¢EGW�N���+l�F�H��W�F��d�T���-�5WLT���n��
$E��/��Tμ�U�R����]��|ܔI'�~��%\,;^���6��q����.�� Ե�MMx=�W�=��E	L�LS?�|��p
4N9%H3����R�2J+����;�rU�[��f�S��{�����:M�?�Jn�����]�1��G�����|�\\��^�ɘ8'�[�w���e�-�&
x.������Q�e���YK��I�����gD�y�{��U�U	��+i�f��C��>��\�~�c�fE��5�T�4��pl�7�I*罢�y��5l���wtz���+!Neo����1�l�����[I����o�%M&�L&:�-� �c�B�|C���Ӫ��n��b��}�l���0Z��W ���~�rي�(�m/8h���@`���F���/�`iӁ��亓�8�"Q���aw���&c�ҮRe(fC���6Y�(s�1��M�f���|>Ȏym���9h;HR�:�����OIZd+�E�G��F�H�C�ph������/�����#�]�6\�qp)�o+��F�aQ�iI{v[�r�����˼�8��ĵ�׋�>��N�+���)b�3��3JIl�>������:��� �dֹT�ǫQb���K���᧎H%=�$��cq[b�ҹO$�<���FdCM[�n�	�L=�mK}��i�>&�)I���y�b�9�Ȟ��rR5��Y^�2�`.��"�	y�&�=2�������h����`���f5��C:���.���@��������F�O�R�T��W�xV�j/��24/�o��a�
���kw鏓��r<53J'gE�ۻ�i㛅3����B�#�7��E�7�2A�&cT+�Ń��QG�X}d;HQ/0P�	�J-&',��k�u���T�+9<3���.�	a�'$^�&6G���n?/p�ͨ���]��q��r�ESBŝ�^ԦQ�:�/O�$�
��&�렒��Ȑ��G��o�� ��:�m�+��� �͋� [̶�ԋjRY��O2eś���h����`�A����|6�fp�G̯��B�ޒ�6*o�u@�T �6ѭ�>���ݴL�i?bY�~�������-.�7/�0qJe�ٽ������o�%9��B�y�+���L��Z��)����b �5�IҦB��[#��%�%�R�6��`2�k�[�^HZ�i*>������TXڦE����̞���AA�TN�`K"��x���9;t��Cm��[�t�ϽϦ���]?��Iw)�����;�z&�+�fzCZ���'����H!W�Ǒ��x�2��L��Qw�-��G'\��Q'׸�O�m�a�����fQ�<N�ͭ"�%n�|~:K���-��<�3���.L������N?;�����J��n$jC풌K.��-[#N���ړ6.yJ ���Wh���f�˯�{z=�*�����]�q�zxEU��k�oY�A���P�_l㬁`GD���X�7�8�Y�	-d�Ҧ�Ƌ�)y��P7�)��a�3��U~T��P#�EN�(C�u��{_Ho���u�9(��h��=�@Ë�I���a�k8��@G �$�� �L�[��}kp��3]��AD�����A��2ۡH�lnm�J���]��7ꅱi��Kp���툶\ mz!j1mW���f5��VHU����a~��b��<���j��ٰ��T�%O��@K>���*�d,54�X���n2��*9:�6x��E�u4,����	� d���^
�I݃6Af��,	�S�e}(ɘG�R��Ygs>k�Ϻ	$�u��yˏ�H���W�ZZ��{����ͷ@��n�����;A��M�s �k��ɲ��	�~�H�A�ژ���P�U^k�܎��
6�6IBh��#m�%�ŀ��a�8�h'"���/�L���.��mO�p��C�I���Wn;2E����5[��fi�N'c8��gHj�M���]��fP��C*D�;��4��r>B��9��r����_�]8W���/�֤3TL,��}�? ��(�4R��pc��d�磯����c�Du[	��ՠP�z�%zn�@��z�mJ�`2u�Pd�G C1��1�4�r�vg��e���<��H��[��	}K�0��>��)�]�~��˾�'�C[���P�C�.JO��g�S�AE5���0��a�YB~��! ��]�Hm��;�4�O(k��3֙��ň�_�z�b[��:n�Ek��&�0�5\F\�@�X3`B�~��굺���m{g�Θ�M��I�Hl�1u�[o~���%V��8n�G�!-�[��pe��v����H���O�?������~NO���~��O�I&W��3�hd�]�#"a�Q!�s�]V ���GT��TlW���I}����01ZG�pَ�p�uz�d$�#�YQ��K�k��T�Uï����y^l)����a�6�����5�Nd��^<ݲ��9lPLa��*��b1 P�X�����`)�F�4�.ˆ��7c �*kW��{��7���V'�{t���2�Ė�ܛ޴:������-�˿tYӋ�J؏��D⟃Q���!�)� �&��u���ei�	3KV�P�����E�\eڿnW<5GE�]9h�EU-��+�u�'vXB��د �Lk�ڦyD@y0B���V�U2� ������M��
�N/�-��}P�Q��q$Lb�ɥ��h�8Q��Ɋ��s��aRW\�K��P��MI �b�0���4�����a8&� �"�c,��B)'4)<e+��X����c5�F�a4	�#�IC{�\��A�2;h��U��भZS��KR�j~�IiP@ET��K.W� $˓�w���H6��x���F��#�$�U^.ȧ��z�Pa�����L�]�D8�EU*�n	#\:�<d��K;��Tʴ��?��j��{��Ǫ+j����c7��rØ��:��k��������$3.�[��f0��e����t��˷d��.\r��PC/�Å��:�(��-��&א+�(���}��zIs��l�Z��5�cHY.���$)a�v��#�I��|gw�[��^���P�Y�aT�;�4=�na�������� M��2ְws�Ⱥ��cC�"8L�p��0�M�b+T0;$�Gߝ�/�d�<�����h����zM�|(�bh�ڟ:^,H`���#��09�3��?:�Σ�;&�3�l��G�g���8X�uO��9�V�#�wL���(���U<��-Y���P��ު��җ�)t�`9� ݲ��͵�+;<K�4�%��an�?z-�^`��7I8����� �}`��:j^Lz56�0&�X�a���"D��C�<�bJ��ua��nc�syy��p6��7�V�=8 K�k�%y!"8����f��ge�D(h�������º����ݤ#�$�d-^3���G&���� ��hm!8}G�f�:f1�\��TEy�𳃉Ľ�o�Oʅ�����Eu :�$���z*�֜6Vvh[�ӽ��҆��y�7���Qn���K���9�辭���X�����iKeS�?fp�Q�(��R��n2��o��RF��L~�;>(_�Q�O���ђ���%(*�N�v0��NG k�u�jƬ�w��d��#jSPV��*��Ĭ"`*���{(K`R��tv��W�:({)\(q,�iX&��!t������c�Kf�B�̆Z�D	.!���RW�N�!��c��d��Ms�[o�4�%���}��\���Y� �R�	�ϭ�(�\ˬTt���t�O��'���ۤ�����m3��?J��Vg�ʱrp�q�d��L����E�0�~N8dt}vj�T�Q�Q:8
Q�yJ��Y�Ѵ9�(���_�����|�������v��`�26;�y��%�3�� V�wk�>6p�4�G�\S�3�Y"�SV�G�h1
�M�`K�Eu�J?�U��ҟ�h�Bx�z��\��`�K$q��]�V�\/��Y�1 ��W�Ӣ.�CF�_/Ɛu����6i�KT�g�-�'  ��鲴�;�߻�U���f�6��0��N�44od\>0z�>q6o���zt�D�+|�Ϝ��z+�䧞NE0Ξ~�mc�c�s� �*�&�u�R�a���^�ss��ǜ�qC��I���7���ױ/C����6�f�������{A,�H~�G��4�C�?�IK�K���6�ad)��g6��?q<��)��q��+R�^�0](�`ˋ�O#��t�7Y��#�u�i^H�; ��wc��h����렒h|�F����7P*ns(�1�ɱW��o/Q�{��R�)�,}�f�������?Ga����+�����Z��Z�L���8Y煒	�>\�[E���1�n���Wq��#E�D�WM)�En��������g�H� �l*�b̟?ix8	ڃ�"	}O;k{���Ɣ7���Y�4ӛ#��Q�
���i���ͷ�iR����d*�֑_�벿�e4�����'��ඳ$���U�KAe<�ʍ�Eªe����ih�G��LY�cO�#Xw�RaʟHeUu�Ӟ4t��(�7#V5���b�=���^ZA�Q��Qٶ����I��ˌẐ�դ�h��d��k�Lle�a����,�f��J�H��R?��6å��ԫ����k����HR`Ha���Bަ�E�N�Y�T� )�X�����Ÿ�}=kx��JG�����D0�=5Ǡ(������������Xpm���'r�Zu�E����I���"��f��ǒ>a���(wj�g��֚V�lv�4�0K�Մ���$\���g�oM�>Z~� ���y�\X�s�:r�7gↄ�#�?���|�F�6d^f���^�=1p��z?G��?eၡ|����Wg���kC0��T����(�Xr���.�03��C5N�*����s����b<��(������)S�E��FSm� u��A�#^>��E0����[�����9�[������m�H�NN�$�5#�JI<���	�..(D��N�E�@�u.m�η15[@A٤L����8Jᦩ��ɲ,��I�:�������1/٘�!��mHGR�=�/��f�*���������`��� �����Zf�EV̩�429W�U����Q�9��_�r_y�Fd����mr�+h*���P����������5b�-[� ^�v%'�6©qf�~a�gD���yi%���	O���2��8f�C�o+��� $|�(~�9ۭ,��}eW���HDkmI��D#�%:T=����?㌝5�5�e���
}�����j���[13��m�����8�o9v4.k��2qWCH��~uX�T����D\���^����$�����Oy#7�	�ķ�i�jY6V4f3��ngd���PE������ ٓz���m�\-پ,o*P4�� ����ֱ5�ｳ��9��Y����1[(�9(#C�W6�������=�)�}�`X��W	1��������6�����s�2)m��=��UnMK��p��=�,����)8	�1���J�'\1���Ȉ����B� �׹�5n��2J�?�L���>Q���Ha�P�9�ٜ*��e� �����'\�w��ڽ�3P��Aʁ�k�vv���\�_�v�]/���`�6m��������]d�5�!b0]:�&G����n�+�m�*;;�x:nnJc�sz��۳?#!FڈQ���ʴn�~�����S���Ý�C�r������b�R3�z�7���aQO��<S�^U,n�b0��_�\U��YƂ� $����l?��F/�@���b;�M؛@�y_�o/oT��=s�謸ɀ�'%�H�P����$���8B�J��"n�����>�Kx�u)nGuu҆"�1Av����;�f��	Z�A�s���\�h�{���z�ʐ�Q�h�k�#�J�F�h�����8���E���u�\ߞ�r8$ 	E�m�>�d��l�b�ĵ� ϽEn��jDM1,1��9k,�z�1'��������Q�mG����e�ڿ���)�= �U�O�n��؍ %bG���t����
xǦ��W1պE��u�ݚ�i>�Y�iKѾC	7k���$�2O�0�pX?n��ٓ��VQ�Tvm��S\#,�
����k.���u5�.U@� �A�l����7�0��- ����*�*��y_Q������=��~�4�h�4	[�J�XP����R�/�V�Q;^�ڜ6�h�pI?H1��w2V���o�-r�-�]�LċO�Rj�19���P��*� �!O�<��Ϯ�Q�DW "%L�eb=���O�����F�]�fEe�}��������Ɲp�x.������_�0im
��tQk�+$|�PZỎ�����N�7��%�V�|��;�є2l�f5j/���]כ`���ˈ�5�ڋ�j]��G\��)�W- .c3��~}���p��k�c�N9Q�O�����BP.��N��[��\}�䭓�FI�۞��NU�)���
lTm�@�($G�0�e@��J�$�X�����Est���v+��K��`{FLA"�����u��
8A� ~��s�0��GG����7Pc9Hm��z��*���AM�A�=�B��$I���p0���!;��#�(�%������ZQb�&�9��q׹�:") � �]�fL]��T�i,DB�m}kf�k�ū�0�mk����'��8VO�˯R��C������.ڔ�lS��Q&2���&��bS���7��<
 �d-�t8z�=n��#�c3Ak�h���Z2��e"or�u�+���-Ɣu�oO�%�B����ك�a�]�s�Y����4�`X6��"��ڍ�u�'Db���=u�4�"$�9�ְ��1{,�ծS*��ue��	gfo�tdȇ�9�H70;O�o\I�5-~ɂ|����Rdx��W�I	��ڈ�Bl��m�2�	>�� 1ʏc�{l�od����@b�d�O�e =;�������?�i�A��:�4}o�8Wz��Ȇ�6U�]5������ ��=uH�G��vl`鼨�.��Б7�V�g)�d��=�\�_56�����S�*�3�t�&�t5�狻�S`��WZ[^�j�Q������W���=����V��D��1�
������m��M>&Zq4zv>j�;?B��Z�l��Y��z�!���+��+k�x�-���H6t���F�����}C��@���:З��0o����Jy��y¨:�'�'Ѻ�؇Y��Mz�%���������:����>�~�4h7�XmI혩�N^��,rl���Yȥ��q3S�H������D?�2s��!ò�Vn���9eLˆ� D?���;�!��[a e�pg0�#�	�Ў{o<����Q���<\|�aeY���Y��|A�
7�.F$�[�>$�l������f]���]�5֩r��Z?՟����<V;A���`ˬ���2q���9��8�:�C�46��+���?�j0��9�|��ɼ.��.E��0���ϐ�w��>���ɿGIK[XY�;���'��;�I�<��������6�s4�M���R����륛 ���1^Vۊ�$5(LNWk<�b#���`�2�{�W�[17�$}��kJQJ!��ʔ�A~�w���s��,�R_��6�q%���#���R��� .���[~���u��P��L���m�����/&�])E��;�X�|���.Tg�Rx���ID�HDT�\VΕ�	ԙ��ך�-s��p(�n����{C�*훂ʔ}8Ce��1�P��_���vqt���ܪ�3�޴�-��x��b����n��ǯQY;��Y�"����>���4�/j���?q:题�UP���F��4�y;��gr�O��Uvx_����m�~*D&8�֡����UfTD��ʜ��B8Gu}��B%�02�I����:8`�E��	���.ކ�f8�hițb?���n�D�XM⟬��X�ɞx���@�������%��*��&8yVU���肢�2�Tz�[۶:`"C];i�]W��Zn��&_�߼L�� � FP���9�;�wZ�݂x�V��� A��ښ��?њP��*ٔhc�8�,Ɯ���l�Y��B�	�yōq�ʙW�)&K0�:M�.�7����'#�z$����$��A(�D[A7d�ݟ�ҡwh���^򢙣;1����d�����Г@<�d%l]����l��4� S{���?�x-
���p�w�oJdv���h��&�Fg�L񮨌�K��{fu{ۛ�9�	��J�i9��R�f�"/HXS��9?�ʊY�u���(��[�k~ݵE���1�O#X�+h�5u���w焅_�+}��H�������$f5?Z�
�-Ț`��a��{���aͪg���M��oyU!yfS�x�����׵���HD�v�����J&*���"O�xh�#~�Gr�cV����+�3wp���p��0�]t�X��?51`��\/��YR�}<��������$�k�8���K!���{OoF��ύM*�P��^~�6/���V��Ã3������PnO,賭�b�ޢ��E�r,-�l��,�K�f��ʼ�]|<~��B�l�+K�S96�p/���L�z�L��S�T���v��?o�y�
�����?]Q�%�u�ŝ�J܀U�X�P����? ������l�^˨����/�/��i��eUu��a=
@{:z:���N�(������.E��e.��(��)����GW�/�"����3���i�i�����U�W/u���fGF*}!N��w�應f|�9bX;n
ĥ�l��tq��R��"�^�5㏐�^�ey��|���>Ro�
n(Yc�F����S�"������_IH�(�E�x*u�jNC����^J�Ȼ�?����H�6kM�5d�#t�$���2������9-�U�B��t����»D�E��/�X`A����b�g��d%�G)[g�w��$f-b�A�j���������o���!ԨY��ٜ&��>�@��N�Տ�wzs�	0��V����dq�{�٢���q!\�,���b��i�2�U���x�>����Є6��Z�B�A��3-b��3dc6�_g����z:�8����qY�i�y��qpd;�$�^�oms��rT�x�����K�`�����*l˝գ������A��R�D��c��B��A,���>`MN2q1��8���B�i5Z��9�������_�g7݁��u�2�봵p���9����Ln��TY�yPc;t[v��$j�o�ӻ��?��.�d!���uHa�{K��3(���'�2�z"7����=L(D����E%�����|�g|v�í"��u��ze��6����S�L��??,�����ą�!�f,�pv���L��(�k�1L
M��|#B�>H�+�7JhD�9��f��b��)���S	r���3���>�5K�~ w$����W{���ޫ�����l �_B�̣�Y��q#B�Y�E.w�
:Q��q	�~���ֳ=0}ԱKzLs:��Pȋ�5a�'��!g���Yӥ�����bQ�׬�"�` ��x�ؠ���~LW�|{�j�3 ���k|Z!@��d�.|��)U��3lF|�0�|�M$���$�A��,e�>���O g�M��zh��_�����X����5�?6��9�J,�D6��cpR[=��F
E�Hh���"[)�o��x9�!g[�U��c���	uY�.\�l�k}����!3���=�$G� >�c����/�zlݒ�3L�lXf�Au���nG��@&rgt��&��G���L��T?�Fe���&����V2�	pm��4X�
bУ�Z��3��L���G/W~n�~�'��
4���X�GrNNz����sa���W����xAL��`.V�:���ev�Q=��FF]:[[��K�nE��q�j
9l�����?[!����3���T����t�'��I"77�>��O���H�N-��</��;�ƕ�F���N/)���ZZ�������J����B�+w��;5���X�!:�%�8�C�{�C������i�jGavh?.o�!~o����_UW!�Jq��|�[����o���*�ؽ��K���CŇl&͕<
}E8�_l�a�E�T��<���d����J�2'�mJ��1x�}�OOʴ�N��:nR�|zQ��Δ�?�	�4���_-X�V�����
^�?)�g7�Ѿ{��3�����nf�nG�-C��|���h�A"#�y��9����0p�I�V۟�ҏE�c=����7G=!=�)˖����CY~Xr�D��O�C��Z㜠.^ �o����/�߸��;�d��M���n������y������ִ=Ř�z|���D�����n��D$ce���"�%��d!t�["[i�7���(+)A����&�5�LV�}g��́	4��=����p4��{���,�Hl��|F������~f�ȟ^YT����rei$z��ɥl0X�k����+ΤLx9|�3ܘ�/Y鉗�NQ���/^N��(��9�X��	��Zr[Z��(�Ů���we��]�%K�
��Y���f:�ǉ�NP���bI8�GT����E*Q�H�9̪�N�T<ٵ���.�(7��m�+27���F�:�����g��L:��G}�nJ�}���� m��(�?f܊Y�%Ӣ�g��B��!�'�"|��$ZhmxW�՛�{��N�Z��纉���{��~��?M�V���8jB9{c�ب[a]uY3q8����&]-=G|�y����:�{���3���b�}k�L�ȴ�WЅ�Ȑ�E���u�%�>9=��}4Q
�yxk���aĤ5dnޓm���zF-����Y��,CdL!l���qY�a�}������K_u���Lc"���#�M�X�"���~���3���+�p�����D�pj�49�K�HPmD<� W��O��"�;��4���U�+C���h٤a{<�k���]���}cý;��#��HŐ[٠K����2�,w�Et��1Ҁ�[`�����m@%~�S���YJ�W �ՠ�L�N��������R&q����!8�z�Yy���]��Z)�v���8^Wi
*K��R�\���5}���i�����]Z�}c�un���w!o��r[�<짙��.G�(��8�lѶ�=5Ϭ4��qL���xp����n�	��B��/r���&Ke�O�7ވɍ�_6���W~P3�l$�[��|�t���w��̴�+[!��96]���4�=����i��-����ۋ��4]�b���Z��P�iz8�ӽ��pe�7&r*~�#�@�x>�������D��"��Z(1;�D&��@?�sn�x�����u�D��e~SA\ǯUfhKdnG� ���z	Lf8�5��C�-=B����;<kG5��Dzb�T�X�-��5>��ƨ���o��J΍��~�+�����K��ĎCjg1��9���<�T��qY���;��ƾ�&}/��z� �&�d!������Ol���.
F�d��pZ����3��"�~���޽�l&��M�6Ӡ�q��˪����!�'&�+U!\a���kDHp����\��(.��9"��m���~��#a����g:xJ:��K��a��꼐�d����~ֿ�����Pǩ�f�I�_D�z���\�����;����"tP�> ��I4�h���05_+���b�mjC@:��'�h,�J��JT�-zԩ��.P$��%y��̫n�����?|^�>��ٞ'�����M��(�nՂ�F��Jۯ�8�+U��]����eA�����5m����*�`�x]��n.x��*h�P;��I�H��A�`���$W��/W��)��{�T|��G :s�j���F���#�I�_�m����م75��k��i}[��=��=_,��Z~����ŏW�.m�"a4�!�T���w��=Y71�ƫ8WYD���o��e�!�M:h"��1���2e#>�t���niY�*4�E��M9@�k�`�B5i���Kn=������u�3��}I8D|m���)7� �(P�=i�΂� �,B���-�x@��֯b_6��յ>�:9���KBo� ��'=�b̦<�xc���7�vx&�/�����ۭ-�p�E�.�Z��I@$eX�<q[!���d(��[�1f��c�J/�H�b���Ή�y05�(���=�z����fA)���ʝfc粀@>-|�7���`y�v�r_:�O�[�Kǫ�,ԷX_�H9?�g��?���ڊa�U�kLIR�W���&��	;�sv�LBa��$�nȐ&����	DS�� �g�;�eч͆���'��&O�dӏGf����>����_9>�EMV�_�L��R��ĮΟ�6Z4�(Z�ο �2��&߾�:I��US%�_��@r'�b\��	T���{�I�.����o ς4�NO���5w���Ƹ�+�/�K�;�ɀ�G���4x�z�~���j���qb�����������<?��Ca��ղg2ϰ�oj�I��2��A|�J��#�N�x�@���5kwW�Z�#8/p���zR��d�����n���wGzK��x�Q���D��u
��*��4���tWMh�ȕW����4�`d��~w�$��F��dY�b������ݳ�a3Ӣ�b�p��J�o�Ҽ\�0,\<[����R'_�N�8˺�N��M%����if�WXx�PL��c�� ��>Q��o�|� �i��ĥX~�^�
(�O�p��A;&��B/�Y�tz'~�y�2@Զ�0k��K�;���JA�{�*ĵo�\�']zR�1�J�Q��FTgI�TO��U���vm�,���Vc�eI$FѐT���-A��r���B/����U앵Ěc�D��?�WI;�0�W�V7;�F�5�;PM��d
��AQZ�n�>2D2Tn��#�����k4Ӥ�QH�b&��y�/8��!���'$P�H��et�[axV9�Jx��K�__�� �m�yBHN�lۆ�m�LN!a��Q���Û;e�v���>��nc�1C��I��4�L�c(蔞$*�q�����*��Y%�<�{=���I+{:}O��!	9s��_��I�%D������3i\u�hxMm\+#���[�k��.��hG������-���+���.}2M,�cx<�r���J��٢_���hqHH;����ʒ��*���U�S9�n)&v���K\��
�v�K�ʢ��/EV] �*t�P
M��`�7+��%HQA�j8ָ̞14z�ׄ�w�ٱ���v�y2�=�����Aa̚T��-���|ーCf�h*y�M��#���;`�����@ˈ+z&")�
G�;˚����y!��KԂ�¢J�%�(�ӦLu�3xE�}4G(H�rHH�c����qN�:�b�u��aͮ��{V�gL��ȦI�Y�U��N�l̖��YL,�o�$�j�2 W���v3��c�:��F�r�ݭn�D/�����Zc�en3�/��!��/��O8#F	G���*f�wJOs�|�H�naE	� Q����V&3�[PIi��j~X�pd� �N v�ᙶY$ڜ�Y���@޽	z���ے��E�,�뎁���&��$�16b���TVxt؂y���,ě.rF�ǿ�{ � ����Ň�~݄Q���c�=�ˤH.ϖ-9��%��ꊡ�\��eP
N螉'K�/lL2��P��g�}O�<��o>ș��BɘMQ_�7�':��H�P�K�����>(�Ͷ����ک[X8���VD�ll9չ����W�p[m]��~�
��R��d�F`c���r�jLg�����ƶ�%Y~�Bv��p�a\�:��DqS��-�ށ���p֕C/��4��w�{`67���������}I��n��2Uw�Ǚ$q9�9���<�w]���7�G�d>h�)~FQ���wR 	Xb�L
���
�6wB4	0P��6�x�	�D�+�6V���v�VI(���U�QlRA�ڝy���h,���+��;�M���Le�q�rB���D�Ô�ǹ�y(7W��z�R��DC@F�kF�i������<t�b[���&���y��ݤEj�*�HC�,t<�%/�����:��+�p�_��H�G8�����PZ�%$Q`Ū�&b���x�M�蹖��f��t�G%bq�r�A�)8��:��8#X+-/��>׼�@���=�X�����>�:�:]���i�����ptpư���H�5���;��h��]U���|n�%)�}��m��ť0�k�Q��ؗGI�	��l>���1s�ڃP�
(@yC�ޞ.�t�N�	s�T`)Q�?��D�*��N *9��]�{1�Ϋ�u9�$�-� B���*x�Ȏ	}��� D(�����
Jd[fH'r�B��[����:�����\k!H�R��u(�?��SOI~ ��?�`�Q�\8�H��z��2%*���{
��ej�7XȺ���Tb��?$ap~�����F�ĝ�����r#�~A�6��|�{Mά����G_�����V����l��Ȟ��|2(�?�#�tt�
�g3�4��oҡ� 7�n����::$�*>������>��y1p�P�+��GP��n��c�}����r�mX��yٞH��`T�Q* )���	�߃�D��,)�]����C�H�c	��x�ۂCWR����V�\D�2�ی~8�'fvY�9������\��O�;�"�'��Ȇ&q���]�l��%O7|&���ͪ��Xw�#a,r��e3�������ڲ����<>���6�촶^�'>�]�(��$�K��|@���mɃ~�9�ɠ�㯜?5�W�Cl�\�%��Ǆ��l������@J�! *9k�c/�0s�+�8�?{�&�cGw".M�[u3C煱�]T�WF:@93\VC!Z	\4�@i�V^��a��|�������F�0/�D����1o�����_G�	�s�����(��~,���Q�{�+�m��_6���~-�G�&��V�����T����q���T���<i�b�U��pa�8�����H��bm�����`Jr�3Ogs)#���&�e��s��ˏe)b�M�zX��Cl��d��Ғ3���������ί�O~�j�!CŴ���6U�F�� �g��Y��MO�7_�i��=�v���%GR��h��Q���v��+��*��I�{m�w�z��t��7�c��z�Mm��͕�G�QN�n��NMT�+�>��1�HQ�0�`���>K�"{A>�l����&�[C�י��� �n��1)�3���,\R����B����%�0���#����#�{��D���L�Ig{�����b�l�PKA*�W����D�����i�R���z�X6�n
�-$��T��o��f��ށ_��[���Qʘ�����MX��e��wsb���|F���vՕYb��Wg���?4�!g�"�Gܶ=��ռ�����\,=�����מ�Vu7��S���X-)0d�t\�1𺾲��Ƥ��CPn|/�Z��*4�.H0�E�-��qw���	����d�r���J.oO�0���^\4d��XZ������!�z$���~.����Z-���Vﻩ��.��}R��Lm�[ـ-���(��z�[kJ
rg����}Wv��KI �b�sJ[�I�@��Y��K�>���k����@��nH^$U,�]�판N��З�-��-,���)���}65�M�
� n�=�S4�=����
��6xז�-42&�~�Fz'hj{�%�jV�C^>���M�U:�ο��)�Ɂ,2è�֯N��E������:ҳ�a_�Y+S�6�-�䨥-�Fg:;a�g��>/=�����P$?��T��T���b��pt�^f@	9hya��C�u�%T ���K(y�﯇T|f���|޵���>�9�X`Ъ;�Wj(}��Q��D%������2K�I?�[	�r�mC���k�N�NLc��n&��,���KY/�Oߓ��%�܀����j�57�t�2bߞ���Sx�}D��݆&���ٺ�R��a��`ӊK�^��L�T'A�i�@)�뀍���)�m �Ce/9~���}y�Wu(�q��K�tZr]@<`Ӓ���s.�l��P�1��E!S�d����yYćtIQH��w�����(���!t8��8������<{�;X�)����8O�#�r<k�?2e�C��j��_�%��6���<��ٸp�Kt�2��dˠ��fZ�x��� �������K|o�\�ڭʤB���@�t��SAɍ�̖������.���q�3�h��協aX�Ȉ�A��HmmD$8d�n`L=a�FH�=B���U�A8���ǜ�I�*�[��#?.����s�S�y�kx��!%�	.�~	���טO�V�`v�,=j���\�`�,�V��'��� �ӳ����|G͂Ϧ��zFR�6�hIICt�7|���2&�����qu ^tP 5��E��d��?ܾ\��������C����.��Q����``g7[��e�������.[қޅ/�N�`��AL��F�4�4yT����ҥ}�����p�;��A�3��TQծ"E9)��I����t��:�%t���!HRjB3K��O٠�����u��%���oGmc(�x�,1�o�}E�`��)TmW˫ M�k�;1uYߒ;�8�/֚��D��$[i�~��Ŋ��γ�6J޾��o��(�R����p'��7��uIiX��P[B2��E��H���nl���j�&�ν���,��RG�W�s�7,WV��<6]���
@&�F����i7&㑯���olx�'B"MB25~��{��"��~m��n�z��Sm��Y�Tx��l�M�#D��ɱ�|H���2R��)�cj��`-P��5�b!B��I(ΙA�;>ބ���rh *��j��"����6kJ�q�qD��'jT�y]�*�C|�r�}�����/���I}C�s:F�F���	��L�͉8rT*����U[0�<{]����+؄�Q�_��Z~]���FժCכ�G{!i�wy{��E���x��U���}A�����t���@l6������u
S<������^ģ��X<�dV�RKd$V��&��aMO��VH�7��z2�T�>܏��j����f�7�ݜ������@ ��<ѝ�����/�UN?����g�8������n�s�j�B�B8�h�[/ȅW��'{@5�q�cr�$�3���B:h��>
#68ױ����(i8���b�ۥ����-�y�m���5�s+=�MٸGZ�wW�������;��,�_�l����?D�7�a0s;y"�V,B`?
J-iR�����x*),'�M8����MA+c5>�� �&O0��R�c-��wB^zZTWs'�5Zy���Y/���Ds&CT��8�}G����lZ�_����	�ȼ�FE Fq�`�8R�/v�~Y�I{�m�a�X�E?
)V�6jW�������cÓ�"�Fhݰ9��G>O�:���, ��o��K�l�:c<S������6���rYhԵ�N��'h��b�����;1��F��betb�R��_ё=�ιY�_i��o� 6�%�&��Y̆v|��wr;�A���Z��3WN��B3`78+���p|���@F��f�����[���*���R���j�|&%��3���ْ�'e�E�9�it,�nC# R-��U"�~�p_���糛���#�Yq����1\�������sH�L���h!�@K�/,.w&;N���I�']ޑ��}�cHbt�x� ���{#tPh����q��Ld�X��*��9�ҁh[B�o܆��r��z���R��3�Wq��M��{<7���<�y%a	��f{DZz�у�/���M��"�I�+��sbJ��B`c����۶f�ȭ�v�gsX{\�,4D���(������E�����<ܪ�8�⮟@/��R7��Fh0�����JmO�GB���$��Y���J*7~���},�x7>D��=�ak�=֥v�aekt���8Q ! S�vJ��F蹸��vYCpey��uB���S�x˛����L�?ũ���
6�� ��~���&��Z3/�g'�MG+ތ�y[�FO$�GH���]"N Q��F��v�D��
q��j8+�8��T��pv�	�.�l��&��JVj��As��a�� ��{^�!,6}~�@뿫.>Kq8M���
�	У�rV�v���T�RI)���Ϳ)�4"��P2�؄�?'e��T�A�y��n�Ǡ6�V��Z�n�
�����~��x'Z��p9��Y�(��*k�$�ۅ�>e-$�%���\j�zI�f-��^���l�4H�C��]T|w�\N�i��j��uN���8�\�1��JrsN3���t�a��^�_>����_<�� Ɗ|[�Zf���G���ZI�o�
yH�>s�C%W���u�W�Z�Թ��[�b!�����g5k7a�$-��@\���{oݼ�ȡ�w��n��C��"�*�I0V��Hħ�pG 0�罎��k0l;�O�9�˦�HcW��/�S0�f��&������]�L���h�c�|����J�f>aM�U�t��
wJI�]H�(��ɸ�2�߱�E��9��x�P ��=��MuT�������Us��6���c�A���Xr�@��4�S�=���{��0��ݝ���� �ny�F�lt��y'���a�5������US��M|�4/-�����ʦ��՗��Y~�b��D;�1��}i�6���u�!r�����0�I��.N�RH`��'�
�g��r^o�!�N#�OUuS�m�R[�ܑ�{C�W���g�4�0ȯMC�
S�nӧ��O�0�;�C�H[�Zx	z�|���0��'}>�⁵�Q���.$���58�#�z�zFF�S�^
	R���uu�Ճ����L���|��"h��^�ץd�۵Z&��/J�r�B}}�k`�d*.?R��S	��rJN襤�)D��&�8����	�,����v�A=����A����PeiM#��>^������hia����9� ���U�'��@ak��Ҁ�J�n�o��|?޳::��Vʡ�SH�0b�	�74\ڵu��0�:�)�{�#'��8T�_��7��4J�Uz5�ѭ�����sz7��x�4�ô%�Dٞ|:��"�9���"&���'��ԣ�|�S�X?���q�g�<�f
�N��7�/o�`U�2*9����S��j��y�®-�R��F@��gJ��{T�Ot����؞�cr�?+'����{G�Wi\K�s��_�"x{{���ӄ��`��L�|zE�K��6��ʅʕt^k�\��#3�{z�[d�t�"��u�	W�V���ΣD�eP��2��p9Ž�`\����t��>0Y� �*�����C�|Y�/��8t��d^�i����ņkWϗ������ �Z�ֻ,o�g/�;�X�����
W��]����*�a�Ͻ��`�mN��g�R���'TZ��]=M�3�}�eeR�SԵ#'�gv����qkd�a��N\��!��������s���5�[�X6����X���.p������%�&�M'�>��nO���ċ���`�`yP����+0@�q�� �A�&�V�>(<�8�L�EFh�yuy���h�jЎ�/��I���9BRz?��E�o��|]�dH��8�=��^�7�9��?�p��=a��Ӎ�j��������e�r��3�z
ꓞ��p�<�)��o�#���!_nd��$�3���eJR�Iy`]���B�/D��L���.�i��>qxth��W��l}�=��m�%�΄�b|���;A�#f�nT:V�PA<!T����Ԝ�����kE\ą���j�,�2�<��_��.���-��;L-5cQ������m�}.DBQ������I��,��-�ӄt6�1���0�EV,U����h(l[:������	��x+Nl�a�����ʔ��8mJ��_��S���T2߀����'*#(����|9�.�̶l��0&����JY�YWK����D�/oKsR���%R}�?���7~��4���E�l@����|��)��:vD�&8�a�*�WQJ�'��k����x~��,�X"�}�j�Y`�)Ӝh&��̨c� �Hb�,Rk�u�z����s?k K�O)�ju��\�M��IN�E��%��KA�b8�P��4?��(���j,+�0^r�┅�����e5��~ś�l�)���8�>�c��gA��Q�~�s;���x�@L�}i��@�tH*�!"��)���X�w�!5��>b���k��2xj���m�]T��3�N����#fs{�Í�B]�D�TK=���Z�u��N�¸�gK(a�NBV�$z :�;�8.%���ddX|B�1�a�,�O9Pe����L����<H�a��l�_�<�H���^�(eh�Q�;�h�����iV�W��g��]���PEJ�pXsj��J(��@�x �f��5C���]ee3rZ2"�c"�7�vE�}�	|�ƹIcV�`���>|U�Ҁm��M�}Ӆ��ٽn�@�ȳZ�bhR��9��i��j����C�������%ݻ���{_���S����M�g21?5�&3W��9����;��]mw����)���v=ٓ���]dIK���^�jo�ԞH�Nn�Z�2��Bg�N��YMv���_"|+����)F.��_��-Fؐ�"P�-`75[��\7�{D���I�>7w���u�i�je�"O�.�KwH3��S�3�ˑ���n��N�
�'�`Ɉ4�rPvo�,�裱����n�>�>L�;����s2�I��.�lS�܈n*�'0��L!���:蹝���RSrcQ�O���xW*s�����YM9n�`vt�s���-6�C��I3:�3���_?%	p*�Ȟ���zI���� |һDl�<1�/�2AO+XL�^4a�2�0]�z�\{~�Ԏ1�;���j�S��e|<\:��'�PR��7��NG�ܘ<�F�"J?<�v��ㆂR}e��
���y���}���z
ӯ�%B-��"���Wsvwr�d�S���z&�+����lk�{�C:�w�N�$���!�t����L�JZ��?���b��l�P��!ʦ.����'+hE�V1�%�3�W)�	5����5
AI� rB̷ �8<�%�`��c��Y���)O�	D�g|�6v��K)�Y;�	F��VJ)Ҋ��m�6�<{܁a��J~xª�_s]�}�W/�u��lmfxw.�*��������_��w(E�p�
�Ÿ������km��~֍���[>ɦ��J�4`=7��&I�#<��H��1�Q�$�w$�;��+<��D(�Ic���`&�'��N��P4T,R�~�Z�g^�&Jsk�0QO�Y-�:��;��_8LŸq9��%�'լ���Xg�a����'�JR����7�םF���{J���
��kҭ1{Wz �81gc�љ{���Qɲx�qy�PI�F�K���"����m�:��D��^�]�u�1����q,&��B�Q���}	��r�R���
,O���	=/:���X4�'����[�E�����8�c}�Bfn)|}�c��Hkr-������; rWɜ*լRq�y�,�s�r��Ug��Ļ1E�DD��UF�Vk,�3R�Pi�pa$)DUw��v�?�2����[�G��}n�s8WB����H� �Mt$?�e���t�Đ���>B���Rӓ���`��o��� �����{I�)�#��FwHZ'�h:���;�I��P��J��B�^2��YHΑ���t�*��3��J��߱$a'�-��֠��P�Z�Zo�"��,��E��qow���{�.��U?�G����PI�~�����	H��&\��m�C~p�0F���n�'�N
{��VK�Y]���H�0����f��xWca֔�v�]~(Y����b�ܻ��[q�
�F~V�M冚��F�q�AɹQ�¯L�D�����<;�@����o�԰Q��UQ�8q�xDk0��D]M��|���ڵy��y	�4��x
ԅ��m���B�:3���q23��yl�ϊ&(����E�2��'�f�*�(��5�U�,�X1}R�]���Ո(�s��p����� ����!1��=4�w�O
��CagL��|(����9��WX�o�}!�T�C��UE]����7 c��K5g�� �l�=���E�ɰ�m�ϡFx����|:�_������*
��{�4ci�[�Y
.Ƽ��{K��1�_�
�X<&3�� �3�� ]Vzbm"��5�څͨ?<Naz�Qt����a^D�s��g��#�<We]����t��&zըV*��T�K���� �m{;���8)]4EA+�@�䬅�-h��|)O��H���g� T��K�έ�I���N���b�ξE�M$�>8"^ ߀���öQ�-����m���7c�Z{�G�#�ݒJe��az���<��E��xu��rsdUp���!u�-f�H�>L����#�*�*������2z�&�)g}�P��f������c�i����6L�52�o��������<�S���5�y9km<���_|�f��T��̚x8|,���Be�GJz�}	W��g���L�!`�4�6�z�׃�Yf��^'ϫ��Nh!�A�G���.O�0����jE�ږ�)��VWￓ�Lؐ����>hq��x}�u/Y|&��хyu�J�v�,~�����!L���n�Z���o4��O)Fhav�?�%����B�La�9��ާ]�q���� }�~�6m�8O�׳L�{������CC�S��q�>
+�������P:A|:�7�"����P6@6t��kH��D��զ2�};$�R�x�����jJ�?�ƍ�h�{V�?W�M�ج�,��츂#���
���|���fM{ay�{�����/� !�AR�F�=��q���x[���n�4��eU��G� �VM�t˗�p~����5'�b�%� ��\����G�ٷi�i����������G���o{��T{3e���W.��6��Kd1�gQ�)o�,i^C@@���:
�plF/�N4���g�y�j�XE����6��zgxX�j�J8X0��`�b*�0-k<���O"¡�ը��߾d��;��,��px�1�R�Z.��>�k2�\�b����E�`�6�*��T)4߂�~�-��U}[IЧ��ZE�K��^�I��2QM�l�Ԣ��
���r9t.���5�T��'�F����q�^���B�
i4[%�c��Mߦm7ru���R�~�ԋa��r�h�A�1"��Q�P,e2���0��i�T����m�&8˲��^��o��3ʭ�p�d��U��m�-�:k�V*v�-��Lm@�2���);�x	��B�1���b���˔�"%��[�Qp_���9�̉��{+{`T1����m�W�Ypvʑ:��(?�kf��)��!�*���p\6.���-K��@*��ϖ����~�	��;�M�ĸ��H�z����D��
ti�q|k���wc1�s�,;����F��^�I���d�ݨ��}]X��VW��<���見!��h�sV�
�?Cr"H�ok����R�r��K����Ox������Fuv]����< 5'CU~L�+=�������u"�2��*ݬ]��>|ʭ!!SX�tM�i}�:�����3ķ �J���Y������*,��x������K����0��O�3���k�iN�$��)M)D��ѥ��c�x:�=��ȥ�9;G%7� ���[�}XH����PG	߶�9���q@�:x}�ż;��	�ԢNy��7����l���?��5R�y`ʠV!�i�{#M�̀�v��T�F�Y��7@�ozs-PV��6��ԝɳc]c⚹�U�.��y�풻�� �~̀9��4ٶuɂ(��Co2�{�qn̖۟�Q1�+ 8ޤ�i@����9!)�N�܃O�v�&y�8N�