��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0���C	�i��E��$��Ȯ�_�� o�0},��e�K�	��D�(��.�ô��by�I/>ɦ����j��������:U�a�Pk�Ѽ�gsm�כ�s���pV��>��$%��"zr���TJ1�Y��tr��@:�>�8$������B؜�7�6"〃����%��A<�o�f�����X�'�����7��!��bM!�i��=دk�b"���U4�����i�0��ٓX�}=&9���1��&';�p^��E!:�6�E�ɆX�Hå	Տ���=��Gc���ˊ?+%øCY3�B�{��'h����v����rG��1��y�/��b�~�-�o�����G:q�WEl�Q;$B�LEUaG7����ş���h�\@g(��#}tЕ�D�:�Ϊ��3�57Ӓ�Y'�����Ӻ��V�o+ʧ_QG����'Tp/=�"ΠUJ����se�W �v;���Iy�E���L�	�(e[��FaV�w�"�vs�<P:�Ҽ���LO�L��A$�!<L��FjY��d<sI��Lh���ն�y}��B���WǍY���)ʿJK�X���2U7@��a���8����-غu�]�g��~���Rɘ�<��/��[Ѝ���Շ�f�u�k��4��	����G`*e4��{�������[�|YY�/�\���h��VD�a���
�-~2�,��5�r�VЦt:;N���@%�Ӣ A���Dḹ��d�ʲ�@Dn��Ǔ?:߾���8�� =����d������A$�E0�R��_���5��n�<aܮ�?w�_K��e�����j�Dy$ݎF�����b"�5f8^���0>�1y� �����S�5@�v
B3�!���<%r��f�#��$@K�2|="b�9���)�=Fkep;6dˢ�ƃ́4��^:-��b /�'o���œ٧k�	����q[j�v�F�ksJ�[��F��k[�^$�C|���a�k���x��֬��2�[�7J���>'c�����`��챌����M80�u��"7��FuX�"a�sM<"֞��F)�$�Vێ���ws�UA�G��_�뢡�a+���j/����w+���f���q���j������Gs^/�ɭ����&k�6H1_�y�R��be�&J�o�����*��jz��\+<�5�7�Ȭ�YBR^w~�rz����A�.��%�d��_}D��~K�J��Y7P��^���y!!��O%�%l���;��d`m��K�MK5��)��c)u�;P{F�!hz���c2pg�g�� ���d�h�����jդ��gF��
:��'�*�:�)��2h�T��q�wӀr	���}�@�f�r��{K�ϛ���v�q9"�eM���V_&��z�ɗ㓓<?g�5֝���/��D����Z6�!�ӿpU=W�E�=����%�b�DG�������|vi0_��u��lU*���5h�ҹC�O�e�V� �C޿�|�}O��6 �l��֗�"�쨧n�3�+��BG���Ż�cS�#�<����%�բ ��'4���ߢ]���� +��x��Æ� ������c���z?|��ɞ��9�K�W>�j>�q&��:�j��Px���
|��H��l�ځ(���K(az6T�����t|f8���.������۪g���F��2"G$t4#���b�@�l��k�@O3� �=TV"R�i���*�xs֙"�W�~��=�y:� �����<���JqL
�k��;�!r X#��쩉3��L�w�|aD�n����(��S�>;!�6��H*�Q�x�^�2Um5���a��z����a��]#a�L�@���A�c�j9"4s�2�@JQt�/��3�c����}��<��^F��1��Z(�d��L�G��RF)זּ�􄃲���d�7ZPZ�F�U��IG����W���3����ԭ�����[���d��ւ�Z�? ���bm\�ͰKv����Sf�U�L�~��^�0ve6Zl���W&��p����O��}��߾�
�Yr=t���k���~�}}O��@&V`�������� �Z>iVFZ|OGT\Ue�p�����3�����߿���r1-�g��&NDЕ� |��y��$kf}�?�*W>Ͱ7�+! 8��
qǒ�k�S���� $qǟ���V��	 R4|+��Np�%���Hh����ߎW�?�he�g:�����fo��O�al��Y��;i�Wۣ�?2*��
Ir�պ�7j8�}5����-����B,��q0*\R�m|�xD3�ޝ��ƒ��A�	��7ߦ���-Pq;�2twҿuq�V��4���LB�NK��Lc�q�L�1b�v`�� �� 0��� �o��IMz���|kY~�4{�u��/أJ�.��sW�m�8!z�%lmV�e1�R�h��V^�8�>  I�����>���-������r�FV��/�s�0�?*pr��H�8�k�cC���J�R).���k�n��NB�ɠ����)ƾMM����%����S�7Nr0�@��>&d��I�S�U������jii��	!T?�T�İ��	�n0�mAK��^���7(����D;�B:���2��C�62�򺍏��+�����s�?-r�̬���7�G�!|�^����3���u|M�v�M6��~�]\�O:������E2ǰ��)1���
��U��6:@�����4B�Ԭ-�������,Em�e�"���c���x0,��/ʽ�p$�p���0<[�E��kt{��z�c+y�K��ǔ�0�Z�8��T�!���\��aR����-�q�1P��p��Ć�
	�Z�&`;i�*�E�as ���Z^��t�4�z����ٙC�}��m/czPj��D����Z�gHF��)�֙_/��,�s.����T׾���2<��*�\��5�4������{�eE�j-�n����-k�b� �I��D����۽����i��clὮ�3,P^0X�S��������p;p��N�����P��Ǉ�6N���;�,�1��J �u���-2��x%���S�FN>+W侮�G�:����T�y��A��_�*V�����)���v�Bk�e�/װ`�YZ��G|TH�Ͻ��=#U7�6%�����,��@U��!�[Pƙ�'w��I9�ݗ��:G���ތ�C�ed�L3K�Ɲ-�7tt�߮@fŏ<����j���!�6/�g
���݃�Ck#����*�N`���&.��ɾ�Z?�Ba�x���$��Pį�t*x�`v����!�����gcG�n��� =h��,i����(Tm5j���`$j�uN�grmQUX>Ͱv��m"��W'/q�v)�0��sG�G����&Tm�/ ��	n
.b�~$L7^�|�\s7m�������lz���M|�g��ûcK��9%�򢖂�S�j�4P�#���gFe�f�ȲD��@�f���}7Q>n�	3�o�o"CƔ�(���ݍ����
ϙy�K�6�U}5e�)��ݮU">��O����TT���z`��S��3_�>���{�~�t&c&S�f�jFe��(�=��5�`BkA�
���o�h�l"K�u�3E/��	��A���(
�N﯋:�̛�I��,��Y2��'�?-<�)�z�i�i�Д ���S��6�Mi�s�~��w�z`���N�nj.���:~D��0-�W'�p ��[�8`�	k��*Vv�|ܑ�x�l�2d?�{��O(G�R�4&�x�ߝ�7���	�����m�{S�_�J [�D�
��Cy�|�o�a���8G�U��>�$©tm�Q��5�~�gq�W��Q:���:�D�)ޡg��T�X��9���"��q���ֵ�Nƫ����2��S�$��X��s��W�����V"������vٿ=��A�M&%���%5����_"��eQ�9x�l[1II���n��1���P���S{�E�Lp�X��@n�+6�%�~V���|B�O�����#CU�h����<�2-z� �d����d��'#~I35����~b�->J��ݞ_�x'2�{hZ�re&��-L�\�iݔ�t04����;e�+�D\�z`X�.����>�F�����a�K��]����9�r��{�7t��NgB;L��h�پbtZ)���4���
�#��-�d:V�NXH^�̜U�!k5n�:����b2�2
�C�3�x[dr�N��U��Q��IkW�H r��c�F4����$��\���<f�j{R��L;�yl�`��#h�ڥD��x��k�.Is�1o .�It-q{��C����>5ny3 	�K�f�gf�{cӑ���W�e���w���X@#�"�T�Ak�T�N���)�S�n���߇S+u�=,5�����C����qrWܬ��dz���`��o��v?0��MzVq��1�u�ۖ��)ܬ ��z���p0�WT�ț��oӖG��J�?!H��A��?"]�MxL�����^4��b���������]�7���G0�J.��\�k�I7D�''�N�3��CH�P?��򒆤�ڍ/��֓�[U��$���mY'��KW��`�(i-e�a��/���j-Ka�΄>�ѭi���F�~�Ю"S�_��`��J��ƭ����=�b�X�PF�+�U�ɍ5��0Vfհ�2r�*�1Y+��nD�9s��5��1���pt���
+h�������Y�b&���
�Ϭ�<�wF�}�1�Q�(k*��Q'��&?+G��GW�OdTe^*u��U�d��gV;�13�}c{��$)�佉J��BZ	6����2�'a�:p�����GZ�;~�ۇ�� -҂����=\�J]z �ig8���+��ҟ�a")�eT�����U_P�Wu�]g���ͭ��W�Zߓ���~U�B��!N������̕\zh'��6ɕ+����e���~��x�o�Mہ5>hg��Sh�l`V }|���MVA��꾥��R�L?b����=p䇠�C.qU��Y���'�ɤ@&�;��.��᪤����|ٙ �BD�Ŧd�+�o���:���^ꜳ��{��<p�	���iF	^���;��Hz�S�7k�<�ոl4�����iNXR~�"�u� ����Y�ʯiXKtL�������T�Q��\HP)��Piij$@�%�Z8����%�q�%0�T��I7b`�@�y��ȩ�c��P��N.S-|�����CSbx!>]��a��zCت�5�	�4i�	�%W�&1b�ƃ�bµ��}Y�{Z|<�k�e���(�7�t���e��r��`��ih���'SM�،Ѝ]1Kȝ����`v�*��9�U�����[�'���g;�� '	�>��H[�}��s"��xq�j���Tzԛ�6�c�KߡL��>��çA�TYQ�Ԅc�v��Na���y�+�N&�b
�_`�m/�^&��h����FZ��Yv�%4RN��1�v>�W�� 4��PW�}.s��w����0Rha��uY�j=��]R2NpQ�-Ә���Ɇ��59ֹ�Uc��_?�"����8/��Y��7��s��*,<7�2�%�,N��P,�:(����X��pp�����"��Syh����'N�q��X�p/����15����9Uf�"6����s�u�MJ�WM:o/� �Ǭ�X"\X��i�W����!�d��`8+�P��x�ڠ�L�MZ���Ѭ|�������vp�ȊzY�Y#~�Fb����4�)(�7�^C9�����+��N���-	o���Tu�Z��kj����{��� )�c_c��[W,�'H,5�o�r�"�`�q��.h�(d�6hI/�N�� +�6ܔ���?�����߬�����*w������ր_1��,����,D4��Ս�J����:�İ�wX���P���.�L�{�,�1��*�˼���!�}iW�����T�0$��i2S�?O�$+(,� ��lF[���)ƨ0s9�0��U�=&X<�P�E���{mK0�O�TzR��ם��%���v�uP�V��{����Pʠ�����ݷ���`��E���?�[l� &k����X`n�(���`"]|�;e�*�lnAM`�E�
��H]�:��Mގ�=�iM��%OuK��
Ea[�wˌ����V0�dڼ��̚�-S@��^�����N�!�s��u��҇������ $�.�HJ�`?wp`}���1J��R
&�dob���md.��@�R.5f���N7�(Ϩ
���D|���I�6��_G���(��J��qQ��)Db�3�8p�$|��eL��l#�H2�v�~��5>�v�{'F����fS�S���G~�J���	E����$��bڦgQG �/o������n(�݊��B\90Qr@�Q������0��v0��e���Nf�>[V.`�h��;̻}���<twq14���EE�B0��*����5@ckiJ���yE��EN�5S���sl�Xυ{C��ԟ(ƕE�ǻ�)y;~������r)9c頼�%�qc��P�1Б�x���D���^�Z�,���=�C��殕�7>Ѵ��2�v>�V�������F�$ȒS�F>Hf\��o��},q�()��� .l;K�������5�)����v'�%�0�}�t�=k^�l���.�d�ȳ?��λ�Qh����^y��; �=ø��?�>��#���r���?upD�U��u��ToVR����Z���8�{�j�!<G΍6#�'ͽɛ_ä��K������p��~l��"q�{o-}������e�%��4*&������G�ROO���6���L����H��ͽV��R�Y�Ǫ�����U�iS�yj���0qN�c�@7f�l;��)ʩ��/R�&��]�o��PbHTب:���tq��vn�`{tjl�˛���U���1�q��2l���*����	���ϰǤ���9J�6�m����B�
S/�I��k�2[��8*��j��:����$lp��ǟ���=Sseq��=�wP�39`���sͅ3�Z�� �H�FtN�|�'�i���W�g���P�/Py�_�U]����k������Ҵ�C�$��Ҫ�{�,�犨M�=�',�)��r_���#�ˡ5)��������8Hɖ	���h��
0���qj�\���U��!+����0b@��%�ܠt<�5�.�OE �|B���S�4�( 뚖P)����l-2�j��@�`P�]�Z7��C^�2w���������VfD�\0Lģ����s^h�}�D=�/��ku��(�^��_$�Y�~��E���!�������d�}�\�\D�5}<�����?^!�o��Y̳���1��¸#Du��4�|�F�ަ��i���2[�Ǳ���Z����V��E���v�X#m�{��*�/��xY'�9�p��P�.�}�p��{��޷�����>A�u3���w�f�4H�TꞖ��o4C��������۶Ȉ�c���<l<GV���>����b�����x�ٞf�D<^�z�����i�nHf��9a��,`5v�ǀ� 8�A��*����NS����R��<.u̢�d�8F�v9���&
ti���^E�xPg�F��� �@��� =Q�F�w���~ȋ%ܰ��I���m?OF�혝���K@TW{���p-��p3D`�Y�F���a���g,���ݟ��w�1EIrt̆�=[^'����x|� &��8u�L zs�7��u&��h�lv<�5��_>�D�qQI �9Q�zꚰN�+H�qݕ�ԁ	
]���C1i���V��Y+zBp]8��2�&'K|�bp��������ڀ�C��_�cR8�����NU��w�Yv>T	m�	�Zcׂ�L3Z9j����~�*�3X;Ґ����x]:����l�8�fn[�M�e�\ȶ���K��G6���ͼ����h�R����&=i��_��%L.~�J:��t���[�@|�צ�N/*�s�@&��p��� �=��|~���
���$?�e�&�x��h�G��[��zǳ�Y#�a�ƹƯ��q��x���q�	BB���N}{��5x���i�Tj��}���
�ق,`��&��TI�<\�5��;U�*2�¦ロ�Ve��p�k^�M�\���R+vy�\�&�\	�M�/2���x��!�~�ZgOk'9t�h���E=0u��x6�i��Nʇ��e b�]��4я 9L�k�	��6>y3�~����9�s�v"Z�ƒ�+�݌����D��*�)	�����i#�P�����"� b}i�:��5�@�#�ˡ�6�ʣ>/�����/qO��x)�t5�SV�ؘ��i�G�-�w�c\DA	�gk��E�3"sV��a��@��^�<\&���v\R�4^���d��ҩb(^��һ��I��d�=��o��c;�"d�/�6@E����ļ������V�'m�F��2r�8����p������t��k.�O�-z��[�N�r�rR!�^w_IQ�-0��HᐼQ�'��x���e��WI�M�7C�l�D}�@��1_�P�)�O9�t���6�^-xi�M��^i��)H·G�͗��SPXKԔ�l;��N�|��B��8�511\�e�e�,�<{(��d!nSu�.�2m�;�g��p�t����!
[Z�o��Qn��@T{*���g6�e,
��;�|*c�M�&̢�ßlJ4 ��q2	D����x��i�r/������Ĝf���k�"p��lj��q�~�X@��ǯ}���(3���2�`���z�9�	����Gx�ޓ�TOߑ�K�|ԕ�K����;�P�%�B�
�/�܊� ��aԇ*C,�	�A�9Q-x�&�M#�.�2$߯Rq�2�轋c����ګ�h<Α�("G޶sc���?�א�y�K�ʊ� {�P#�"{��߫�_���%Fo�$��	�O�����=��_28�l�|�|��D�F5b4iSo��Ƴ?s�|Ű�R�_����� ZI��ݙ@����H� ��T�/�n0Xp
��@/����^�Yڵҧ�ؤ�d]J��E��P	�1�_��P,�ՠ�n�hִFn%�z��
���`��~M������3��)|�[� �ya�q�)#	��jl����0�!��?�zH͙u�y(��H��]�,ު#d���ѣD#\�A�;�?� u���,L^1FB2�Mo��[�%5�UϮ0�ljS�/���P��uq*�	�{�v���.�=�h�iK�O�O��㏍��{VbhKK6[�CM�`���e�n�J�������+
&F��� ҇�+�M:��q�Ě�S:c.J��~jwBI�ԉ9�j����.�c�`����>
�Q�_G�6i[�8f�����f��lJ�`��ݳ��^�E��'fw<�x�n��$@.{\{g���c����n(�UTw���LRvS�4-�(�;�O�Vڴ\l8���@�=�������u�7;�ҵ���U�D\Es����9E�7W� %__��TM(���b4X [���p��S޶�?�*�8�[���|1���$ױ�8�1A�
�Rc.&�uo�!}c��Y����X�C|��b�m��!Tsߓ��=O���Fdr��7��o,�s�;�����(�($���Rλ����>C��$A�D[��z�^zA�r��2�J�����	شY�%J����u�6_��Az������k0!�C���j��S��Yu�;�#î)\�M�E� ��8�q�- ����G��z�8�G/�3����甑GJs��V�G,?�|�|$�-��s�B��y�l�\�ؽ7\�x�g�����ӷ���;'>��&q!��3��/8kT� >cE�B�׊|נ�aXzc4Ϲ�L�r�	��R���{���g��μ{Y���1*h���,)>z�5���±�V�*������g@I�������\����W�\q*3�-�PMQ�K��Fm��Sn�n��EK�hA���]�}EJg+��26�D�OY���hZߍ[\&�X�I@�S�%97O�������p-�� �p�HN2�����D)ϋ䝅l���>E����:b!}�>�7�q��Ϥ$�a��|���'[���,�\'�R8/�]#1I��)��.V+E��"sAs���s��s�bo������RR����^�h��2�{���Bi�D�a���/.:��Y,H��y��@΄=���?���`VxW`�A�S�K�Zú�Rk~�g�6 �Qꊏ�c�*��+�?;�D�7�����s���P�R�2�f�F���S>Fb�"��hN{
�P���& <��2�қ�
�j��z4�Mj�e��UU����Z�z!>�V���^|)Փ���A�R�����z���ǝ��Yp����� ��������w�5�}Tv�2�_�������
3i��:��y/#��z31�8�6�F%��Re��]`d{���d9�w���N����*�}�˥��+���>�Nv�ƌ����?����@��P�DF0���G�d�Y�pY7��	Kf��l_-BiVS.�4[f˅��I�4rg@i�ą@8��u�-xnK �XK=��`�jO�ľJ���ꗇd/0_��!�d^c;��c����-�2����v q�>�,"�٭h��n�d���?�5,��肍}���Z�c��7`��}�W��`��T�T�"���̎�[֜�TM_�p?�]���;
}���s�����8����;���8(BW�	>:;��1̫��Hx-	�G�f��@��ɯ��� �����rj/�ȇ��	�K3�۱F�C�����n�x�H +ܱ{�H�����f'�G^�y|��}+Y�Z�y�ػ��ߦ0z�66*�&[�y��_Ղ��{�4C�v�.�A��"8O 	��s�IT���]/9�_�����K��؏8^��XR��TTyFi����#T2�M�7��Yxʮ&by�)U#��2�����t]Vd͒}"5���DV~�nq9*�V�o����ne}�I2݂Ȍk^0�4��Z�䙔����u�}t{L���o���R��f�|IyO���Y\���z�5��W�u���-9�����8�X���g`�� �p�i���M�� ²:��Bfd��v_�D�lH՝-/>�$sZ���j`�:e2m��nAv؇��p������:NEx.i�Sr��v���Vl·�E�;� e	"sc�ecQ��zw!���jmO�l��t��,+\�=�C�dѷ�M������@M�v��]f2����t|����X��-�u ��I�GkE~���jRl��e\��Q��5ӱ�S��pX(�O�[X���X�3ƠΜ���^�ɑ �G�h�1�Sګ��.�෭B/M�b@���[��:�3#<�������\|ƣJ�9M���X�^j��[b:�S��Ao�&��H*#5^�k��IX}��{�Q^W6d�N W�\ֺw�|)���-X؈'���׋�Q ����\���P��giaޔ�Yt@��n�4�u���d��`'^�V}�bi������i"3AE7F�%eln��3r��yڣdq�j�� �����7Hp�abk&�D�X��r�6em�|1�$�;8�I4aP�{>�,�戕9�Au+a�-�nT��@����!� qktIF��7�棳�Ё6�k#��z�n�'W�a��^/w�p%�O)�S��*�kS�)�f^ �s�np�G�&ךH��7�ig+����}F&�!nvd��
��?��&>|h�G
�\5�X
��(��q�)��g�	}�[��{�,�s󳠁t��p�%Q�<��΢&���	qZ�}六t��r��j�Կ>���JJ���`����FE�.���b�Q[Co:gP�U�;��+V��6}�d��-C���O�[qU�A�|�Ѽ�e�dk�E����D�I���ܡo�|DR�~#o��L!�Y��FXG�5����\��:�JHݒ�N����6�"�ڽ��I���'{/�2�~�Y`�_�]��
Myw׌'Xq����"cN�N> �}�����)$T&r�{࢞�"s�LKx�'� �~����f����	�=.��󣌂���c�`مb��D�ǩ3A��xoN�A֠��B᳞��(�>��}��D��vT%-n&Q��S��#��x?? ��#��	�+�E��-��3�8��n�)��nĹ��c�}h�i��Wb%��	J��'B�n� ��E���h����!$��}�T�z�9���z�e8�ٝ��҅Q@d=����Y��*Z�@C�̦ٿ[��r�=���>q�����tXS� ��*�K�m ]�}��8�#���t��+����ųL��B��$n�$�/K+lY|ŗ��!Uu\خ�ڀ�J�S�J$.>y(9�w:�%�U�7s��4��gzQ|.� ��PR x�k��A�a����r&�G)gh幩Q�� ������˒�3ī~;�t��Q�Ɠ��&cv}�1!F�B;3��ޑ�7���!_�T�v�D��t 5GJ4'�y��Ps�LG�\+_�W<~�m�������,;TM.	�b]x;�ϴ�A����������n�ĺ21]{�Jb>4��:���=l�?�Pa�s��eҭأJ� ϗ���`\*u�6ty�g�~2����K~�^t�����n�<X�V�# ��>�ˠ�o��]{"��(�W���O�O������w�K��2��b�v��r=b���%�ny��tL=��&Y+�G�4᭶��,�;�W+�'�%`��K)`|�(-�WQU�b������Ew���r�@�z$+a@��,�[�.}g�| =��~O��<6�%���s��e���i7���-?e,��/��|����_�Z��,����@Xŏ|`$� 
����Fbv�*�L�lE�lb%#m	��-7*��_Ю�7%�����*���{*�v�%�^s�I��y��D�4?�^�@��e{�\���Xݔ�2�P� �8S�%-?r����]}{�i��t�M�X0:��/ɯԼ���V;��%�Ϫ��86��Y���-�7�G\�H���3m��ʭ�1n��ĝ��b���.���8h�;l�g4�c�`��N_�@"FGh)�H���S,��}Ap�b�U��.r�z�-��0�1P��c5=�l9�~t�`F�Y����1�o����.�U�Ry$���*�h{nWs5eGVk��U�N��$?�
I�,�[��Rϕ4�23��3���+_�B����Ȅ�[�*�8.	�ǁ���Ԙ�xV���>*���ñ��@�ڼa�x50	4����J�=��D̿%��M2T��$�	����u�Y�x�
��	��\񴰪� �Akƨk��X'{������?�؊��q
�eZ�R� 1-V�#�3�#A!)�T��[�o;�D���#jvHc�Z������	?ӊt����ȧqm�u��;�Ң�9�$D}$ّu	�'V�ʺv���A�毠�m�1aq�4����Q����t�#w���]s�b����Oعk�js��E��� �2��/l�b�ꌝ*�jtv�3úI�?�9�H�QKX�f��+��:�/��4��3��bW�_��&��3+f�Xmqܝ_��.;@�.��FP���@-�Ƃ矈P�j�uc@�4*9��H�q���CnY��+"af�)�Gxpw��8���*-��RW�u�&������s�J�}{�%ɞ�qr�9H��E�Bv�e��a���I���ދo��ݖPC8�&CYz��b`5g�ڟ<\�G�j߀�ĵ���"�f���+���#��-ecf=e	���'�3�S��Q�n�lrc���v�`���&=�܋Q����i�9��f_��e���p��r�H��B\���a`u�+j ��)'-���W�O+�~W�Y3���b�cd��&���(�x P�x"Z�J6-C���Ye�7�r@bn�@��h��lD����7��eBJ�V�T2�x�D)��.�iG1���-��bTR��q��zm]u�pѥ:�u��������b/�B�-o��-�J��Ԭ���Wf���"����i�p��.�#��J4��Ϥ�=�*���&V�5���{�V���hg�rx�q�4�&�M	�z���Y�Y��߃̊'��[�n��������Q���X>'y��j�a�ا٪���{�&�l���W4�q[����1$�;��LR��s��r_LQ�pn�[� uq�=	��܈-,�u	sM������I}׫���tj��vDS�؍)%Av�:/�;����B�<1ٯ�Wo7�+�CT�_3�n�� je���o�|>�z�q��:�2��@�L"ۊ7�㕱YhJ��E��A��t���Q�o%����X�V  =ߋ�Ψ�f�'{&��8��C5h���#��LJ�j�e�lt�)Q)��Y�x�#�)۾���X���w�#=َS�8Ѝ�y+O��$ڬV�_P)L΢�4�u�̇.�N�v��B��u=`����������Z�3��e�RN!��1u��=�陸���A)����u�b���0xXM������3Ӻ���`Ҷ�m��:���s�@���Pd�lI(�@^������8��|O��ڴ"��G���-���v�p���o����8<��� �`a����e2�w�_n�u_!�b�h����o�����XBKW��Z��VV�)K�"�L%�ƨ-�:T=�$���������2��L�;�}�Yπ'w�����Tɘ��T։�����R�N_d��>& �H�j�?S@��&���F�,��2w9�m55ұ�eԗ��T�ħ�����b(O�4�=8f�gS�K~�JJO:�\!��b�J�� Q	_����>��(:��i�=���CƗ{�p<��
I1�'B����	�o�<S�K��C#�h��#��e�<pB����i�a�~�;	3W�����8$��fL��vks��C�B@�a3�D_�	�x��&?�+\�V�N&��Q�W�,�t-�xC�
�ܼ�5�����E��2�����*��:�Q�oS��IM��&�����zN�8�0i�4mrdPT�q�D�}�=�	�&̳�2肭$9L�*�wD����6��b���}����뎅֤�ү�v��r���D��H��܀%fm�p�Xtݠ�Tv�Blھ��̼�B2�����g��&�7��\�����ՔF���Is��P
�u�J02\�Wxc�����t-��d	���$ϩ���8�t�Y��0+w��`_6������FUVF���g���1�� B��|r�[23�;���0VE�v/ �,4m^�{� ��g�7�ʚ����f��)�����w߰�v�S1�&U����ċ�ĲC�6zڰ�A$~S���J���0F��� khR��P���-���v6��� Iq��b"��ˑ�1=���EZ?�$��]u�\[�:tr����F�8��y���g�]Zʤ7k� 0�����m�AP�$Y�>s��4dCbi{�eVl~��܁��li��$(�+f��,���Γ�N���uL*�o��q��\A>b1�,@/D���T���a���qȐ�7�
�ӣ�����Uƀ�J�D,zO��(�`'ezB�:c�)S]w8�����[�����!�/�3��f	h`��5@�z���{b��Dd�$ qi�����L��ߒa8�d��ݏ�S�$(E��@;34@�2�������PvJ�����N8z�z'���9�jHb~����4��~��,��Yb�,������gxwi��":�^��?�K:�Wmې�V	��1�Ag�.�XB�6�ʱ"�f��g�fveI�����1�!M�O����C��k�� �i��Q���87ב�L�N<>O�����y`��/�K�����C��aAF�bf���B<�Շ���^,�ڬr�s|�M3ؤ�ʄCG{]ۈ��@R�X���tv��Kv�1�#���:�����+1wVdŰ$�8��{�{%ZtQ�d������Y��éE��������`�*�=h躙�Ju#3��!ϷBeS(�ޡ�S�d}`yy�|��&��#�SY���S�]���[�o�<dj3Y�x�4.�	�9l�l�FT]VIhU��V�fp����NF?ݝ������� ��+�������}�)</
�+7��v0�(*7��Sq���� ��%┱���+�%�F�L����3��xJ�k�żC�a�o�a|%R:?��3-� *���1.��|0#2W[K,�a۽���F�i2�~WBc�*��n�#o}�J�I�Z��/���6e6�e(�^�9��k��},"�D�)Ds�2�e�g
_y�z V�x���TY��Y%��E��0��![8��35R�-��r0sZ۽�N>�4������X<MF��V�lE�`C-��x�*l��sx�0�R'���MC��Z�E܀�������Q �Y�9O\�ק.e���׬#[^7p�YqU^�#��A��[c$ofaY��Uj.�H)��B� �p�`�E�'?���������j��[:�����k�W�A<��mZ�UD(���w����N�� b�x�s���Ȇi� H�8� �������sZ8k������^�
S��B�Y���O�\j�5��1��8��S(4�SG�{�w�ƃ76⥮8o+��f��)�p� )6��1�&�vZ�nYJ�@l�2d�{Ů[2�O稣.�K��K�]ԛp6���6+�a�����ȋ��Н	��Y)mW�f]jޮ��W�����5�e�8�Z���	rM�ܹj�����,V'}��n"ka3d�����H�/�%˸���}�M�釺0g!@0e�]9��;z�C�Y�&,�;Ӻ@J����R¯U:�_i��38�N�}�k�y�_/�/@�К�����S�,�u!k�;�o",W����9.�+D�3(rZ��J�8iI�
6�>N��?�4�c�>挲�¨1Gų!��<ǰ����8.w'���f�v���]�_�Y�},×��X.̯�յ��d��Eɸ�/i�G�D;'2�2�P��Gm����ߵW�Aq��L�����99E3W�䦖��C��2�V�/�����h��ǐ�\����п��B!��z�5��L-&P�#⬹!!_��+�(��c�?�5�i� 
�辋o&	v��Uطq{3[��x�%�����(P����g�����ݶ�dhXKU�	RԯKF�s��|�feiڞhs	Ccu�Q�b�tK-�,��g�u�9$��x�& ��bT�,�X5�N�ʜ�l�9����$��y���,_д�r���H��x�u�qS�
7%�đ���(t�/���Ü[
��'[I�x�O����C������:N��&瓗��Z�(d�ȃƻ_EN�l������?�=#Y�C�fC�r?�5�1��u�&� ��Y��P�1L�&9�9=/�O�D��'Ə�QgX#77��P%HU���z�h� ��+�	J�fMZ/���ubV��2����%_3��`�o�i�/`���q�2U��i���%�.lL�MSV=�8��^�
��5�e�� �����c�U 8�V] :gw:�����z�&��|&�6JYJʂ��j4��6� @W륜B�NT@ Csf÷����ڔ�h~��q�k�Z|������G�D��Xы���&��Lq
`�����6��RjR*S#u�Y�S(�q���:L�)�f]	g�s%�r��͒&��n���e"���.���v[3;��a#���)6�9��u���}��@����� ^I��6���G�ެ��%#;�B�|e��z��H�p"j�k�� �r�����I.\��Q"C����GhqD���Yv�̴IT�T�ǜ����)�]���~�@�s���n��X)4�$G3�_àT5S�"�>��U���S��?�◥���p	2�R�ׄ�����#ܿS7�Z��N-TY �Re���� ��"�q*�H9��t������H��Յ�é`���u��^��� HH�{<l5/+>9!:��GH��_K��L��Q�9A��k�Zh	�`��r�}} �з�&3O��ٍ��NR�A☹'�J;�d�&���xo�%Gh����}4�
�QS"@j:� 9�o�4����S\��)9���J��`��Nt�;]kk��kM�d��O�.��`Ց�,����pW�7j5W��������?�:�ߚS1R���*���ТG���R�ODT�lș�:E�Wn�'��|��tqOt:߱V4w�M�,=U�t�!7C�W�4�u0��
��z��S�#Dq
��l�oض�gX���B��#��jR:��t*뒾(O����a��M�p	�8�c�
�}@'LL r��,���C�4������<wQ�76�o�����Z�M��`
S��jN��p<>�n�SB�����¹𪛰8@$��Eh	�1�x��}�[!{����<�o`���33~���GS|&�|-�k�&��2q��Q.3��ӔHB�Ţ c������%+w/,���ŀrw��R	9�����f��p�¦�3U]I�c��6F���$�}eאq`E�mҟ͊� �@�?���{!������O7y~�:ڡ�sB?����_�h��`d`tW��x�N����:v+~5��Na�P������+JO-xI�1Kt������`h�=�,���g$���K�0/��'���v+2��rr�x��? ��ʹK\~�>*��\��X����G���È
��������r�r��t�O����5�+��lz���342��d�;p����w�
 �#�E�q��PO�ttA\�2Ɠƙ������p�0�*�=�!*� ����	bx����(�Y�,��V��]���3Һ�h3"���C�:��D�����wÛ]3Z�^�Y�g���G�zL�$+>k���c�o���D��0��\�%2>�dt鄎�W>���>X�����>U��#l�#�ǎU��V� �l�����Kv"*�8�d�Rt3�a���i�5l|���+$Y%��z��Ws����W�_��XBa}�����c���8���Os~�gT�&T:�-W8d�ة������O��Fe����r�\;���Ӳ�p�2�h�8������X2i"��DI]���C�Z�q�� /H��\Z~C��D�]�IJ�iΘ�I�_�2=!��_��7C��Щ@���/_��<(�i�d"���LX��3�"%쁱�|.�ʓq���x�O;��j>jĆL��U��O���I��^Q�L6^���x��BC�Nn�~��-"�3k|���{�8�������z��⽯W��cID��dt��=h��'�Əx�J���>���h�`� ېZ�!h�+o��XX*��Ȋ�G>����E�Ϥ����(U�  )	���y|�O�;���Q��Z�
p����n��1�0��&D�)���KL���5�`8R+�]��ۉ��&}����QƄ����!�;D���F��Q��\���c��#~��)s>I0���92�qf�� �?yj�� �Q[���)�	C˽C�ɾzp�d���t�G=�,��l.���'q��@�ues�:êW$�����i���_Ҕ�d�/�g/�W[���,���
��.�hʨ�U^�x�����}�D�\��8����f�r7�yru�k�ɚY3�"X��)e�p&�V�����}Nꤳ�#���`�yZ�[4��*�!���R�5E!�!���p�8]Έ�������e ��Š���.s�7|nۤ� }�YQ���G*R�A��`n��Ax���T_{i�K�9�nU��A��b��ՔF��[5F��1�h�}$�:{8Y�?V�$z*�%�c�`֤m�;���_+�����V�04-3p �a� fe�o"�Tz�n{�o�c�F��CX4EQ���;f���'/0vAi����K��5
��0P������v��X�d�n���^pOMj_w�Q�6"lZ�8�^�i�ؤ@T��й���q��q(\�M
!W�
�
���h�����})u¿��4E77i��iM�Ԋ]�c�$��΅8]�H)_!h��"��H��tO�"-�u�|u�U<�qu0O�h:���&/v���^\Tb��)�<�� *�f�h0�&/^a=_.����ΉV���p���ms�(�:�{2B51r��X�E;�V���Z��l]E7/8�Ef�AJu�7����'��8�7�O�qM*s�?W��(vq�?���nz�t�_I�z��&!�"2����W	������(�@#�A�#�n���f����>Ȉ�9n'�����Ƙب������Y�0���w,F�V&\9K��F��/�j����V���w!��'�T�4N��O����Cר<�����!��ˆ;��䑖���vCj��˟�����&������������ϓ��o���W�����]N܋/ͼ+X�+u�v��~���*~\S'�(&�Jաȕ���_���8��'{��3�g�W�Y�UX�˳�_h�s��w�.�����'�?�4��Q�k�1�z��|"����p���f���nmi��f�W���} NͭmA�	#3��@�Pa��Aŗ��0���W�L�Ԉh>�:Ei]�R���?��)�X�{`%""(�#�Qj����}��*����,���u�c����c̪�
[)�_���Y��V�VdP^$Y1��`q�?�|ۡ%\+�� 
�
�-�C�s�&�Oklϲy��mCp��U�����q��н�nI��� ;O"�o���zx��r�n�}	|������qj��=C�Et��qS�֑��bK8MMV��+�ώK��)������&���B���ou�}����}���d�?����Wa��E�-�$�Yp�qm�lJ�d���g���0�6�5��*�8Ӡ����7̢f�`��S��I�2��"����v�#2 ��\ Ay͸=��z3�U��Q���k
n\���n�X?R��M;�n�k����=��~��r{�R�*�3G��R���$������W�ee��72T�m���)�a�D��v�3��y!���^6�_��UQο���y�7X�(�.�����i�B��̔l%
_1K㈪\�T�Y`�zu�m�ܿk_�u����`�:�I�51��IJ�t��f��9�|��tX[IU��ZÜo"�$�D���P��.k�DU{�5����B�)�H���\o[��1�.d��0�i��;��N�*@��g���,��$��x�.�F�d�[���80�?�k�\�J��g�D,5<PP�src�yP�O ��<�@NAq���ֆO\D#-nA�o%��ņ���T"oyQ��!����v�c�r1Fz�,00�dF�k��"���}z���?���x�$yl�1�[(��-fP��DW��S����n0��`��Ys�|�������N�l[R���T�g/j�R��ٹ��0s'T��<�>�~��b��S�?��(V㻛5eT9V���9��58��I��A8���r��٨7�6��`_6]����"q3H� Id�@"� J�BS0��<��I_���QH�M܄�*��4_{yhD��!�&iy�Ǚ�dGO v���[7�����s�$e��f��"$f�OcZlO�w�ڱ�D�/+�%�z�����)�/�0����l�e�����B��Tq�_�{��Y=y�%�Ȼ���
�du��K�0^�H��Td% �:T2�H6d���C}��;����b����ګ� 80�:7���"�cܲ��{sB���8����A�82Ǐ���kݻ�:�s46L|%���#K����S-%U��ꅢU2�:"��������*��v(�]~v%,��i���Hk7#r�Y������2�a&|�s��ⴀ���1t���p6]�<�,@�l�u���Z��lK�XI;V�^`�ܽ[�8�����_�u8��S��.��^�~׽��j� ��4�C_��V��lS&�<�<���Dt���s�k��!�5�����qe������7��k�����T�H~ASG�Y�{8Փ�4����0�Q��^��н�����t7���%���q��м���\�����՜V�k��\W��jh�L���!ܙ��K)'X���+��A���OG6`5��eu?�ҕ�-�j#�����T��Gعi,��$�%x7����<4��m&�D�;v�bg&��W����;Ϙ`�H�������"V�z�Ȼ�����/F�)7/So���A�]{�щ�6x0�$��^���_�@�����ߦ��)����<ԧ%
l�\��._�T��!׃ky��I'�4��~[	�m|@:�Ѓ?׷\ ���R�|��Ω@���ELqΧ��y}/�����:�e�5(������xq�Z��&��y�bST�Hk]�L9<�2V�H�/�%�2vDK�N��D ��,	�֟ьt�Z����PRּs�*�~q@�ȸ�g�@�M��`i��oV9N8�!a�7��'�J�!�!���%I2p�T����o��_�{y�([�R�e�D��N�0��+�uzh׾Bk�CC�J�"6����W@�b븒Y|גӄ�i�f�?�<0V����c�Yi^�4Mf7rz����,�`��%!�=��Sd�ȼ�E䘊%f�'ʒnh8�}�����\���c�b�{̅;Rx\K�\��.e-���3D��ZϢ��SX<I�B��M=�?��b���	�7�A����O�Dֻϖf1f��	i��["e1%Bg\���W�b�p�u��`ն޲�ZD̕L�`���4bQ���V���1��6S�Y���溑��P&g���Q�z)��-���f�x��ߛ�Z.˚Hz|9YM֥0ޙ~(�,(�=�h�'���ƍs���(z��g5��x��'.�m2��6��֦�[��,����`��7�q2���F�^`��R#�X-�	*g�O�"��A#�A��2�chm���хַ]�xay[����ۖ<R9��&���B'ק�����vTS#IB�͗���F��;�\h���J<�����J�K.��.ڽ.�0��)=��o���`����*qF�2��	���5ܚ��Y�Dl\d�4��s�[>>�1x:�[G�����K*��Gﴥ*(J�B�#:z��9����t���h
)��y�zt@�,~ܓ8��A[�=Q��&�����<,WȪ��Xbq�d�_���?\��(i����� ���@�cg���E$�|uO�9l@v5>V��b'\��M"�~!���4���ER*b�'���^~��[�+�M�,�8��M�=��}�N��|j=x��5D7著���K�Cn�7�����	�ذ�Į��9��km�ߛ�������3m�9�b�]EB��N��~z)7�$�V�a�u!Q��a1��ijo	��1���9���0�oX����%��M�������6:L�}�LM��}��c��|hp�oU��I J?NB8���	��ᦞ�5�km�I ��pѾW�s�e�NА���;J�g]�@����P6�/��,{k.r��Ĥ���ت����n5�� č�\��fO����Q
؟<��Q����Ն ��8mw�IuR��'�s��p���dZ�C�wk����F��^��O0���;ZU`%��J`��t�m��*-�f����A��LD���x Nt��k]�@S�C�fUM!�o���j>����[Iv?��{�%��4���\Ju����V��$,���)��&�ut�SD}�H���*��Չ�Eɢ�9;'�'�A3�K��rJ���fdl,/��k��rq��|A4�8}��K�Pf��rV�!.x،]��yD�9�=��e2[F�:�- ��K������o���;U՗%�;?�D��oP�oB�Uj_��Lr+�p/ !������=��I��_���	�r��k�V�N��<ϔX��z?��G@��:�ά�<�|�fU�6���<(D`~e>Ҡ�ݺ��qn]�&��]�ҕF��&@��&���yH�L�NԠ�����!=�(<ܰ�?����#�n"��?�5y�ܷk-�@L~���j���|�pC��?A��. E&���&������2 ����y�7�Gphbx��r�7��ns��yi	�~�D*�l�f1�Ih�����pD����+��t׾�&9	[��:��30���_�.�/$��kN )o�L=��v���5L j��T��:��.ͬº˹_�e��(����v��Q �S+;&�|rSs�W�Gt�0�3�1�F�J��&�#��^����uyV_b�!d����l�q�/�͇֮���w�Я����VU�vCh~g,��D�B��ˊ!E�����Bހ Ɵ
՜�����.?�Xo	���5't���Z�`!�����|�`��GO*��	�aF|S���Uў�z)��:Ɯ��b��^�S��<8�d&���U��b����MV�.N#ּ�+5^mE��a��g�x���R!�5bSą�5v���h����H�&qu%����^j�%|�YDn嫧-Ż3>a