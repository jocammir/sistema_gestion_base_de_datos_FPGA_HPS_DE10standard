��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0����&�#��A�>D�#���� qX.�[ �qB�FG-w�~��N�<g�3��*�u�Ji��9�������_��B� �٬��*�1��)w�|{����&ɵa���Ԁ8JF�ͶM�^8���k�+ˎ�lE��`q��2����ߖ��F��t�7 K���La���`��D����v��ȟ����XyA��p�*��Ҍ�d��J�pIy2��nl��h2�T��H�I?�^�+�jD�^��,����ڶ�o�����V[���w�+	�H.�xa�/j��z�k�9/T8Y{0���Y��vD^�1A1�0'Cx��Y$��BUZMOFϙS�H類˦�yg�}����F�b��t����7:�%`vPcaup���J޶���,"�|�K6��x�D4U�"��ۻS�%�q�@J�F+T%2L1�)�v�Y�;A��?�����(@]bH3�CipA�_jk�l6��8������=_�#�M��j���6�
p�q竂Թ$�ؑ�^��Jl��[�S:�Q����MX���0_O�~���#��sL<c�l%�����l�gFs�$��B��m��'7zK���	���f�>�ur7�n�5#�	QQ��%o֐%P`�D;�6ݾ�l�j��,~�P���ێ� ^�_������ �RC�j��Zˁ!�ܧ�@:C@
�Q��z�x�5����W���#8B$����=�3��K��vH+�Qٮ���.�Tl�pG�U�*���)��5�b�bEu�:bW9�s��/�E)�>���'`AN���fOߺ�ZF!�g74�WBw�t��9�VMm��&Ѽ�`޶P���$�[�/��{���׊�.:!U��ܔ(ră(�ݕ̃`^��U��E�\��y���8�]��)=��|����5�W��VAI�c?�z������D��=�^��w�r�V����^"N�O�`-�y(Y"�y$�D�Dz��.d^�Cb̬���Î���a4L�W���Z� O�5��E��1ߋ��o��.���p9��"p��bR&`����;Z5u�e�؃��!�t�T��.nN��/laM�/�=� ml�	��> �>U��4L>٣y,��F?��,��V�4(�������R���)��q���Y����е{��L��/g���7��	>Rto�]��L�jq�{׎,L�wFg�kY]����|�rl����F-����	�t�|�T��'�o|6i�.���z�[
��(\�2��OG� >P]�&D���	yxܺ�xJ׃���ax�^�~��S�8�m������quE�Vw�V� =%]��B`)��Y�t[=$��I�RЎ+}��b|��ć�j��D�K�\��-��*c�����ZX)pE�Ї0���V�0�0�/ٮT{�wy҃�J�?�@8���䝕���|��Т]\aa.�8F)Z��rh��q�&*؇�n�U�$��ZM����^��/݈M�覸5iU����}>�}�zʷ�,��C��ߥK`��Y Q�ת�_�y����-A�%W߳�]/o��D
���x��ʉ��3:d���"���¾��gZ��H�?&��=\e�O;|1�`�CG�	���2?
�i)Xǳ�gΒ�X�>�A�wt��:�Wn�aMB�S����3�7����Ã�9]�s�ͷZ)�& y~Sl�~#XW=��h�jZ�����1�k�=c5#���������ଆv�J���9&�Q���t��/؞�,�9bH��|��"�wCɗw�z�:ҽ����@.��D}�!P5��γ�$B��^�6e#ء�>�^#ТE�?�+3��qX,ڤN?8f��7���a��'�:���@zV���w��m�_�=�i�<�^�isk�	H'�\�B��?* o�H���!}�x�ĕߚ,?�W1����B�n��@����&I|u��(��_��L��ԐBXS?Z ���U�����!G�w��i$]�(�'.�@�2g��D~��!��d�Ӵ;;&�&ґ�$�p<f@��_H`�.V��A�L�Y�W�������E��E
RGUa����`��0���j��ՠl�N�	����2��ՙ��wIiMu�]�Ԛ�J��J�����lD7m�Ew���X��*(�S�':sY���j��T���AA˶)�7�m��f�u@�kr����*���X%�p�r%���br�>�$kIjs��0ڞ�L�s^��s]����8��M+е7���B��~|9H0���5�q�Kh�F���,�t��J�?5 �e�ׁ_̜M.�ξ��G۠<�;�x��knBQr����0��R����oY>���kjpx��==�:n6}�In�Z���QĬ��������*�D.|��#��F���̤���5]<�LW�8���U:��>��C�4Jv�g%3��ƭ����o(���M �'�  W��i�@��Kq�+�W<O�/�s�uT�x/4��������
Ɏ��C�%��i���c�J^4�(��eV�$@]�԰����U�_�w����+�Y4Jz9�rM`��P�� "ڰgh��YO� x�|���(@Y�{Lۿ���ݝ�~æ������,�F�����m&y�����~�����gh��(޸�C�Q��Ӭ&u�1{�,�-
Np4�:_Cfūoꔝ�$����j'j&Q?6���@�&FV�V�ӞJs��1��?lʆ�D�L���owF"�;�b8�$�8�pH-!�-8�!qɾ�/���0����2ύ�R{S>  �}^�ӏ��iӏvC���=9� �j�a��E�-ZR�d��|�ܕ��YJ.E8Ӭ缒=/+���
V����ul�-����ڴV�<�����l�O�\([��,ah��ݷ}_��o��1�.�����ǈ1��S`H�RK��
�P��x��s�yT��?���tf��y����!����W���h�����bzZ��5�jsa����X!���@�tFPgA�v�@B�;Ul2!��~9�~�H��5o.��� fE�U�a��]Bͅ��.%�q%�ED�
��u�^�J�3O���5���L��C��d�2 W0,4������w�oT5�<.`�K�u<�)�7&�v�I�lE8f���A$�b�>�cP@��tM�F�`�5�4;o>���"�z@� ii!;U�HD����@�-�6FX��{>9f�?2����ƪ�p�h}�\c冣���h�O�/L��kS�* 
�=Ì�J��bN��0�ۻ��iq�E��GƆ�`q�;��boq��ؼss�q�ݿ~�0)��c�bu�;E ���M��֣�S��yb}6� ����{D���5��>KUF�J��k�U�H�B��&A�Ah,�"�>�^�US�[�#����U����h�|���I�n���	Fd���FG�ś 6Gl收��O��-4�EcC�0�*������1lb3�Naϥ�5Ȏ`49�kY����J|�)��Q~5�ء�FU�6�MbMTY���c�Ot� x�h=_zD����� �����b�$^�?�?A�Ջ��{�@�jve�_��I4:��w��l��v�dV�����#��}Ov�f�E*�g~ݛxW3�3ߦu��3>'z���V��z�`,M��.�H�@�$=r|�9c���}h?U
v9�
��-
@,p���)���P�1%Ų
mA�9���Q%�6��[�Y����"�c�G�]�Y����T��{|��.Y��\�=�>q��[����y��H���bO
;KE'���E��D'Y��z�2�p���gf�j�3��{س^��۝jq�q?Sd7�����Xl�0���a�$l���
�a�1��?N+��D��<�+�@�� x�c
����Ϻ�3nZ����7�����c���хQ�'z�V�8��Z+��K8+�ł�B<��܋�2O��;�+�r�p�7�?�ooM�37�1�.e8�+8&��NoS�q��G)�4h���S`
`�2�9�|����j�{�pao�u�wo��i
��ssT��Z}G���B�{������t�?�П_����A�u�8�]��$C�k��F�Ć�s��,�X����| �\�D�q��Y��W~y�ƅ߈�$��ҳ�?�5��j�"㳎��Q�I�";��`usq������/����7o{�4�k���/�`�;{�Vn����a$/�v������a3�Xߍ�R������拉hh
`���*�]�v�L}�Kw�R[ N�襻02�寴��{�;��n�~B�+2��� �x$mT�-��J3�wma����F� 7�oX��7�:|�-��OfU��bBD�����M��Z�Ti;4|I����?D��H�Vz���P
���Y�0����?%gJ���-��;ΎH_c%��$��.N���ry3$_����D�H���V͂�T$3�f��kk�B+�����팴R�\AnEH�~������;D�vL��˿q�l%�z��#1͈�8)\��o�yy�M�g7}	n�3e��ʶ>��sg�	�򣗢?(���x�(����\wΪ��i���j��%M?�C{5�����Wi��Vlc��߾ a��.�o���v��D/�W���YD��'c�-O�x?��>m���%����4���ת�\�ջ)�ʩ��p&�#���T���������n��n_�E)
sՃ�_�"��6���O�,��J���V[[�
G��hĀ3/��IO��r�K���T�C�O��fT�`���t�S�P��/q�mw�:�'=�f���zg_A*���%+(�# e���oGˢ
̠���o�PF�"m+�-����P����)&rBW�����x��&��G[f�ox�dYvnٱx](�l�+1����`���7/���'x��;|�;�tS�~�JQ?��Qz�lS��ʜ�Sh'�)��8���?�Oc]�&�����)��K��Ay��N|��H&��n&$��� �$�M"�q���x����kJ������V@gɀ>~��N3$����%��>���i1��~�VJf��d�7fg�ךgK�b�:�,�J��L��> ����X_fx���0�S,7���8�uA�&z-��w:+����Q��P��F�f}��X
k��p��V%?�0�f-ݭT՘��Ǥ���_i�>`3b�T�C������СDMhX�8�a8�:��v��&�\&�!��Kx}B�޼���i�V�uj�:��s�I������q�HP�2�oE<Z�T��@��-�Q�JS���`��S����mӾ�C��ԥ=f`�&*��w��f�i���G��TSb�hp��Ș<�V=�9S^��(-����1-��de`LFi���"�w0�ϖ1K�p�����V]?:݂�e��Dp�f?Y�w���H���]�S����P�i���V���w�Y���є.]��2οw���ӑsp��ge�#�h�\��=�hNS�E������g��������Q�h��%ܞK��P�}Y��I ���?ޓJ��l���80�RD����Yw�HVa�ԛ9G7[��ި���v���?a��	��&:K}C�PH�؊��÷�����ғ�d<���D���S�W�T���A��>�zÀ=y+$�)-�44,�����Дf<?A0g[/��2p�u��5Sm�_iZ,�YJ4��E��bn�������IM�n.�����ɭ�&�ģ��K\���OM����.P�N��!r@T��)M�F��?�� k�|o[��?�۟��, ��A�ئ��oJ~2�\t�^���_~,�)f-,Y3��x�x�n3���7�v�����Q�Oq��S�bg�/���d�����V��lq�q�����~���	o�l3A`� ����$���Xη�ڲ���_��K���f��Z�"����p{��H,�: �/QJ8*S��H%C��IkP| 2���7�[[6��%���2��{Rb���o��)(d��J.��P�^��*��_7;���I��pu��u�O���2����n�{ZZ0L��0��Ҕv1���?;�����rv)*~8J!=�8��&��j���Jl H�Dd������%4k����a	�Ƴx�+�ߙB]=tvv[�`��l:���"(ȕ��\�<z�|̼�w��.�is[��GV�6��~�ä��#9{����r���W
)�%�i9c֦i�������d���\�@����y7=�
�n�=���x� ?�_&aww��C���� �\�7g�
���7���9ط0�)�����I��t���jW�����9e��@J�7ye�]'^��g�sL=d�tk��}6I~h��z��e��>�#9y	�5�#�dS���sȥ����)26K�!�O���e�h}`����C���I��K�W��gn�4(�P� ������j1tג@ã<�M��>B�lݤ����M�����]�j�6@�ef�K�ɡu��"���.Q���K*sH��8x�H|���� j����,��U3[�4&�A2,h���0����a��&��~�o�Y�8���aŠQ��'�Q�Cb����uC�(>�1��Ta��,��.�]��J��E����
���Vx�x�̡���.�lWJC6~�hG]64y�FLg=�f�!MS�1���p�&�d��ࡼ"��bTs�s�Pb|ܛMA�+���,�|
P�C�~������m�u�O�<-�D�B˕iH~~�8�&�B��۵�8�	�PƔ�q%����{����Mx�cL绊��N=��q<=Qi�5d��t���.�H���Y �]�����}�(�;�R<׏���멐�͔�\G!���[��eNK8� �*IoJ�[)Cx������F���/IHUW��j5U�]��+��<��U����8�Cy8�WBw:��|�9��?�A����[]������Ҏ�=9�H�l#�m�YvRւ�5�
�L��Y{o�姭Q�_�����1���X~�f�Z��W�|�dE�H���lX��%_�θ����؈���A.������f���$��
r�Z���F�D��=iU�I���X~��V��-7�[�;=g#%V�f���ojLg?�p��Z0Z�6oѦo����}A�Or�i��vP�3q�#r���G�#g����I��2|�`_������ĭ�j�\����X�+f���a7���v���އ@���OZ��0�4�U�Q1"\@N���`ܲYά�5:d�K�>��^�����W'���\%[A7�����5�(����l| ��Xo��Tݣ�CV�~Y� ��0�	��,;�v�k�0�CKe����pu���lj\vz��C��2)��Ջ�*i @٬dE��Հ�~.F���>1�.���_��7�B�I��]v� k0�Pû��W4���H�'D㣽��%p9Le�X�$k��$��,�:��˺^S�_�y��?&ZC�Қ��W�\g���c�o��m%����9�������fR��k$������O�w������)�||��p}����v���e�aUɍ�V��K.�����{�F����`;?��\3gRv{3���؟�Pl�
*���ֳ@ �=@4�.�y{��NW�]�v��^.pA��u�~�h&���'2��P��[�M�0���<^�����8����g��0ّ#�iD��QgjP�T��"c,yO�QK�'�$@��}����ph&���񖴚<���8| 0��A1�Utg�GWq�=����x<<��
���^��߇~1iO��ֲ�}�i>� Q�����*+�8A�ߧ���� o$h��	s
��f�`L�oe�i1��q!z !���B�a�u�+dt�17�9]m6�����A�U�;E�Qϰ���瘿���z�3?~!mfܣу� �(�lu _�3sI{N���a??e����*�j��5ty䵊x�VQ�[�01,�5�VRB>�邴R�x��_P2���_@�(�4�͓���,8�e'��c?��q�A���(��qc�g%�z>$4��B��;9ܢq� 25í(G:D[b�Q~���	q��?�,�d��!��Q�4�su�R���F�P�A�V�����`ߟ��X-᜷PM��l��hMڌ[c�&Qm��Ye�y#� ��d�K3�g��m��é3d1p,_ˎ�	OO�Ak2"a��}�,Ҙ���㎜�A6�H��d(h���|4�W�؀�CHæ��_R��T��d�R,��@&WG�[�,�Qg�7t��;{0b�2�OhH\t{Ɩ<�����v�NۺKO�P;�;?��dJN�hC�ݶx���ז�.k���y��-�:��+|ym�R^�z�b0�e�V��e/�R_�]D��z%CIkoQͳQ�ѣ�G{Z�%��D�{w-Ĕ��z�������I��N!�ڇD��+���=ܤs/��Ƒ��ѽXA?���e@֥+A㶨�\@�p��\��^Њ�W�G �?�n3���	�LX�����7	�_ޮI�
�T�>��Y�3��9N���UnN	6�U�Ne������e�sϊM������`��sM�K<1���@�/ķ����l�S���,���%���l�`�_����?j��v�Zc�B��B����fǕ��],�=X
D � �үK,7$Y�>P ���K,m�pg��F���P�m�ؙ$ϛ��5�w��Y^�"š��Ɉ�9��j�0�h'4��3�?���u��mZ�:��^Ґ_D��\q����G�9�2 �ߛ����v�=v�nۇ�[��`�!�k��8�Nx�)��FIZ��f4� ��ڮ���g��ΐ�Rށ��UC���.�gk���B}��PW�ek��.$�5t�Ć�aPΦq�֫�Q��}�O2��-)�l�#_y}�~��a�͑G�Le�܉ N�Ux���O%ʑ6Ajeҥտ�b��qZ�x|`��:]1�|��MD�kC����&��h`Dx�G*��%	>���h�$�i:�|	Cs��+�a'�	@"O��˓��4�2Oy�%1a����HU������ְZ��nk2���s�qj���D_u�y ;IvO		�<�|i�1�����4EZ�]��L������P
ف�p������|��)��А�uU�klO��L�Y�o�b�ώР����7�2�A)?5<��y?2|�1:�b���^���Qrs�C����֧�7Q�J�H�?�<\$�;93�2�?I�a����� Ӯ��,<0D�n�{�Z�y�܍=��V����>�RM!Ï)%�[?�����w#����t]0�tʴ��v���R1��#{��EI땂Vy!&V ��O�s�൭��fC@�[����Bt��.��J��A���	������P`�1ԗ�%q*�^��ㅘ��c|0�\.0m{�=Q?Z7&ˡ	Z� ���!�L[���Í�R�ڀ2�Kbch�L;��
px�d���hP:fKf
%�<183��a���	>���Mǿ��6�?2��������t����U��,y��=��t��7ө�}�GB�>��%�!L
�I���ݣ�����b�����ҙ���ˋ�̆��*�T/��|$�����A@ukKh����w����EO��&�K?{<�<�c�W���?1;ߓ��ؙ�v:�7f�7s�4�x���$�޼zz��l�Z 5���1`��+���R��R�,���ν]���5H;��q��_����B4��>�_K�y��K�G��"&�����=���B�e9�*�:�cB���B��ӒBk\<}������&��K�Hn��"���h'�_�z��., ���k�%�K�g6p�|0�o.Ӻb�\����Y�ө_��i��Y�CU���E����Ea)�?��5O�,�Xs�ȭQ-¿M<5n67��;6�2�)�yRd��%��2���v��L�����TƗ1�o�O����cV�fl�[��-}�Nl���0��E�g<>�i-��Pa�<ٍ���
uŦ���P�-p��m�U�RhS���=��i��u��,?�U?yYB�q��Uy��*����S6�W� #ri�.a�w#�p�z�}^�yd�
ET����'�OpI]T�(I�
1,AzR�/0/@'��IJr8�_�oЯBDȞ~���h���xV����r�yS ���lZ��������<\��I�±h��QC�/=?�mq��,��ۇ�衅�?x�O��D �S.R@-7=\����#ڴ���ż9��T��=Y��g��Xb�Rah"�1����4��c8�]L5H�]J��2�'�D�/��3׳(��I�G�6���Jcld ����is���s4&2���Ƚ
?|1X{�-w���wx�n����H~�����t��SJƱZ���E����v��|�>��y�I�Y
Ѿ��%�ؘ�㰩4Tu�$��^ɠB|KCjL5�lru*�����E� ��r&�/��?۳�Ǚ����q�[��H�x�;^%xF��Z�e+�N'V�]�P�3��g��!&�y�������"�*���m��;���3���t`JVRiZՒ��rG�q6�'�*�����
zg{������t[���,���\�ykKt���d�|�(�꾑����UMmw��s��Y/1�U?9`����Ŭk�JJ,Emҝ֜`_0J�R�-��[x��w6���t:����	&$��Y��5-��T$y��(
K$vQf�(�j<k�3`�Vg����Ћ<�\���1h=��=�7Z��!��%ڹ(���U_��'L/���F�F
%hAE�px�^�����7ܱ4U�ͦ�BF[�"���`P;Fk�����>�1���������3�Oħ�qgcV��8��ock���W�]��2�$����m7�	O�W�P�,��`2"gO=�)���T��}�TaQ�#
R!t~��[�͖��
b�; hI;�G,��g�[L��īx�hĺҰ
Dw 6��t//���B��c\���B��KC}�:��hr����ZQ��DsqK88A#��X��	}��͢�g��|Za�1@0���e�WX��g��*Q�!�58���,2g� �dH��Цށ!�L��_:����:T�������8�
�qKU�,|����{x-�g�ȗ�	YB�q~�|yxT_�����3�/R��#��@��^��D�����X����Sݓ���DIn��;�q��J>߱��պ���hS�.�5�Q�{���ɪ,�r���,Uh��ȏ�f/��@�� *__�*���q���n��<�g6y�����iJ$�o1��m���or/$0�Q e���X���g)�i�0�D��t�a�)R����*,��3�O���F���u~"�����m������=ʶ^YË������0��䩀 F[L������}�;;* �Gw��3��ͯ�tO���j�`[��zV�4ԤP@�,1��^V708gp�jco���R�KA_��&}�Ҝs$���C�T�i�>pj�W<}b?�����

����I:k�&�ge���,h1�Ic�!�]ށ>��#��W
ӽE)���ܕY`�0u�Ȕg%���	���R�1Ӭ��9����o�dkRO�u�}�����1�e� �ɷ/'7����!/]u�?���E�%i��:1mr����������ͨ���m�l���;H��ڂ�4��2�r�Z�CN~bv$�Ȕ��BWhA�?6��糜:�-KaKj����ʈ��-��z��(�*��Ղ��υ�1i���(����[s�p_Tai�3qH��l����U����{}�1�o���V+�3��i3�c��yˁ����x�����7�e�PѲ*�؀2�H����"y�n)�sɘ�/N���\�^��U��V�������v�E�?po������w ��jZ҆��ބm�_�g��oPT��c�Q@�#^i�����2�e����	��eB��=�d2٨*�H;������d��&h9:�q%�H�=�kp�j�7am�5��3ǟ&���y�k�k�� �'<�BL��"��ga�q��~%�8�t.��R�09PZ�U,���iޠ�^b��|��K?������kj�m�4Y�W�MeCO�m��8rg,�]*�j�2
� ZW�.4�wh0b��|%�*�|_&+�Qt�%GҬtWbKcib�/27���*�r�r�,tDW�������T�����B�]D��d��>�6�VŅ�����[E���9T|$*E�8�$��/9�lڳE��Ձ��VQ�8{\ ui*�uS�H��u�_�jN��K��ӈ#f�m����,�I���ڤ<8���;����7 t銎)t� T`��7Wkz�
n�U<�	��w�ɹ��?�o���a�N�U%@K^�+.S(����K�������ק̨��6 ������g���|3��"��\YN�&��砞�0�~�0p��&oʅ�`�����ٻ���?v���b}h�G���dSzVGX����/�	`#�7m�Բ���z��aLV����,���;y��*xr�2���{M��c`�� �i�ɭt�8:l�<$��:���.O��������I��%�
5��p�M�h,�Y������^�b�*�U����Y���dR�.�{��K
e_O%��ѡ�GaT�Ƌ:���}�F&�2�3�y�t�r/����2�q���2C�4䮶=]�w'�V�	���T���9_hMI�#B�RWQ�A�ļ��5ŲZ@Z;��O`s�z���ڋvo��Z.�"������3�]��D ��|'�=:�"�������}+?=[c ��KѼ;ݘ`�������$�L�.��������Di[�h/���O���V���h3ɻ�3֮��;�-p�E��"��kH���S���)��%|V(�ے?H����K������<��\�D0sQ�iQm�KH�S�+o�t�i���Q[�⫾YV��������������:F�yV�`,d��`�8�])y�Jo�)��`$�0N�M���Jy�]�B�W���� �3�m�U�	oƀ�n0�M�C�c`�SM��{�q�JW*��<����a�r1p�+,�e���6�!zQ����ˏ�.���3
���ZC��?)��ۣZ�O!:C_�w���9���g]Q��(��8,��	�A{Bs}���m���]�1�W���������!�x5D`[^!��W�ABYջ|¢}�[�(��H�X5��e+H�B�x�в)��F6S��u����<�g�,���(b�솨�u\qa.)��P$t+ε#�Xߍ9�J\y^�{<��u̅CyA~|n��Ti�!h4�4���={���7Y*b�b���:�*�M�+�߳LL���1���+�9��N_��d4#/H��$�X	����
�;�k>�,s��~/�$�U�O��~��7���M����h.1�7%-c�����O�P�fbM�l�@r�������E�	�b��}�нu|ӟ�V���� ����4:0��-�6B��/҄=i�X�O燥�J��QELհ�+�%a�g*��c��<B_W�F�e�=C�*�ޠ�t:�E}���'�@V�����6b�7\$�Ӝ�o�����~�"T ����t���ߒ��$30�t��M��cθ����Oԋ���NN�E���8�#n��՘����+�<.
TO$��,t>_V�Y�g}��0_}�cew��B�5�&� �&��֟�D����y-o�O���)���KB�ߕ����t���\5�^��%�f�-'y$a�E�2��+\飤|�#�{��`齥jeIc�~�TC[oW�rj�i��ƈ	��i�k��-i��g�5T�u�ַ٣GFь��8U�G�p�}��mu}�Fd1�=yn^|������Eh�Z��}�\�L�vvQ �Ro�q��'vc�퉥�7D���Q��hH��+@�&p����(ri]�MW~DJ%5`.|��F<�R�5@�y#	���G �����n��YJ�[��	m�E�@-��O8��] \O����N6�Ci��P"�!���w�P�}E�ڒ�f_&�Q��3؉��0A^_��[�Q`f�FJ4�ned�r��z#��h{J��P_��
����r�'� xiL�
TC�3U\��1׽� ����T�~bNʇ`
b�������!d���� 1[�u�6$�i?�I���x��ce.N;�/��LC�i �b1�B" f v���~:�X5:
�&A�糯���D�9->zZu�p��>�w%n.lf��p�0��5?�|�f�=��i�}�����e()VP���H�����b	'���u{�;��i�(0���{��hݾ��Q-��"�f��mO�6[m(�:��&��:ȓ&L�ٔ���v��x�}zu�nK����u,�5����Pg&�ǧƫg��{�S��)�.`��?�x0�Lwd"�.��R��_��z�WM�[e��$��W��qB���*��7���V�Bł���Q�#���Ѷ���`�x&(~j���Y�nk��w\�6�N��0��@x��W�5-�a�Tgx��Zqg��FL�ʜ/)=E0n�g��+��L��g�K��2zǃ��!E�l��>X}�u&�)}�-��kci ��V\Ǖ\�ϰ��7��\i��lݗ(�x*�9�K��/cI�>\rN�d��28	7�>���K�~jx.s��M�`��x�.:b0I6ލ���S+� ��na+�E��E�˾�.ѫ�Sq-ِy'T;Fm�;0V�����L�8Ho*Gݛ,���B�5,��K)��Fpo���s��p���Kp����Zio �W+_yWl�5�2�
�M��W�l�)T2�ˍX;7:�����24���.�Ex�k�~�z�2�O㿠��~�'w�ʘa��oH�8y�����
;���e=�fl��._�H7�`������	 V$���3cV�G����o��gy�`U�F����*;T[1cH����;� ���+!�ܳ���;�4���p�U}:J�Ҟ�Y����+�L�Y��Vdq�����9o�VB�ऩ8s�Vs<��}�J�J4���74� 6��g.��gf�����a467]����@u�Lt�Mp;�~׮�O�]���P����djJ����䷨�m�o�˭	/Gϰ��:֨�������f��9j����Z�4�t+���u��>�߿/!b\ ��=���Fü�Gvh�Y���O��|f&����#D߄�|ӹJ�$Y����f�Դ��j&oҐ��ouaGsj�sU���/��]?#��b��wN_[���-�^�
i�g��rX;�?ý ���ƿ?;����1i�-�=���}�ӌ�jC���>��`�I��hMCmw�����f���hU+=����Z�!z����TP`�� )�R�#�I��nڋ"���hE�J�����}P���@�/���_�Y��on������
3E��z�O_A���>v�Pe5��52~�e�OZ�Q&�PGb:�@�?}�0�I�V����J�Ol$�_~Ck�'�::8P���tȗ,@d�#䅠�+�]�+{^��*�g$t	yG�HD;VI��������f��������Ϋ`��a�����|x��\�Wٶ��N�����y��^�x2KmTJ��nxM�B~��AXy���k4�}�j��w�L���B�)<&��+
���x��a���UԈ#g�$OJ�;O_ɵ�/�;�X s`�{$Ӌ�)ZmXq�*�8h�ʭ��W�LO�U�y��7�����I]�Ɩ?`�g���8#V[[�Ÿ����!�������e����xX�M�?x�'Ze�4�A�!�>X��{�3+�t/d�6n�,�QvB�����3�'���>;u�x���yR���x��kJ6��kV"~��{�/�݇�!�rk��9]yT�'[��c�w�v㮕�����G�φQ*T{[S�N�"�[�K9]��e#�@������ð~�s.b�c0� 8)�#�%�p��~���PY$�Az�#��9g�� uѳY����)��`Y5C��Lϔ�P��D��;jR�x��1)�C#*>��w+��[�gS��*i��?t�[�HlE����H�P�|�Z��1�Z\c3���U�/U�<�z'��S�嚰�N�o/8�w����GD����Ч�^�b
~&u�{i'!��ݦ�.���u��^2c]�����->�r���[$�8��Y ����J����cW��('�	z��:����o]��B�m"iϰ�n��*�D��O_��L9\`r@V�Q��&����,i���Ȁ�.@�����+@X1��/J��MxK�4���q#VO�T#Ԁ��l�[�/������� ���x�p���R#'���yѕh��a�<�(U�s�n�@\�� �`�̊R��~	(�S�ǘ&je%5�$o�a+�>���O�LL��_W���6��|�M-:��w�'����8Sᒗq_���f���<�,&pF�c4���^���{�h*���-}Q�X\4���I�J6�����HuG�#CsLȸ[Җv���*���i=���U舍�|����V�L34�"�{X��A�r�Nb�3ǟ�`4���Z��$p�[�Y�?7λ84ܿ��+�B�.\ ���/<=�c*��ژD�jl��ܢ<�UQ-r?M׍�L�����i�3^�D,x}��B���5pe��U��΅�>r�B�����`��E8"�2h}͸��rk�|��O4-���/��82.RGԥ���|�!��
o�Zv���й�,D���e��S����?D�X~��!Z$nI�?���F�v��r�`ҚZ�pJ�K=�Lp��K�_�A����N[vy�O�J���S�E�T��H��S�P�*����:�f���V�O�jtëc+��Z�D�Kwt�v�9	3�e��� ̬,�䥋m��;R�!�̄7֠ 5����"ͽ)Dk�\��ӕ�;x��bL,.%��fF���s��@��S�#E�`u�:Xm��&k9�j�j�B�x���N@�E����9�`/lӦ�C��S�c5�(�`<Q�TvgPwx2}"����,�ً��iK��˯�_"��)ƒ�*����'Q��s�t�=0z������L������L��k�A����I+��2�>��F}d2���s[�5�\�_� !�-0��8Id���UKb�ٍt�fj�|-U�^�9#��0dW5��0�N��>SoO�7�h�c�_]Q�6m%}�DN/���(���,F^`��a7�3�+�X��`�k��K�q�y!��]-���`�RX3��� 4�� @��b�-:T��d�Wѯ]�g�<t-��Nxr��5�T9@5M���k��~��=�@�?=N{tF����ɬ���f���Y��3t������x
{w���fԐTt �;��*Đ9i�˹z^ns��)P��3�>�H�{G�B�z�TC������ҿ�D���b@��٨~�$�(B�c���1�P���۳����p�->�����F���,�1鉓N�WTT���31�#�K���Cc�t�"�q�������u��6��DnW	A?�e���,�d6@В2]�ǧ;
K)�B;�����o��c6z��z�i�̸�6�#��4�!�V��u웲���b�W"��Gh� ��1F[����Iq�ت�5N Vt��,�<[%��Fzy{��A Y�%#���ͼ�;��9*Yw�Y������0x��m&=41Y�zz�+.��Pm��`�"�	�(QP����n����D�T���o�e��j�����F�~X�Ś%�O㽒6��e�"���.I��ye ������C��/�Qv���ep�x ׮�O�pη�Q5&��~�<GH��b܅�-pT�U�����I�试�S�P��G�?�����n���=����׀ź\�� ⤇��J
��\r3p��8`CZ1�o�k�R�K#۳�F>�U_n;=3����D��P�%�$",�>�����L��
�T�}w,�`)��҉�V�'�:�9F0(�f�
�mUiK����i��i�����a�g��v2�^�\���r|��P��@ :��oKM��9|��M��X=c���R�B@����:(���h�Ew���N��/������∪���-"��(��c����0�G��V:��ǃՙ��d	�>\�lz%P�B�MU������B�L�2sq2e��+(��Y7bQqKʽ�I]����a��|��*ñ�|'V?��P��dR�6g�[ʫd�7����Ѹ���%T~&j��QғȲ�L]PÐ):G���4���X�y�MH{��{ux�R��&�)�"���oz=��ASJ�Ԙ��ce"�}��B�>���������'c����[r�I�Ey���j�t{vJ߯9%��UL���o�s�W���U��!���P�?�p(��.y�ú���ɘ��`/FQ�C�_94�z�m]XVg��Ҡ�H�itwT7�"/�N���:�LW[���N�\��j�lr� 4^��)�iK]�r��`S�����]��+a���1�A���X�j����
�N>H���>�
�'M������+-h(�~��vl 
�}&j�X�!���7�@�5�H��S`o�٥���G$@=�v�Ș�m]CV٧���
�St`3���z]��R�/��D�Q��]3k�$Z�Pg����;�m��`[R�3�Ө���&��۱cWIM��+j�F��H�\���'��3��~}�TX�K�㸛,%���-'�8k�T��!Q�K�<����xqDjG*ʍ�뎴B%��z`�u�����Y�
������lho��Uc �F���������~b�L*"��K��y�+l�ۆO�������u���cq�tZ�K3�0B���j;�|��"F���^������yRU��e���ňY�U��$}ǰ4��w��Z�$OROan,�����p��_��:I؎U���@��uEy�����C�b�#�l`#S�����1�'�O�[���&n�C��0%��q�@��/IC�*��
POT*'Ti��w��������������+K�n2]oΐ��:}�L��Iy��jY*P̋��L�5�r�y+�u*̠7��U�T {K�i߫��$����f�d1x�����ΠU$��|�/�Z˩�=�,­����gZ�$-�`٘&η֠����e��+Ƈ�WX���+�|VgSw1���������&�r��*#�q���wq+�]b�AM��E-��Ī"�輏MU3�c"�����?{S����5*�t���R���/�05��ϴ1�٬o�+d�	��Z�ډy7�j���F�cT�%LP�V�>P�ŁS��p�PR�����TT�V�H��m�J�J��2�.s�Ay���:��o+֫��~�|/�Փ��� �K��q:���%�d�kݮny��ZAȺ����k�5��h�nc��b�������'ڒ�:�;�!u][}F~�� �n����ì��#���<����B�X��ig2���V{�H `��a��~��/�Ɠ�� U�?�ۖgR�k%C�@>�4�ɑMT}e���l��8��~��Y��2v$ʘ|H
���d	m+���Os�^Oڹ,,�����|]:Za���ɟ�j��p���������ñ�ޥ�&���7�.�K$^ٮ��LƀM���~�MYh� ��=֕(Hי���H�kEk	����]-8�sU��~�N��(|�L����[��J�fC�Y�@�կ�Ѧ�6o��$�/NF,�dx��À@��|��U���^؝�능�S��h;6L'�����w������<r|���	r��ٚR_�$�~�����t�_���ۂt�ĺ�e�Y3Wa<�{�D���Ӫ̧�)�g�r�U���FBT�����d�O��#e�/K��Bs�'�õ.�?>�$c�����%>>��ZyGξ���K1��b4����#�,25]�n7�w�YQK_Kݙ!Y�@L�����\�J0XEJK��I��!����t쒌�''�vc�x��C��S�s���1T�h!�ô�T�%+k�>�6�"�a0T��@����0� �Η�
1�Г��6�����F���
k���Y&��pe�)�
��brHɚ�3bk��Q�;q���JnL�Է��S�r�r���j���Ts���ǨH;{l���k	o�|s���hI���v�@x��v���i�?���96�BҒ���m�<T��==���aF�c��� �h�Ns��D�9��5�9�qZ~0��wܼ���h[sXa��, ��b��޼�}�����x
4�J)�Z.�(����������Y(�G��@fd[��
l�Ci���~D���7T`Z.ؓ��"�����=D����e����&"8���aG:��#X&U>��R�6��Ϗ[0�\d.��A�ع4�ɨ
3c[�2�^�C��b�y������M�̻�{��^qV���Ӄ��g-p0�O�F:�^���HD�k����ҩ�@_���Yp�<�8+�s�f�Y��ܗ�uP�� sp�94&���/�����Q�^v�4��pN�$!Az���<�rȶ�#�!G>D�zX�s��Z(��YF��W�~|���-�k�\�jAt
CP�W����)$���#��-�|t��b��.a��ʔp�9f'��y��m�U�ekZ=o�ifWG���$�P����z����*Xm��{R���B�r�4U����*�G,�'.^�6X��89��QG�ۿ����a�lKq�����J�>�6�~�V��T��m�;���x��DY1x>@8Mk���i�R�ީ�8����v<��.5QU1�ʚ��В���G$��L��D`g*K�^��wV��xR�p����U27���9j�KGD��
�<ĥ�'�Epdn������v`�k��E�_0�����~4�cbgi�r�������3y5eᑺO��`��Ġ�����٨@S_��u�܎NC~�'���W�wl��(dwD�O`�Z�Tv����	�PL ��h�ƳZ�&���Or�z�Ap[M��$F)"."�A��BE�9ϑ�h����I�K!�6a�GJ��]�	G��	7��d�{.1�y����bk>lf�#�I�|�( �7�z�@���=��&Y�4��]]4$^���z�a�s�1α�9��ؤ��]*4-^����;���˽GM�Jn�T�R�&Df9��Ŵ	�������_D��2NZ��Pe��8���Xwp�-֋iȯlԉBz�MDVj-���u�R�׹�)GK{$0%��6s~��N�t12z��*�=�&��7� ���X�h�u8�®Ma۷�?�؞��61/��.��`�am��zqzd��Z����A���3�5<�f��̡]��J$ͥX7&�A��c,*�W��J��9淃Z�ڣ���6�x�T�oŲ7��{�E��4JqW���񧀢�#�F7��g�U�[�03����b7�2g9*W�c�;w�L�vϒ���m:�3�Y����~m���3��7���E�_{" ��ӄa��,�8��Rև)��5��8���U�����<xY&q�ƢW�[��d{KZ[Wq���������j�]f���4)lk��d��)2�C���B�����U$b4��cj||�fuXQg���K��[	�%ƿ������h�a��A���%�ԕ�<�VK�W��p�Eޭ�aE��4R�1��ެ���.�`_ ��p^�� �2#/,�e:ֿQ_�w���W�q��p�ӂ��\����@������X<]�]�QT^m6=f/Ȟ���V���r�9,�R?lտ�G��r�<�x=��ҝ=�An��k<��g������I�A�&�@h��15/=T2H*���rfh�@i�Q�WrבR���~�#���O-V��A@;V�5N��v���/���YX}����/�x����7@�\6g���=�"eS�Y	��^[���~P@��~ 8?�自��Ļo�ӉM���>�Zn�7}/�؃A��8��Y�G7�� \�%�7�(�H�9F�\Se���2�'�Ґ�M�o���]h���9���]��]��+��6-bv1�+���˔�,��t/�(�k	HUo���:sf_��@�"�E<�q
{�C�7�� Z�{%�흺G�$9�H��I��]�j�g�>g�'f��&��ׅh��j��~+�+f����	��ׄŘr���|�+Qh7���7���F��/��232��l�:�Nn���D=��0Q��ګm����$��xz���<���24C��e��o�O.���<x�z��j�i��!;[Ɗ��NE#��H��y�ɵ����1���5YEf����$a��2��}��7�"�ܸ+��<�wݫ�LL����`,_Ն�]z�ӏ���*�7K�p����Ѭ}�"��V��ҤW�m�4TP��+�F�����?��$��v	�F/��_��1.���� 3&�J���T�²X&�'S��G�TcwtGp��S4��#BP��>��D,�o桇��k���%���<���J�?�뷪���鑲OB�PX˓7�)P�T�}��=0�3A`^sݓ~�X�Q�碦wG�Y��kJv4#�7�^K��=��#˘���R���zZ1EۢW����,�Y��,r
� T0j>�ZzԘ��-(����n��E�($&�v���d��-��㻿��� ߕ��{@^OX�&YTo.�#Rۘ�RCx���!��zp�0�`�&HE��\�3uF�σ����e�Xf$��YN�A0�G�c�>-�4���l���*����/�*mY��[w�"�p��;��M�2#�"�;��d�2e��(��b���
�ׯϱ� �M0��S?SG�� R\��6�bF�����6�j u=g�:.B�u���7!���r�!F¯3@j"ん}�dL`��X�󿸳��B�^h�z[����A�x�<�|Jx��āH3K&�'1��~p�m��-Y�J�\�< g�FlN���еO�{�{m���^|�RE��_����I��W�u/���M�:���΀��2�����@�0�H$e����}A&���k+�0_����}Z�_�!vm����b��<��&��g���F#��)�#�w��,���ai�|�R���uV+A-Q�^�َ�����B9a�t(�����Ff`�AQ�ϭv�Ѕ��b^`����a��˪.��(�����[渕����Ʋ�f���0��4i(W5�|��.����ϐ�h��@��h[p��'ػ�M�b��F��O�TC���[�6ss�a�I<�bg��hH�H�l���K�����:Y�H�˭^w��vO�'0��b�j��r����� 9�J�(�b�xR

t.%Ja�$�д�s�w��7���x�;ó���ފf�5>�=!�ﯗ2�<���RU���"�SM������&Ι{��n���/�#����
��x��������c\��/���7��	�g%�����8co1�RCN.r1	���T�����~:�{V��
��}6���5ޚSǵj?�B� �^�p~�Lو���!<������d^��������Y}���fd����S��K)�\ԛ;ܐ/+��` MF2%KWz�\#n�p3��xKP���^1�G��'�pt�%���@�Q<��?I�|��� Ϛh��N�5^��O�yB{�0�
;䊋ǈ*/Z���Uz��aC4!WA�7�395��V�����j4�Ť�� �T��1�[�3�0&��"i߰Ý9��Z�d ��T?A���}�n�>g�z�8��ƚ�=�P�+J���]�Q�l\Q	��%v��ZM�QX=̪���
�~;a��L�yK�N_��k�}nJ��'����U�b�_���JF몥t��F�8l�>�y�~!@�%@�ɇ˅��ט-c��`������At���e�����@��]���OgNrx�=�MH�yF	p&�����e�1V������n�F����9#�2QId��F��g�mSU.�/�8ma���Y��w����j_7�Y+re�ή7�/ٳ�|�]M��-âkE9�Sa`���b73Ek	�!2<�%�.�@ɔ#�r��)_%;P���]�DύTY��[��ׅgxC����b����6X���^+�์F�5��c�|�1�oQ^+A��3W�)nid�Ve���(PĘ��CH��`͇_r�,���@�ޭ�<�!%���N'Y��jN��2v)�7�AT0"�_��=�>�C%���Bz�����Q(A���n�Y����h�H��i-:�3F[�y���S�%%�G��0T���qq�xl k��#�u��D�)Ap�;��㥨n��R��@���~��XB�g���,N���0����o��)��\�����y������Y�!���f�Q[���ܼ��1�TaKGԔ�y$��I������8W��o��/�b^>��f��lT2�g|���0B^�b�3 D����L06��ڻ��'��}���>��l�van����=��EeTQf�q3_&L{�n�D�f�
sKTp��p�j��jI���Յ�J������03�3�D�
�U
���㊨�<��<�r����~n���
4��������ތ��a�tl4eW�zX����btg��6����(g�
"eO��z�d.<͇W2���ZT�xs����oS�{�D�c_Q%��?�t�4���"�r�yV˳&֗�;4�Q�K&V!YU5o���߾(W��~�V���x����d��`r�B���!�]]���r���l~l-���z��@����/�RX��km�1������Z�3�o�ћÍM�Bc�+t��ߡ��	�[�<��*#�oۓţ#��~�w=Q���f!5>�%�y�� ������9���M��p���{�<�<`�I��o��+���T�\��Y��l>$��D�jF:��Z�j���NJ�-�#'�ʀ�P	E��@����*���P�u���o�'
X��6�T`�M���Z{+dFu���?�R��� �hu�s���I�Bsܸ��I'&��cK��ʓb��`y���J� �ؘ�� F�Z���B�xyf�2O�NF�M�݅������Gk0p���R�z���c��(��k%�1YZ@�]�<�!
� ���1����"��],�j
?d��fRB���G�	�1)s��=I��Tϛ�s��m�I��o�^D�G$�Ad�&����^_�SE+[.�E������Z�T떙��,ŷ_����LO�jo�$?����y�,���,i�uk�M!#�8@��($������#9��J��y~ʟ�*��A�7lD��4:��6��>UV���+LsV󧂂�T�.ݭ�i�=	m���{���v[���}�o��lWE����]��f��JuV����Zd�������+C��;����pu���45�nx�ȟ�B�`��i�!�͞��n��I̥JL�;�����νQU@��!8��9[�J1��~�<��������n�2h#�r�fp)l�>?R<Ѫf;�˹�-���LMxt� O�@������0��hIn.�4Ƃ�@���K�;~k�$�iޘ�����ɩ(����|)-�ܓ/�i	�N��fx��Η�Q ���1*7M�]{3��A��Se\6���-��р=<��5$Ǫk�Nv�F�X>9v�[�k��D���'�KT]� �·�m�ڴ���=E�"��/A�q�O�8����G_�j��:�@-�B�onV�����y �U��tR� o�Xս��a�%d$�Uz ��b]��{1(^=Q~� ���{�)�"F�C�l�A�ȣu���q�;��Q]��P�cN��.����:���t�ؐ�;�ο0B�����+$�g��J��Q�tsĴ���a�%4��<� 0u�|���6���"��x�Nf�#��O݀�VޯIk��H.��9�s̶όŤzX����,�߱g��~�y*���h��g +�oo'	�;UD���[���& ��{�3���^8lX�ן�}�.�#�͞��b����870����W�1�7�0ZCC9��n��O4D��������-�?���Py�=L���1�\���}�V��
��ѝޮ{X5�R�k��|��1L�I�1��U����p@��_+�O�l ��֠��
)�m�6��\!�0�?ܵ]�<���+���5�˪	�,p�u�'(�B������.K�Ja1�C��
��:�=���mB�'_��&TuHvGr��H�]����f�5�Ȟ[����w�-I�Cr���Q+�Nïc/2�=��Fep_*��'���R���Z?��8�Q��L���]�
.���^żr���ƴ7G�J	[2�2Z��$y���_�d�s����tEk�%b�f˖+�. �?�q��ƕ���-�����J�\���IM߃�����ǭn��˸�5�� 7��lrDl�*o�TJ9q���	�	�#���[K�?'׀^�k.o��)|;�[�i��c��N��"��ieZ�)#��G,A���{C�&�l㪎�4�"4�l3��a��D;-�ɾ���ctbᛊ l��x�3d��RLk6*�#≯{ÖD��52�3��k��:H�T�Wt�9j*>����"�L�J��pFlAvFN6>�pq�J��8��X�$Ӹ�X��=���a�MO��H1[%�z�	�<�k2  �^���x��B�Ɖ�Dj4�lQ�_ω�3�I,�^��q�7/���v���͓C�/�,�H?e�\u�Kդ%��g�7�A��$κ��Ϛ>��'ミe�����ҵ��2�V������B�AU���o��l9]I' �#j���~�h�#z��\|����K�**Ͱf=����3��Y�J0ڔe���/�kK�k�m�w��D��i��ZZL�?҃���!�l�n.A7r�;6p��o�Sq	-����u䖜�,vᦴM����`�-ê�1��ZC�f�ݍ�]g��n��y�%X����x�c�+��t ��I�H�g:�kD�ϗ����:#�~�q9?�e�	O�+��T����V�i#`?�D�s����YO��v{��R�'^���[~EB�z�W}{=��Xυ�=��e �쪅�h��,,�s��ˡk}ͤ^r�
å~K0��Ƭ��2H��ϩ @.^��Ѯ���T�1�m<ّ�8�|o͘1.|Ub�Ե�%��S�L����4푇Z�}������:�
<%y�� ��@��em�M�Y�'S|H������	��.�Q	ҷ��1Y|�}d�-������gr���֙��m��ׂ<��t>��ISpը������&P���3�)�$��s�{�rxlt���pb�^���hY�z*E�^[�$a<�̕s���|
*Þ���ɜs�ըi��b ��M	��X7H�Uv.s�Q/��I�s�&o?�׸݈���$����zS�]2�>f��D�}Q�G���q���(�~��@�
�%R:W��|�+��tp�g�q/$����oM!�۽Z�g�z�d!�28	Qz.֮�I��d�>*�m�����v2K���r�j�x�º��tp��*�8 ��Z�4�B��*�������&JaֿsD�+�݉ӟ��w�"pߝ����jM�H^<�X3�AV8�xtu���@�'����K0hvz��ڳ�j��&�X������Xnw�=�ټ]i��/�E<�B��]O�WѸz�e 5F^{�q�i���R����u�hw�E�n��x��t�
�&����SY�)V�A����g�&�=���n��	_^Wr��X簪�F'Վ[?y|�B�E���C�0®y�'	b�Lo�������n�Q������T
.���:�-CP�`[-��Α ��e��lɲ�"���������Z?K��[�.r5�ե6�p�i=R���%��s���[�&ڽ�����t!���ևV���ߐ�.��5����7�g��~Zo��ݨd���,��鞒�S��!��(�2>|�_��9+J�N�g�X����.gw�&*�xW[7�}�hv:�[����,}�b34x��e���+�����mЋ����e�֟�j����iDXs(xۼ�6`��Qf�<H�׏��"�t�&�	(��/<Y��8�B^f������05�������-�U
�f�o�1%N���>W����Y`BR��x�����I�0�����(��P}�&��Ds��y��#B��7�{ʾh�s
JO���9��|�"*�U��j-��=GY˂-I[�t��8�$�����0"��O�a$����
1��V���I+���]��/�n��Q�m�+Te�N��7n�4
a��x��Lf��I�e	�+~�X�5;�G\�<*��X2^S�Fյ^�|G����f�P
��]��=\r�f�@��W�/��\d_�!~���^N�i�$�����R�_��9Z�^ɘ���.���5t[����x�����d��5llG�c�+2�d��4�K��i07�udV�T�����E��Ě�ܪ��g�
�?C7�
��7�����7����u�}�,�YK&��J@)(��Ŝ��vL����f������=1X/(iV��+Xq�{Ls	�zy�(L}U�<���(�<�E��c��q�.49䝿�/��x�=`'l�ΕX�5M�j"�P����h��FP�r!
���-1:�d1nTQ�`����"5\=1zΦ�����U ��a�,	e�D�m#E�B��X�â�D�$i��r�e�*

�eFO%b��/�Ǡ��2B���h3>c�e)�xfZ:�������ut�߮fi�{6bZ��f�8�F���j���2�r�[�c�!�@&TT�-x�LAP��^��b�g�2K�� ��H�M���QX��ua�ꯎ0��~�\7�8*�PD�@;�|�l�w2�@׮!�ҩL�{��?�I�t3�{�T�Q��4�C���oK��lxV�~�\tv>�g
���ڛ �}f�
�iZ�-]��ʬ�q�+�G�h&ĞsƝ-s&x����x=m��E�P�3�ĕ�ǧ��@��
��6�8�{�u�ߠ�
�9��Mp^����e���U�b�?5���d������Sp&�^�f��z���yi��=�|�:�,�� �pZ�/^�%GK`��r���xt%(%�Bx�
�	���|���!�_���7J�Q]?�?��$��ۡ1�����ALq�$���=i��~��n��Ysu��z�j?��ĐmN�qY9�ҍ��p�������&uᕼt�e��Iu4(�%	�gY-A�G���0��/�f�*�3�?6����G`y-��W�I�۹�@y����&۟)n|��f���Ţ��G �?6,��i�1"��L:D�H� G�r��b�fJ�P�j����Cl� �w�����Q�h#��d.Qk����U��$*ef�����ƒ�F�JER�u�~w�*{+V"���u[X�>�s��U��OA��G���7���<3����k{c�Y�Y�65��C�0]�:R�oBr4�D'߰!�_���K�D޾�pÓ[J�/zd�f�����^��Y�Y�V���#U蝮�k��H�
I�T�����G-���"Lн��)s�Ŧ&�*�:x(v1�>8&8��\~z!j�R�n��I(��<k����1�*�T���@,��X��c�{Qn����?@�]M�CNfl�2^�&(�P�N!�'~V���G��jjR-
-�ژ�=e,�B����������A�7U �8K�_�O�	-�o!����p#%ɪ�M>�"��C�눗knvS��06��~�9f r��\���5>=s���ɤv)B?���u�Tp�� 7���NǛ <�m�&������#٥�	�ug�(F�z;~w>,��tɍg;p.D�%K��sZ��mPL����[N�ٸ�Q��C�]�u�h��e���>eU��F2�z��7[�o�]�w�s؇5���7P��6�gRٞ���8�BT9g��5���G/��9[�Ç�[�oWT��-�ܮ-�k ����HrU�{���U�ks[���܋U��	��4~�߰+�����;�J�<�g�4{��Eb�s}�.~�<��@������j��l�1����aK���{q�#y���h�^�ę�@�:��ۺ�r��k��@J�c��5���9H�9q	D�y瑱���	=�Of�4#�;�0��'� %��ԨT�Ro%xB��A܈2Ѵ�
��E�AoЈ�rHѨɮ�2��p|�f��H�3��?���%"�X{{3�����;U�{I�J;�~g:p�v}P�t���Ep.)88wU���{����|��1D,$�0~�Ƚ����Uܭ@�9���s>����|��G���9�x��^k���}3p��
3Qf_�����S����"!��[W^E��ܕ#XaZ�P����6�lF�l�}H?�v4B�4��Q sC�n�J�V��m�����R��,A"t�5$�$�+.��*Mw�񗟇Vϖ��t`VϖM^8��1��z���D��7���-<�[Sp���ǁ�09��^@�b �VQ����:����ӱhB���*]��5u��K��'�$eJ�ȵ"�W�P�k֕Ժ�y1�]��0�7��&G̡���Z�B�;���96Nc��!ԏG��7�4O؃/�
S�}&��>5�	'�g;7_,%+�~#p`���1����Y���=�Z\@Q��g�qH��	5>eZk�� M���D�暨2�u���wy6R=Wn(#~�>�`�є���^m���z��:i
��,6�-o�>���FXw��?\wp����Ɗ�����E�J�`��=���.uЋ�.�ًv.W���z�v���F��b6�)��g�(�#7�>�d�ΐ�Y���>r�aid��b�v����M���H��ѶA�Ұn���)΀��M���屔:��-~[�`��B�ވv��N�	���O��'�4�`�d�z��v�؜�@+y��&G���)��U�]� 9*M�ʎdOGg,(I��]ܼ��K�Kb�����p��˪e�E�p]S���(n� D5K1c	���wSӧ(S.?���=�3v[���_�ݦ�.����.횁v����ۋ۾�j�fWw6�y����$��Q�u,�"�_@�m(�5`If�19��������+?~N>SIE���	�,Ջ�t��@o0��_�|�u^vPYްL2���}�Y�;v�C�ĞV�����rxM?�
��|S���K�OaS.������|q�YB�c� �(�}Wao��_��f�#�;W���st�#.NeA�~�2/�g��AB�,@��>�-�����g�'?8@�H�o�ǋk�PלhA_#4QIE�M�2Vu��o�u�2���r.q	q�}��y��������?HW�w{H�����8�4<�K
�+2��ZY�����&^�O���4�L/]aNxc��+]�0Ѭ��f�Bd�p��x͹O��2��Ԙ���!c���O��yǷ��$�D��ڋt<��qJin@ԅ/�����n��!4��p��Ͽ�-�����C��C�� ���g\L8#�*	�%���oG��P��R�z�� &=7��6�L2�_���HrY�&ș\�k���b1�d���������/TAdMc��-����g������� ��k�߬���ZT\��4�Q�z���%�q�J22�]��Y)�N�$���mL�!�5����.pЇ�#l�6sҏY�m�X�`ܒ�������RԤ�_���gw��Ǜ,�����V��
=�t��1j�k=A}��g�Ȁ�4
~���_�o�}�)�����q�r�Ph��a��!������ ��ֳ��>5��mQݻ�Q��TV�{v�������M���Ŕe��S�q�����g-���)v�
G�b"8��O�R�1K�!8W��~��7yd��5��*뙻n��HL�v�h���Ah�;X���2"T�D��7��c��W<��[v>;(�]�]�V�, �C� ��[���e�Cl׉�z�Qp��y[8��p.��Ҏ=�^�'.�(�Q�p]��or��<��$	4�=��>� ��{��	���N��gt:m�KD(���.Q�/�����XP�m������ɱ3?�*�!u��w�#�oa�o��ɑk��l��5��)�i�0�7��H��s�;�P�R�UC�����T�/򎬹@�Ϧur��Ec��6c�����ب�!
/���:T��ؙ	(�QW�R�&���� b��뫓���Y�1UIor�����D>��R��=Ϡ��Ul�ew�?�0g��x�~:����b�ow��Yjʅ����CꝆW�:��vɨi�]���'.��϶��EX�F;�qI,�p/�����0��Zz&1@��O`c�;�f���:�\"�a�.儆{
�G��Z�{����
�~_e�ّ	��ҍ8| �1���h�>y�6y�bUI��fՀp��g�b�N,G3��4�]�;Y��E� Zh�[�������NA>d��u��3�/Y���8�Q*I�=Ƒ�?#ͤP��I-�d�
w�#��	u��S���Z���qNʥ�O���B�̲�l-�£��n0�ԏ�!��=ï�h��}�g�kb��I�t��(�s@��_ a�P��^ԧo�����4ճ2�AO! ��M!�����-Pc��NGБ����4��G�i�`��">��6�R�SM(�O�%���ևI����PBj6���j�������¬ �� �����X���Q�kݬ��E�B$
; O�a.���f/+�O]ŀ�Al�e+}�6I;��HugΜ�18�a [�dϨ�R�)�cNQ����*�F�Z���o�G�泩�BnR���O#����!�����
Ǧ)wk�^Q�l}i.�%�	����g��e)VB�ଢ଼~]�6�"ʶ�1]F��i;v*�-R������E���U��G6�ƊT��ڗH��ӟ��Q#4���P�߿�,,��;FC���jg��SX��zF<�=!��B587� f��t���=�{g)�������B3!��j@RK2F���u5c
��QU�i�
�[4�ׄ��|�/TO1���fs�2��]�|�fh��,�$t��j��U��H��W"L9��m侐y=!��dk�l\B�����d4`xô���B�8]_�cs������(���}Φ�@ �O���*Y�����;�V-fj���M0?�3&���c^��{ɍ5.���F��e�����^yn�-	>��J��<�y����q����V���PL������>i*3U<�DG��*LA+eA���_��vh_�ƥb��|�y�=8lOb�@w�_<�S2eI&��g��A����O{i��)�k��ҁ�M��&�J�p��F��V�G�` n�'���5v��ͬ1���Nl�c?ן8�_-"7狺�'պ�p�{�D�(�uPƴ
I�@�uL�ZgBJ�%���߆8�h��c�DI^ıf|��i�Q���G��[�]K��UN1�8�����0���{��q�bk���1`%4Đ� �H�L��o�g�$�/�<0�ŭ#��Nά�μ���4�}A�>Cd�0փ���0	h��g[U�P�����ǚ��>��|�t�Ҏte�rXF�F:�������yC��h%[�u���/��֑y*ŵ�N�"Dl��S�l��X�����[q����!�~~��= ��!&�-�+<��ww��)��n4��Oy��Z+"�An�Y �1�.����$� �k?�Y�o#dhB���Y.��gT��w��I�D@t`]{k��h!.-����!���|l�>�[��ݳT�r�=�N�H���8{\/���X�T�T$FB����,l�/Ǐ1��tY\�����P����;� ���9��ɐZ>�c�9�~�!h�IB�]]����-�5	6aK~ ���|C~> y�1��e�Z�.cpr$�@�$Hl�(w妦�Ͻ�
���;d`���4�L
�n*���)+�ioHC�M��I�X��΢#�tƘ��Z�����WMrk���}�G���(�EyeB���m��mòG� ��#�j��ܼ�(���)F��^��`�$6S!�����ֳMo��ۜ�kp52�x%�}3��@?�/��O����m{����5�nv^��!p�>
�o��շ1���H��9� N�xYT�0	��βG��͐7�40��R���,��]��)�e$��-Oߕ/���U�`�l<�Z;3�s�M��F�l���NG������� �ؑ*KN�Ԡ�D�s����޶��C�>��a�\ݘ]��!�%?�W���w���RD&�Z!�(�:/�I��1��9��f��4)����!�X|O�V:(I��gp��gdm&d�R�e�pR^VQ����,�x{�ix������5��~4�Q �Tpź�ˎ�ȹݡa�f��={|>�~�݀���{�����=)-�I�L9��a�7Ы�֒acj��_�y�9��Z7������X<qPs�AL�I_���8/�{��ɇ#H��J�I�U�d���	�8__M��0�D����OKa����a/�o����D�^޷L6�_��(L��P�p,X9�W�ŵs�l��n����es�:�	MB"ZjJ�S�4�Œ��ö�)~ɽ�p_��D␆v	^�ܭ�}���v�?�j�U�����`e�(�1�t_���(WBt�����j^tKW#�/~���;�9옃b֥��c����s��}���T�ʎ��mo+w�]�_�ƬJh�9��8b'�ۙܮx�*���ŖV�e;�nX�#F��6��wer��xW?�o�0hk>�jj8��sF���}Dڪ�<6�0�Ea�� �QU��D�ur�����D�h�&Đ�xn�*GSa��jgo�&�[��W���Nsm�
uH	�ô�C���0qAilA�1�M��j��d���U��5�R�X�b�S�
�8]y����(j�
S�_���v�,��%k�܉���d���ȵ��X�J��3�}R�9�ʓ�JrB��Q6���(Ze�ܹ(�P�kG��}������& ���'�4�L������GM�_����Q����s���Z%�(=�����Ӕ�ԊOn��`.U{�jB)1sm��<9�������1��4���}ؾ���:�|�&���S\�@�6VP[M�!�.j�������8AOʜq��0x�N<K�[Em�@�$)��A��ar�Ն�����zx�Yʭ,�� �z@ks�/B�Ǫ/�8���V3�k��`&�<����RѲ��
ƶژ Z��9_���ev�j�&�v���� �������/A�g���N�&�Dc��$�3��:�^`����aM�t�%���R�2��{#��1��[pAf�52����t<�c��+t������]Y��P���pC��Z@��Uo���=��Ǒ_eiYu����IA�����A�J��p��z{�Y��2;��A*����쾗z%�u���r�ӏ������]�o���U�e8 �O�{U�Fk�i�!A^+����LK8�a��R\{e�$��Ǽ|�4��1[��]���W�븮]�^W�$�9�m��5*^ꏆ]12��Yp��d4/.�Tl�Ć��ˌ���$����2���¼�4�1-N��M���:� �::A��c&zpP�,*l����5���9�E�k�"���!�1d�T�мpH��6\�v��f;����
�m�o�1Pʬ�q�4�|Gn6���SPT��E^X=	�X��ժw��7��2g�����fMAG���@G�@U}�wcL�5Pt���������.�h
���� �#j>G�#Ge��]3�o�����X��jq��(�7�zqԈ?�5_oVU���+h�pC�C�aGGW~W00�ƽ��H+d��䂸°	���sxb�Xn�e��K�zHs�"2IH��N����zD�j D(P`C��v��y�(��kC���Xn�}b�^M];���9���F��#�{� ���2��M�`�hC�6o�]'-\��mN��8��������97��첧o���C�{Jog�1�?��H5���8����S�7�K�J�b��b�����Ԯ�����sU���Pf_W��$�:*`���Y�%�g��MK�3@rfs�Y .x��'�%���86lٓL�|pd�+�.�bu�NU�aD;���V`��>�Aw�K�R
�ש�3�=v�L�֘��V���[�e��{I�f}u��KYh�z����!eF��GX�G�*��0ԽѠ�Վ�l�X#�xҵ�w���Ǟv]���sxMn݋Ki�_��D��5��d�����A�Q���?k�`o�Y;��e�#�*y����Onw0��k+�M��`��y�$XrF�@sݩ��:U�� �!w�0�%���
�
/��%�6B)�^�@�?_������X��O���ed�GG�����*��Ʊ3���`�XrKW; ��,��E��j�������N7�-5��0�i�R4ۏ��Cs<Dܞb��h��ܻ���op]*��>�h�{�sA�d,���a�$xe!��fڃҨ�k���y��<���\$Ykf�'�c�����X�ЂY��Q�H(N���%�P/b�Λ�����{�:W ���ڇr8�󞾒�2z�b���E<�1���ׯ�� |�.O$/�>�+��S+�]����ɦY�?٘�j�n��.�h�_�-��#��ٳ~0�$}�&gF�Yw@�4y��2
x�g�!�r��4r�%�ڙ1\f'�����N~�� 7�]�%��Nș�Ş2�(�S�K��h|�qv`�����gQ��G����e�h:�A���ܼt*7�`�{�U��8C�Gf�k/�v8F��yaHu>�������4����r����H�O�a�pJ�`N������]'I�b�z��i��Mu�n��GE�D��#�X;+�d%�RKOc��[m/�L&�BZ�R���t�E
:5�X���������mz�d�]��G{3�F3o������KF�ӈr,�,'��#:ʎI�tb ��D؉�~��?�m��=��ڡ�%P����C�;�}le�-�t���BXNh��-��&F!UR!�{���aH�Ӭ[��8�Z�l��G��&�c%���Hk�����B¥��p�����ɦ�f}�N�鍎{2c��9F?$'O��P'D ��x�%���-�h��m�I�E�����j�|Սld����/�Z��8b���Ty;��9y�͝��V���q�w���j���0�ɐ�I���������R�ye�~�=�� �B�#��7�����d(g�3f
�k�Sx��7��q���r��zM�1,���d�ɋ��d�15�*��-�Mo������L�*Bo�Ю�ة��rʑ���/��B�-#��3Àx��9�Wh۫~�#��(%��?qg��@��
vtr߃��:��[�>l}1���Ue���a���*��	�ն�:b��b0}�Ն΍�To�݊���@6��_�֗��x>A
�����n�tſWUR���/��SV��<Ac히k��X(c����\d���A���!Һ��滦���j�j��d {@�n9	F����ڿ��x����y;���>���Mq��J�YE��c�t�aC� }\�e~T�9�lm�����ײ�������������- ����09���<e���"Ǹ#b���@��胟~H�m�-���-��!�M���ⰷpԁ�,S��1��X"q��ι�P�[�Ԡ�O�m��*ي$x��v��s��q����SǢ9�A �W#����C�}���+]lv3Wo1V�m ����!�S8\��b{G�yrpg��
�o�=��<X�,]��
�y�V�N��{�W�j�����_qJ_K����e�҉i"z.0Z	$Q2b�IUP��l�*i�T��7L��؇��w�VK?� �R�=�6�*�rE�r�z�'|���N�=�; �� ����Ŏ���Im�e���	�O���O�1���:b*��5���:L��"�.�M <�٫ޔ�3�tː�9@j#����{1��������%����,�����/KY�r�#�h�K�׋rI�lB[d��$p׺��N�nߌ^����z�]���W�pЬ�g���=�����z�@��NJ�o���ˢw��^@9=Ne�Cu���k���oM$��Q�;)�sآ�!wC�mp��R��σ
[� ���h��S@ r��,�-6�n]�i ��d����@�{A%�4G�����K�Ot&ЕLˌ4����oa��
&$�+���K�Ym�2'��9T2��Z��y���#��t5�H3��35���ԉt�'@4�0�揅����P�K�Z���Mr��%�þ>5R�#ԓ���N���Z�NaE��Ʋ�v��y�<�I��9�=?�����Q�?!�L��)�6.�~�;x�c�V���R]n��HX7�LG���g�Tɳ�䂑C��������"J���ws��{���Z���� �ad���t�s��?S�Q@�!˫sh4 ��i٩)�i�J�����z������8)6�z���2p�߃�l��m9h\:��:�(��	IQp��ږ��ψI������a�H�?E@ބ�jV��1Z�Fh�vF]����#�j�5U|,�:3�l|Lq�,�l����B�a�gO���]��|N-��WO"�
r-���DΪ4h�4�d^�KΆ��@��˽iºؔ�8�zÅc�D�k^,<n�K.�^��pX��q/�Ŷ��J>��]ʚ�2G`��Q�Y����8t���0���5���Đ��:;=��{�2,�ȓ�ud��B�Hy�l���ʓ�J�C��d���C>�W5�[�u���]F]�����G��tߣ)����`�f�ێ��[l�OWٙ��@Ri~V73d��׭'߸�bH�iƩ�g0���Q�`��2�e��M�����J;����kv�����F V����KeD#�A�Q� F ���˾ �ZaL9_A�}�����!ڠ��XW.h�S��4��?i��~1#b��B��uY\�k���-�7�G.K뺔 ��Aa�MqD���ѻ� ��bU����P����Tx���+�ֺ�����G@�d��^���nٰٗը]�?���ҟDuk�\L~��k�۹����	
�/V�W[��O��v<���3YV����S�����StWo���G��� � n�����N�آ�eL!����|?��wI�d��l��Y��˽��E���&&�g:.Ϫ ��۸���s������cA�[�������t�����J1��#�(����Ա�ߗ-q�k@�p�g���c!I�?[�P�	2�<3%JJmM�Wy鈤+>ɭ�-�s��c��A9ǐ�}��x���A��U>����U
���Z��[��l�.Cxv�z������h�%�?e���_.��G��	<��s��A���5D��׵����$�������p�&s��p�>?b�\��wh%5t��`߽�ڣ�aW�g	�������5
�}���1M[�^:��׾��1{��O'-H\��Ɇq�R?���Z��3�O�Y0m��$)�Jj��X��%Y��
�����7��oRu H#R��NQ���G�/�rc��v]ؕ�'� L��R ��_ʹ��z�.]�\r��p>���F=��z�w�4(�!y� 
޺�g1,]I|��/�W�� .��kt��ޅ����l����6����ٟ��������F�K	 9Cs����l"�+I×�*h�0��V?QpY���PXw�{��X%[|~�!��6���x����j-k���BRv��ș���I-Շ��;�	��A~h)|l��&@(���}a_r�ÈK�\"�9���QC���T����Ok��P���d|n-�p�d��>FzHf���>���f"D�=T�Rya�m�E[*�/���)~�N"�ܗe8[���[#|P��N��|\I)ͳ-���h��ьoL��1�����K6��i�M09�n5���V9��.�.}�gi�������/���UK��1g�4�#���}2����jR=^�9ǣ��D�o�5�[�b�4����]F�SH��l���|%��K{֏�����=f�,�&9@�����J�w�Ž�5_N*�0�noub��g��] 6U�!�PAx����5���4&x�xl��О���̼u)g�lI#�ZD����q�1���s��M-�$r>���\��\滍��'�s��z����lxH�^i�bb�t{zO�g�6ۣ����ġ��ߴ8�ty]L���io�G"&?�T!�GX���Z��Wug]L����@.f���IH!6^eA��J�C�����u�L�Գӄ�;9�D[5��VP؁�B���<t7�z����xe���m�E��{���ͫc�p/�[� R�aB��c9�����q֍���z(�;�W������b/SW���&I�8�i"Oc7�]q�����zTy��U�	(/���w��s���ݓ�N�C�C��,���ǒZ�j����~����"�*���y���^��(�?~�����3�sTm�k'�T�UA]����O �0��j�wY�m�ɍ!�.ݲ��`� ��8Q��O�D�d�z������L(g:^�>��C��bM�3p����"��!
���
�\94����k��yuܬ!:{�_Iy)R�#��&�ts�~��%�[���@z5�{Ql|}�OA9@��z������=��d���r���X�x�������Um���̖�4��n�;/�G�#5��z|k18'�g�C��q���2�|q����(�h"�uF�����G��N��pކ�z&�=њĈ�v�L��J�BcĈ��!�Z��Qe�kP*0鼕�9R����L�n�H/Ssp��>G�Hc!3�! Y��B�M"{�ʤ���O6Hߚ��Hx�wB'W��R��}rL$u�$��OW����wX��Oemu�Npڀ
�!������菖�+�4�K8�2���|�Ԟ%(0������m'�US��[t ��3�\Wk^�|�ţl�1jEj]Q�`0D�������4��u�$�F�3�}JF@H"ˣ�q��*��)_a^��#����۹:�b���u��L����B����.�����N���+�&Ť�)��i	�J�Pux� SL�)����p9����`��SX��szB?Jy鋋�<��%����M���Ε�Z���I�kX�%<�&�v���4H�=���р���~�G�\y��:uQ��r������'�nI�n�at�vLD�˧��'Q�T� �F��0#�:0���^�Oyb_������t�!�W�'.i.]����v���-�7uU��L�|O�y9�^S3�^ �&�����`Grq^���3����!e�G��� G �(�bN���?֊g���K��é(_�y��7��Z!��'E�<�$;@��V��Y�!H��:	�J�5��S>�\�n�G�����޸�0	t�K�<����S�8Y�#�I\
�m%Ҋ
�u]��}���qo��Kȴ]�7��#"ή��Lq����^�\3[���(�JRc��G��4C *�SH��_����w83���:��9 ���ͦ�E��ǲ��{N�ޤ�SJ�To&�_���X��� 짳ߨy�����/����$8���=���A�9�r������8c�1۠�>�N���L�Q#��z�m��U}?��-w�{	+>��淫��,*��S�,ؾ<����1�l��]�-�ٺR������3�cz�P�F���c(]��h�'��Sb���\�b��m�rTM���P���-L�g��X�E����}�r�h�H�{[sY\���,�X�k��)KO�}"Hߴ��^$�Z�\g����xDo�]p��F�'����n������ce�J�%����4�<b��Ʃ�Rs��Ǥ--:���L��C������m�(}My-h��v�o��zɺפW�^]�B0��\ff�3jQ�9�LR�'�â~�wuɰ�Wj���)y4KV�&V�	_]p�:~�ʡ��r�E`����ӎE,-�*��T�d֏�Xk-��rfL�$ xX�ō�^�5 ��1�)�������&� a\{��=���X� ��s��r��j�>Q��oX�("n�Gz�\6
�w��ڒ�Ps3�\����|�a�e�)�5X�����N��q%�X�ھC�����Avq�(�Ժ����GO��B95b_��D���}�Z�0�J��<^/�����bmuqN�r�PՒ��9�}���9�V,���݁�'XJ:?h�� i�]��c��E)����!�F����w�{ـo�e�[8�iÓ�љ����������a|T%�� ��[Iv��V�������k�a ��%�dO��j��/�Xs�tB��*Q�ː��I����Kx��]�;D!qT���ȹ!�"��;st�q ��F�jK�����,���!����gݡ}��RS��d�!W��f�Կ|M~D��/Q�=�u)�X�V�����Y��^���t!�M~TY�S��^_w˘T��)��"��U����y]�P=���$܄}[�Ee+�[L����7!j��,d�Y�ք���{�a_l>��n���IB�K<�ԑ't�&�d���}X�2�۱>�?,����}ݺ���98E�����`X�}@��7-NQc�.p2�K�:}�b��]F�o�u��,�J�4��K��0��|
�͗��O��Ͽ�e�~��)9�> �KK^
m0�F�^569�¡�@MyV�P�o�֡���;{�s��QX���e��ˆד鿫��b�� NP�=���l-����w�(1s���>R�b<אPg���qK��<�r���Ž���╺��. ;ށT�v�'�>J{�q�z(*�"4B�Κ��,�9��SN��Ѫ�j�*ntv��o�=ŝ��t�ߌx����<ReR�Yߞk��]x&�Acu��[�f3�۞i@W	�.��U?�ϑtp+����bi���U_�X��ħ@���le��4����]�-l0\�����@��3���kc�0���현mh�$�C ��J���L���d�d���0�ꍝ����c�,z�;�J|�z/$���fj�9�|_P�7��(���i;s� Y[�!,>���x,���xZ�_o�`�UigMi����*����7���&k���vd�j�3�22����ȼ�����̬��Eh��Bv#�ڹ1Hm�Nm��H���U=�������/<�p�-6J1i���[�S��h���k�+��?�����.@Q�YS ��nE�B�V���+ 3`0��v����-�qߟ��ތ3½t,K����\�w�(2��%����]/ׁ���b�4!M)[F����`�@yS4�I�G)	BJ��*�yUMI���8�i���l�Ay�ٚ0wPϹ�&�s��Q\Q�Yr\]i������zJ�7<Ȼ(�P
ν�ڀ4i9��Br�;��:�k|��|�{�T7C�b���",�^/�a&�����ɠ6X9�r�!�<�2�¿7~�A����ь��[���(����;�P����*D��a0�M�OK�?a���O	>R�gv���r�)�UG��
 -���֑��9�_-��b)���tzf�VB*��q�<��gJ����N'<��RAP�������D^�0�e6(�0�3�`y��6`��Yɺ�'��`�;�z�� T���53Q T���@��n1T��0�:\b}����y*2�%4_�/dA��a8��Ⱦ�l�d���jQJAc�e�{� �T*�!Dk]^i���U`��/i*%����_�/= |[�IQ�t���9�:�4�'������*�Ὰ�ytwg>��B�*\B�6���{Qn�ɞ�����"�:2=�?�<�����+8"Fq�B.�Nޒ�b�g
�l*X�����ec?���jP�f���&{JcIbȄ����g d�Xsw�$���w?z�o����-c�3T� Ca�	V�c5��?���Y�}<g�/{N4�|5���)�Q�j�֤"�)枷sޖ�xq�#���G8�E(�ߑF���
��|U�U���L݋֟�����8�#9�n$�����d�ᱼ�id�ġ�F�<md� �md����w���֡�]�F�F"(u��u
�q�$�l+ �:Ѐ���������Lۆ��M��S�i?���Xx2����NX��\:I����>���zL��Q"c��L�7�%ް���#�d��\!�Vc�2�iÈI���n*�4^���J�z��.��o*��H	�VZ��_X�J��
���}hd�c�W�����Q�2V,v���f�b`��⢚y׭�%R/�C�pU~[�-pztE������e��x-9jRN��%H��>��D�m�P��ط�ĕĢ.���v����؈0��m�g����~�]�
��rd��ݵ�
PG2��;�`�9SB"r"����\�i'��̊��}��]� {~�A���R����k�tA��7> QZ�������`9���:��%��07i�d��+ULy���`>5<<�@]�_�Q���Tl{��WB��=l�~���r�� on���x�b���� �2�6ޣ|.�F�G}�[�G3��+�*_��+Kn��]l�k��E�A�f���)�k�)���-wΘ�!ي�@���p�+;���4ﭷngI��y�0�[>�d5聳%/Qsc'���wmv��o���G���u#/�r!�5�ܼu{m,�7���ƛ"}��&[����g���Ln��1���­��i��z����4qg�No�rߡΞ�c$�L����Q5�X|��-a&k�'�#0�X˙��_C�yL�a$�� >&J�������)̀��=.���$�<��%ǝZi�;]�O6�������< �����7q���Zԝ?`-gn�=�Wc�&�C�y_"�S�Jl\oH��1� �|O���
�;;کh�#}RbZ�]UR���%��S(�<FGW��= �G�A�RΥ�Êͮ��Yf[���WB�b@���>�� ��މ�?�
5����`�È���@$+s)�"x��3g�C�� � J"+}�g��O#z�k�Ȑ���Z����2z��� O�"?�������Cm���������]�ı��v�,N���m��X/��,��F������(	�.��@�&ӿ�� ��,��8��.��C�4�����C>���B"3>�ZA�eQh&�������獙y�Q��{�1�V^e��\+�i����M��Y�ҩ@G�'�!�4��T�_��5v�c�t��������\����IRt�" �ys���<㱞"jc���W=��;R�HÑ"<{2�cN� [��9�H��$W��荸'{w�� �qit�n)����U5S�`xUg���ﲢ*��~�x���T"�ɱ�ؚ�b�蘄9|^*�H�[�;
[<%$�B^r0�y�����OcnM�d��.�ӊ�-mk!¶���M@�@9غ'�G�9T�h�f�)��8�â@������`�����$��nRF�qj��Yu�����S*�T�1p��<du����	�����7pD�u��Xn�0��X�yaxC�Q��K�k/X�묲���A'w��$+������7�ç٥�h��g�c���ul\<�P�뽝6ȌN${�w��BU�rum~(�
4+����#{���b:ɩZ�;�N���Rʫ�h�Aj��j��5���{}�������)݋t�A�w:m��M�Ʉ��n���=�E���jC�;��	.c�^Y�=�ŧk����.|T�����,��|�#�Ƭq��N3mR�`�
Q<-;��c��p��x�1��P Hy|�$T��������������i���1�[���RF��w�M��a���-��~"�s�� j %����Mt�I�ma!3���X�zb�Ԓ
�7��%��Rs�ص�b�-��كG�ׅB8x�?MYɬwu������_ؘBpnd[�C��v��A��!`#������w��^���cz��Q%�S�c{l(��o�y���c�vW&#k3w�Q��;��C7�|���=��o����>���_5�X��m��pr�ρޫW:E�	\ٻ{_J��HRqud{�K��O�>�Z�,��7��x����2���$��ؿ%�.�ҫaWs�{�b��<��l�WR!A����I����%��0Vz��N�]V��E�-`3�j�,ʳ����˱���l��.?[��"[,�D����X������a�-���� ͛�,����A#�%�>Qo����.BO�_�d�E'���˚Nky`P	��዁�|>�ռi*���:�HS�[�=�R��!����V<OL|/�!�~\0/ٳ��
��0(�n��AÓ���e��+ "h������k[�����Dj-����U>��bK͠��Bnr�E��5�Ck��G5��Mi���	R+%B��7�p�0��j��b�&�?�-t;�(wG�+ i����=��u<��|��VV��;@�H���qc�Y+(sKd�I���o=��7s�R�H?-t����q��x�ǿVol9iB�>�[|^c�&�n�ܷ #�6ʯ�09�i��@C41�}���1P���*(z"5�q_��*Țtv0�7�m��fG�]���ʸ��mW�^Ўő�`m6p*���E��@�u(�Ȋ$����]ː�����A�֌���S������h�Pw��Eu㴭Uj���Ä�OCJ��QZ.qB�N�I�뮭7���=(w��L,F(/���