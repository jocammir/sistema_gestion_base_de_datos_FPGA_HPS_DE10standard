��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0����_���3e���ӌ,nF�r9���Sْ�?�9��^'��\���G^�>I�W�UN�gsچ�݄�oڽD�/�k�Q>7(s׊�҄yU��Lʲ�Ƚ��A�@�u�3l"��ܨ�Z������f���#����z,r'_�cK���JM����p�V`/򕅞��*��F?�-P��w�T�u6c��GM�%=g�E�.K��ń� 	����e��X=� ��B_�n?i�T^o=��
���X�/�\���E�b@A����׍��ʵWn��^B;���b��z�Wh���P����͂?�����z��zD�axoD�LnʏSL1��w16J%kP��g�\q����kc�DJ�j:9S�L\�z*w�Un�$4�n��z��p�]��`$�\d��
U�Z�Y<��Йpl�����`3��u׌�[���۶�,G�J�����;m�#}z!3� yc��] k�w�����ީ��=��Q�c���l>yV>�y��)u�Z��W�<�E����%5œ�N~L�� �L�,��'���~�!��c�w���	���f�@W��������`���d�P�
J�r#1jH�nl�"5�V5~٨�@=KP����֮�{�$����c@�)�*���e��HʒeG�.����7Ø)8C;,�
��O��tG���(#�J1� 1�b6���aH�M��u��BG��j͕�q*��`X�ql�܉�ּX�G��˗�wqC��$W��@��,�_�?~Z����0�~h�
d�"����0����{{=����1�J�~"��l�^����D���ހ/����f�1y�ўR�#�b�1c8����Z��/d���չ�u���ؓ�kxSR��߆��p���r��]�b�ӌbͼ� �Vs7GEs��$z��Y[ $�d�c�U�=�2`du�؅�g۟=���������Db�&�k%��0��ڒ^s�r�6a�P3��>�h�Hj�w��� ��7������D<�U�>��]�1�d����1�O����5AU��.�o/ܺm6NG�Em��}]C��e������P��fฃfG�|ì�d�x�%֨陷��j��8�G�(����j�.gB�gV�CF:U�����`_�%�%ʭV�;{�V�����J��G�k���e��elW��"�H���$ӵ��YB	��X��C�R��J���$���U0n~��RSmM�����и�c};/A��K�O�iID�=�DW5S�s.��� l5^�d09�њ�m����Z�D� ��9-Q�XB�c�",�{�������
�`��v�ԓt�0#��`�*�s��������{T9����&�l�ד�'̐�:
��N[n�."M���Y��l���߉��Y�է�D�QZ+�]�֠z���wt�_���ol�u����W"��vX��@�:�C7L�%X�<1Ð���ge6���biʂ�U�c��Gj=o�:�M�6���
��A���F�ܸr6�r��e?�Z��.ߡ�Nʐ\H�2�Nn���'��C	�9��'��L�xBp-���	�]���L,�a��-}��Ca��r�}��-����#{�*k��b9� ��8\�_��4�
1��˒ކ�Y�d����3�ʵ^�G�l+���{)��j#I�,%+U��,>����+�N�̮��>νp��"^�^�:`�p�ܐ�i�	i�`H����E�<�Unc��n<��~�Tn����s7��$�합��FA̝�|�8��£�uB�� eix}��7/;�)Ǟ|�P�Oǖ]�����-��轞�Dq��{���g� n��?9�t�I�n�k���c3-2�S���k��k�U��(�Yb0���)�C�jo������[P��L0�Y~ʘ��r�w�L߫/�p��Itt��	ʰ���Ǽ��z���������-�.�Xn��҅��S�u���ѣB�	�jOrAL�o �-q�ӟ��\+�6���O�w�{�@�r=�mf�|_E�MBTQY���IUV��tP_m#Ĳ��KT*�Z��ԓj��{Z8��2�9��oզ\䄵��h� 'Ԏ~�l�2���oHo��̽L�)3���T�����6 <�b���bT���du����lEY�5f��>$PHe��d~wt�t��<����[aFha[L�?nH��� � #
�U+5&�r��C�XR�Rҿ������ɩ��^E�;��pSt2��"x�_[�'i�c�V@*W�<���"b{��<���gJ�
zw �"���\���|���B�oB�:@?jVP9�V$���EL3�����&����v�����$�hw�a=�ыi�x���I�8:~*�b�x�j�&�%8F���a���w����(�q��[�e���'���ʜ��8�QT����c9ބ�e�C�B[�A�{E�c�i<�'y�U@T�.�K��iT`N �L�S&6�n�m{L���P*5���*�gf�������ל9��t�\#�e�~�)>.�p����QՈ +�8N��N���͞息$
8h�8�=$(<�{��T�n�9֛�5�f�����aE�O��������8`"	��S�ld&R�u�qv�y6��w�]ۆ�&�-�YQ���@	&L�_��V��e4����Y
^��w7h[m��ν��o�[s�8,�����k�|P�8AcA�e���������V���.���`y�@�%�A��_�кԑ�����<���X�W�e���ݦbW�
�l��\�*O:A�j�ߐv��>G0"�_o���ֱ@M=��^[�sxf�O,�5ܓ�Y����.8��X5���ʃy���Z���b�ܢ�Ku��L�fW��q���evY�����?V�gtz'Y��!��"4kkD��-�HX&ӧz_|S��m�p�4���=J���!����Y���G4�h��Ϊ>��WxC���sHL�/�Y�)��)X�.��������tfV���]1uU�tyK>�GdB0X���ŧ?�U2N47�q��6�(}�M��\��?�M��Q��8~����G�u����KTk.w�P~P��W./x1Y�W�xΚ���r�ܘ�bL���t�y�N?�둱�(ˑl1����Q��貰��Hl)��ي�15:�&�:|s(�X������@;�v��@0I������TW1��.�����D���=�787p $��?�X'ȭ�<&���-�Jk����(�(����A�9^2�<��a5<�x���#'n?8hL/�����ȁ�F��#7P3]�����|B�w����4�9�/��͚U}TeՁ�&��U�3|�\��a>yZ;V *Ϻ�*����vR��}�2z1�^���Ѻ9�O�ߙ��Zy-~绨����øZ֍[�c]Q
��5�x/;�Xn�7��'���w.�ξ�g���
!
x`J���D��5j��z-:��	�2(w)2�Ѳ<��L�
	Q�`jQZY�b���]��i�Uw��AL�b�+���E,���_[E_k��e��3����r�;�z�X
��ЩRx4*��VƜ3^��{���r��x.��Y��F!��n(nsl�
a��M����";V�F��s�:��sR;$�`�ݝy͔&���Թ���L�"�d�!B�^#�D-h����F�����D��h2i;UX��6%�Y�r��nB����Kÿ�HJ.�Z�%,�@x�<>�7Ϗ�XW�!Ҩ(��d~��%a��VR0���R;	1��`p	�9`F[���Z���A{�ߛx3>��pb�K2��i?�Ϯ1�Ov�qEʿ9d(����k��B $�H��<�T�����u��{��%�=$��9`h�Ǖ�P��^��"n(\��O��vz5H�G�tr�`q�������:S�ͬkI�橓��@r �3�s>��Q!�Um�y�[9(���Cg�ۇ�LY"�1�vnL�}�m�PC�+�t���A��Sl��y����>'�=چ��3��T�
�\�����ɚ�"��9��77.����mw�-����#�E[焠�fn�D]7#L�B�ZM ���T��G ,��������b�����='�6�������Q��6�gT㎓9���~�y#�ſ�SO�8s��v�OtNbb��g�c�U,"u���L����b,������3�C�s;��7Uk��T�f�	�K��ӷχ��:���bXC$�Ηt���]}���"Q@rs�"=�ޏ$�4�}�$)�R��|fm�+����}d9��O�M���oEZ���)��ݽ�lƪ�r����ιf3}03Q"�N�����6ځ��ն��6R������ԛ!K̿;���=���'EÚ����	;8�	������YT�D|z�h���E=��`���܄p�<㆞R1,L@��G���ۆǵ�\�������Jo/��2�z���W�P3se�+.[N-�q�{�a	+�l�FpxԠ�!�������렍�L�(�hlFf�mYD��"�����s�	IC��'��@��b�9w��&����F#��@����QZ����Q�E?�Y��*)t����^�� X+Q� j�}�Έ����4��]YO�����R��~�y���C`�I1�n��E�q;kx���#x:��� ���WZ���g|�O\	r�k���:0V�v�I9�z��i/Yb�@�u�DbX�_�CHcBA2��\��Սj���5p�mGS�p�u����+�&5�i�~ܾ\UF3%�
E�څ��q�g�}�p�MD�BJ�R�d�ʗ�6Ů~��D~��ݸ��Á�4��N~n,���hj���o���ħP
0���8�wX�QIA�-�v��C����!�p�w���d�^�;�ߝ4$�k��h̦���I�����j�ӈ�9p�(�v�+���|0�ڋ�tS[��%�;k����������`�5���gVӞ�[�i�b�
�\���p|�]����9^-G���I�JE+��|>���*U�b�=(�1�ۢh@�k��pz���R��fE����Z[I I���QpsB��p���18�Tm��P��cQK����G�=;^L��A�8O��f�s��S�T��sX��K?)�z�7.��r����4<'o���k���(�͠Iڄ+O������Sb��8L��G�>44'[u%b���[�)=G��7�
n�sX�k�W&ZJY��~�pr�2�$k��ķ�GU�?i\���n��������=���K3Z����
G/ur.(�р~N����Qh�Rn!���$>JK+��{�Z	2^�/��:u�0K:���j��_'8X���]�{"-��D[�d����9UƠ�X��R����9�^ |>埔] b�����ZD�ұ�0�{/v�q������6ڡ��P\8�ل,�e=V�-D��VZ)���
�wS�(�/�l��S�QUs͊��@溨m7�Z�1Y�UAF�]��d[�y�@%GjΘnx��T!������^�ؙ9�D�BZ̮���N�u
�p��z���x����(K��_�2>��U�����^��P�s�^�� �Xߛ-9C�M`j������)zW_�i�
G�����_=	�
2� ��?����jN�w���x�1ds���٩�*��pqP�Ȕy�Tf���;ۿ�(T^����7d�l�֋��1O��J�.H��s��x����Nc�^�f�+u_!۵�|�v��=S:Z�>�����Pd8\ �mz��P]�V�čѡ*�E;��\�_���DN�'ֱ��o�k�:3^�`l�u��k�[;�'>"�wK�@��1&��u�x�Y\r�Gٹ �S�֗��v�H�!=R�^���e��T :燱&j����̕��am�5q1#�������˄v���D�.U�?�$D�����a �m���MS�$��<�%k2�����z赹����l[���$� If��ovPz�I�)bX�5�6@��f�ßCԹ*�-_B�l�%�,U�jB��W�,��F7��R��+<J�= ��>8)�\��i���� N��f?~1b7�bvs�
��Z`mP�7�0�{�뫧xLTx�����{4�3t2�s�λ�ӧxU_��F��Dbˀ5!(��NrTko��zL�ee�������o3 �!nᲉ��y��A�����$�� �o#Hr�����_���Qk�O��@3C@
g���5řH��^W:^z\V��T�͸V:l��L��4Y��\�L���esy~5�\��o�3�G��G]���G�kvu%W\��2��7a���Q׆��K2�R�v{rJ��q9�4z<���N�=5d'���+��������̲���{�B�"�eS�P�՗�O�2ZS��H��đ/8�N�9�Q�Q���cO��0M�4=g�z���fӢp��Ȳ@Ag�br�:����2�+�ה9�k�Jɯ�و�|�f�~ZU[+}���#zk���Ra4�*0y�*�gtg��U��aa���_P�p?Q���_�g��9)���ϬG�ϔf��k���H�X�8����F]	�;rDPH�Y~�f�o�SJ;����{dp�^����/ף"�����0��hj1:���H���`��.�07���A�.{�"�+(v�+�}�x��������A�q�O����3�u~���Ő[`��.�����"��d�r�}�DOnnͼ�~��r�%o���*3k(lO��v��x����ǐ���:�������5�5���g��뚇�aUr�E�x��a'M"V����#t�yʕa�`�Ն�����V��8�[R��~mi��7 ��?��S�Ɗ�B�� ��ߺH(*x�ʷ#!d��5}�)h�Ka�L��	�Tg`u��0�,�!.�S�m�W�
������E�^��v?�+2���V�M�?X�9�p���tyRyJ8���Oߌh�E�=z(�^�'!��ࢍ�C����6v@�@M�L���\%��eM�$���H�=�/�f� QgS^/�6b����Q�0�M�.b���Ba
a�qv����2!w]t�5�`���p�?���i�!�e0{Ȁ�F��� ���}�~-Z��e?��� 
ݸD�U�*Mo�� Q���Mnn툵�.�~W���c�*��˽��g�qB<�h Ƕ!��;~��M�4�@^�� �1",�7�ϕ�F�J�����_�V.���:͓��2�Ţg"f�� + ���i��WG;iϰfu�\�@�2���vCV�)Vu�����+����y,��_��qn���N��}�_p�y��g��7�!?���!���e�猩P@�{��U�8'�P���	�W�N��F��I���Mg�M�:��i�4�nc�,	�G�9�
�9����P"���	�i8�{�R����L��i��?X/��i,]ss�i��7V�Ń��2`��/�Wy�i���B#>��h4M�_4��GW�[*>��{��5��`<5���^�i��K8���	`PM�M�"|�97�p����	%�b' ��=;!�Ó0u+"|�ZTP{�g��,������8�:0e��Vu7�rʕֹ# ��-�T�Ŝm����G��"�/��{ġ���-"�(I�`�c�AAb����\t��\�~���o�>��N8'��V�ܼ{O]Ԑ���a�� _Cz6����M�S�0��W��x���:�/��b��O0��h����h����4��ĦBv:���5P���Kbʙ��шg��[Ȯ�d��0������.l8���z������b����o�����)g���EB��Oփ�X?p����p�۫�S}�k��hcg���]E돸^JX���í�'�@��_��I��۶�;�k����K$�~�3ɽ,� oz��A����.��"�R� ��4�s�7���Ŕ:^���T�C��N� �nH�\A�,V�F�A#_�
�`�@��{���0�&����r��w:�}��x��M�MXou,�F��`윤��7�s���{�m��]�%h]��E��^qLD�\0��i^F���\����l��Э���2���-�G�){`�p[��`
����Ӧ}g�Һ�i�(3��)����IC�������n�/R��D��~Ч�#4nVy�:ܣ&o�#�=T\���F_�n�A �<$���=�G��"�ɨ`F��b{\�>n��&�c���#|��5@�s���}��!�<TB�b:Y�Dp��~��B�CK&�r�ՀrGI~����Dٻ_ҧ�э�9pi���;�%���t��B����.�}�Q�Y�r��#޶�V�eDʽU�}��L����2��1��\�zU��:��构1�Z?�u�گr�/�S]�ۅ�d�K�m%	|-��D�����!�i7�d�ʻ�Pڙ��}CMp����8��L#�X���]/ ��X�<��𛋜�$o3��21�u#2�O~B7�9��x֩�����3i������Qd��*�Ǆ!�a��"���	la���g�b#�M�$X|@��L�	d;���w�]���7���^��ۚ[atT�6��_߃�^Gϩ��Yx����~����̴s�t =�|2�`���i�b���j�|�����1J,�����͵w>�rT�e4���	HQ�h�e�O�!�.>*$�`9����磌Ɋ<.�4�ӎ~��}��|��us�M�@�&d�k��an�a=��`<���2?Eq��!C�˫H�m�3~`���G���X�]�����K�
#�TOU%Y$���'
�l_��[Q+����N�2��,������" &�vY�ѣ~:�"��.��[Hy%g��O=k�%wI��}�ӬG#��4���q*36�7��:g߱�߿�4�n��9�ib"��P"��j��lY�T�]�h�[0 _2��k$��cԄ�XZ��|\�A~�#rd�]O�+��P�N�g��+H�RvG��nנE�;%mtŜ '�C9-�!�ē_�íE�g:�\S`�Wi}����"퇱fyl���<Fok���4U��a`�O�/a<�����3��>�$���ڤv�辮�yǿP�'��������ڣ}�đ�%PJ+�#=RS����U0R��s���V���5�eD咸3��*"�8��4�	F���G�ť,[N��P�T�,z���R�)�'�Q���7�y7S�n$����#����x�������5y.�����JTS��F��������Or�����7w��x���H��B���DF4���=I�Q���YE����NQ��X+*󝂚*��C�ĝ/8�T@�a�Wږs���J$éL��zEs��i��Y����`���mU���pW:�o66]��G����1�9�E��,�c��4�ǴE�"���܃�a�y��Q��C*�\@�I�!��#ҋ�H���B���!
{���q2�w<ne��7m����=瞳�}?q.�5ȣ;���Mm9�cnw8c.xW��HP��(�>���-���.��["�q�(���e��~�,d�3p=�W�^�_ZM�q4�M��k��\�K�����g�q#i�2����y%,���V�0.�(]� ���.|�W���6��������5*l����q���I��Y�B��è���8w�wU�׸Fv44�VR�^��[�mq�tIT|wƱ���Z�X�:�W`8�%��5{���Z��ȋ�Ss���
����aW��9I�-ŽM�n̎��,v�J�rrG̿L�9���_�:`p�K��Ä׽���!�I��C#2�����pT}�ln��@����=d%�S]�7*���f~ZL�1�ł^�&�䙄�t�c����NT��0*�q�sc��z�@z(h;/��YS�����թ����0A/t�����`p��4O��ߦ��kGVO���-����?�z(H�.�o4��z/�qa%�^zo��{>��F�!Ϭ�[������TǁA@厰?I>p;'��_�����ْ�3�F����`�r&��׆�-�*��}�?�PĻ�C+�h�X�����ٵ��`e*�x&x��DiJ�Z9�o�<�x�O�b�l1H�%�<ryǦ���u��ׅ����~D��)���<�k)O�+�#?�T���z��>z�Vٽn*�H�j��z����&�Q��*d�o=�wu��K��ۄs73�H_y�r�0
%?]��"��w��w�]�*�,{��Wԍڊ�(�2Вuf��� ۶����#�����5˲�O��o��	/ӕy�Ǣk�#=�@E;䞉�xr�PB��ލtp��� �����🍉��]*�wJg�|OB^�K	�<z�4++4l�F�t����tY<�2\G�i�n��g�u���Ts���_Q��p$���S������"\�����N���������'Zw&vUs�8��ƀ*T�������CI&��z�C��	�`׸a��|5;����k<�OdӅ���[Q�l���7���E@���<���������c��{b��$Ff�����5M �\l��1u�@�n�� ���h�2ɗ�Oj>g]	x��	� *���D�'���ZߜG�ˬ�s
Ӊ��Z~�R8H��T�@>��R�W�[�"���1��W�k����5���i�e���1�Y���P�,.��-$��a����'��@�:���f 0s�Dn�&]ˏr5Ø�!�~Z	m�`֢�^�0l�?��+;8�H茳xe�kNgJS2��mb�����5ޢ#3<[~��� Q(�*�D���B@�E���|JT_N���(���.�qꅨ����cL���5�W��R��k��(�84Y��Dz��B���F�����z6�Ϯ؜;�幃覀��=g�6�&Õ�n"���"\�$�I�6|��3�������=:��)E������^��5�4/�O�Eo$��@:���<�����+}��N���0�� ��<���d�i;��d���ȧ��F�*~