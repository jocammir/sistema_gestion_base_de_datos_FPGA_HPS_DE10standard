��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0���p�?�gu:���@�6h�B 6���+�Rw9G��KĿ�n���4����]�����"!;ޯ	+6|�%�h�JOe�wX��r.�s�7�)�c*Z<3���ŷE	o;�^;V'�gn2̡k�q��+A�\y��ʶͧ1���v΀�,�k񉷎H��+�*A+*j򬍵쐄��s�sv�2L�
��vc�QkܭȲO:��J9�UT�4°rVH���1���N1��O5@$'�A{_k�_�)�&`'�@�ff���{�ʧ	�{r�"c��|z#G��:�jM�`���A�p,3��oކ��/�L��F��vp�?�7Y���%��!���ej���ɫ���"��%��ɤ�#�E��c�����W��$�����/��o��;�fY�3H�.�~oA|#[>�l�\�{�&�Y�a}�e%iN�[?TY\��ުV"����������_L�e"v�D�q�~��,���!R�z�q��Ͳ��J�=O%�r�j5��Z�Y�*��ܙ����~��K�4go������8�64�ߞc��Ёo/�C�-𩁆�.w�mI|�#a��L�bx�8�;Ղ`b�����xwN3��}�bC�,�Tm5�Uz�w��&�V�~>�~���]�f��B��g�E{�#&SԺ��Z��^޽�^qBt�/u\�2�촪|���S�=u�^��)愈� k�͗@U�����<C\R�&���
/>b��|��(��9�LK�ɢ[ S|������D�Pe�NRb_N�odX��}(N�-��
G�Dh@����~�7��ܷ�9����&����oLl�}3�Ń��|ׂ�]D���JU_����\9�bҧ�c&�%�?�<	DH��Ypr0�6�9n���a�pH��2��&��!ж+��6r�@6k�g'BK����S�3���/� L��?:��Dl�6W�IK���J�5^���� n��6�.-˒
��O~)!�ءB��%�Q
�8::e����L�&xD�2��ڧ����@�,*|ѳy� �<�
��=	�j��᤹.��'�T�"5dZF��]hlD���/	p�h�66~�`�1;���S�K�Z=>_����z��˩�<t�k��/�y�z<坂���e�]r*��z�VA�gՄ�,�5l�.@�����Y*�P�
�`��,};��Q���i���-\#���Q�DDu�`���9�k���\��^�ė��q�]ƺ�����뛉mص��V���}3��B�����8]�j{��Pxw���R��o�|�]jH���ۘ�סh;�D,B��O�*��Ӷ�7M�*R�������$�ք�}\E!~��J ��Y7c_�8"�As�dwu?��K�������\�Loc��0�Z���W�ɹ���ؘ�,���q�|y�?V���\��/z�[�Z`J;�Q�K�xj����p�1C�~d�*�g��eQ6k�^���bq݌�ɓ6P�=�l�M���Ȧ.�$i�iZ�'9_(:��T��YǱQ�8e��}��Y/a��9e��YY���-ػn,�lh0�g3ll�a0i��V��>�ʄ	����e�@���l|��J�I=<jf�p�3f�y?�4tQ%�A��B��y�Ȗ��J��t���Ck/[������Z��CY������`b���3��RuR�����9Y�򘢇	A��h&���}X�@��6N��H2��:F>L}�#��'Ꝅ$�7�����Ƭ*� ���4�>[�W���	���Tء�������h䇂�J-P��]� u��g�5���]{���� n.K�¨���W��3��aI�5bV���¹����0�N��fgҜ>�Y�sj�Ĥ}�z�T�=Cޣ[=0��H��������a#�r�=A���z��"�7�c��Xʄ��	�VkA�`TN�
�Z��B7��K5�M�����LI�D@��coq��u�N��.���� J$�<?��G��C�|)��tJ��xO����C�j�x�}w�#���*��`)J�5e���oLgC��i��0r�G�\�ztT�a�i?�Nh::�_U�/���y/oK(�Y��4�����8�ԅW�����IZ�LP��1G`��QI�x�*���Wv�~u?��G)49T b�Z�g��8}'	�_�3�?��nq����ȁ f1琴S�V�FT��ܪ+��{q�g�aw�Nt����!���X�x�;䴏��V�-w�}��!la��|��X�(:)2><V^�%5k����j��T������z�{�2ý�������n���q�Q܇8��B�"��GR�0'Zq�h�����o)��34^s<o�)�`�:��`�/��Ԓ����#��M�o�X`I[$�*"���1�k�OQ��ě2P� �B�D�-i�*���u&���c��=|��%;[.�\�߹�$J(���@UІ� �Ch+�Ԭ��ȣ������L؈����]}yA��O`lɯ�#��eP�����E�3寬���(G ���f�zև��ݨi�GI���0b�}Z娌^Vb���9�V{c��u;PN�lU=����J�$�ҖO��7��s=0�K���Q�v���Uzu��{aQ��8��5��M�Ӄ�i_b���xТ�߈��E���そm����=����c>��7�Y �:�h�R��Y�15��8�B���E��&�JH�ee�i�(��m��vh\ǝ&�%Aq��\>8%ŏT�W��g����H�� YD���Eh�B��F�4cD�ǟ�p3�.TS��"T�&���!gxZ9ݐ8�,y9>J܊���}5� ��6>�4|��U�[ؖ�E�?�V�i�� K����u��+7(�� "�M�vHx[�8��Y�%e1d���(R4��U>��%TN��:)�.Y�d����z+�giU���k:3�@�4�t-~�~7�k�vN�P�Z���*=��сF�1:�����U��8�_-jn�m���k*�HF����:�>F>�*Gj:�g͓ʏ�\�=���5+��� =����j��Ɛ�/:�h�'�+v�������������e�<UP@��	u��t2���g�pG��Z��؍?ܱ����ӳF����vy7�5���r=ሷ%*��u���J.a��+���r��a4� ���-c$��q��G�U��-�C�Y���R��D���>r����}��Um_vfx�G�Tk�.}�qV��[>�a��<?��U��e�W�~P=�;[ߦ.B��樱��Z:�&��7J��~�h)s��6�g�LoC�AeM�<��<�m�.ߺ}G3c�_�; �/~¬P�C��|�W�q;�-��gn�FZ΀�'���قD�xpjY��(ߢ6�4���<	����U�x�|)}����}'�*S\��u��sa�z�T�#��pP��e4�����(��薸-�=���K~�V9�#��Y�'���c�>��9���VPX-2B���`BC�w<�5���*,E�o�;��S2�=>_�e���3uI�ɰ��P
Ru;��(7�sn��y������nz�$�������˲��`:L:b��>zB��ރ�K#d����,����WW���=�h�0�I�gN9=2d-,=M)Enjew�\6q���:H����R'?��$
�/ &r��C&�����=Ju����Hk�fE�Ԙ6�-�K%럑X~�' �BeT۔1��C�űucJ�T�4�:*6:&�{��$ԮmzN�BR'���E�te6���~7N�δ��B������Y��Y���	i	�D�Z�6;��Z�J���U�4Ɓ�^��
G�x�o�*�>��;vÛ�`�:�n�HƢ�\] ��������@LU
5�k}�Q��lK]� S�ׄ��U�ũ�o�Odb�N��)N*tg��˵�ƀxe@`�3BqRq� ߸p=0Ӄ�F����^M���S�%j�4������ii�Z���R�����P|Z����*�`3��[&�����&~��]�o�NRZD&Y�3XNCK"6R�|=^��9)g�iհKOn@���j�Ä��sUI�'�V�˴ r�:�ۡ�r�n@H��s9��$��;ߕ�~�g�;���-�e�*/	M���Y*����3О�ۂҡ�U�/uU�U�'ҟ�TYض�:[~A�O��^\.x9��va8���ۡ�a{���H����?�M�6W�.�f΄3�3x%����%zϭ�3W�W�z�U2a��	mI�6	T�+�⤊��jmg$����NAf�[��/7)�9���O�2�q�z�<�K݈[��'���.�$6?�t�;P�?�y�U�P������I��P�џi���3u��w�1��|�k��U�]/(��؂5����7|W�rIs��r��R)��7�XQ����N���±��4����p
��L�+t	���խ@��:]��͜�z2�p���i¥K)�cq���������C\�c��M�i��ߚ���֍Fd�� ���0d��	������ڝ�B��f'����*�~�ƚ�G��}^�@��7�M����St	����yίjI�bc����e�b���:��+�j�yx-�f��n� 5]�����w��:C���5�}�C�׺�7�i�Ώ�ϡ�p�����K y��-�i�1�	O�K[3��28�+�D��T�93���*��������y��F"$[
����	y�O��YU2$;��Y�R�aFP��.�{4TRo�[R�S�k�[�������h������n� �k��$p�$���n'?����)24^u�=�葡��ss��zxUq��Z��K����[�W�4��z�c3�Q��p��d����'7�
Dq�h�P� \%���Y�%:�fM	#�@�`ʶ"YC���p�4��w�,0#�JeZ��ב��WK4��z�I3 XJ�D��0��~�mn�8[���OC�zE��U"�Yb`H��bg�1����h�6Aiw��R��)�a���j��>�V8�O���7+�Z5E�����W-�\��0ge����q�T���tQH�S�;��)�.B����o�3����#�X���<����>������a�5kG.��_�ѐꝺ2�
.:��D�?��"�i�O�p>6�>�0a����³X����oT▴�ܗ��Oa���S��~$D�ܠz˭�)����)Z������)+�@4��'���)����,��<\���r_>���4 ��jt���c!�4�>$C%\�k'ulΗص�KѴ��\��tzɐ���-���=(
k�I�fZ�K+d(Z��R\�m�r1��-�Y���F����zs�V2��s����h���?�s��I�`�N)��Y��ɨ�)�����̕q�6L�R�TH8�	8��m�.'�=3�����s��ą��