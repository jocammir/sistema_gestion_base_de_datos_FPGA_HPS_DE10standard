��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0����_���3e���ӌ,n$85�J����D����(�j����R�c{�s�ZP�D�d'`�L�j(Y)������3���02bcm��:O��.Dk��/�88�8h�!�,*�ow�;ϞF�Y��T�#s�X=��V�$���6ߏ�/�l�ص�$+�H� ��J����~��
����΂�i��s��;�Z�ʳ	F�@����d���پ��lO&c����<f�:��/���3,vt�W����\."g[����ߤW��8(�M\iv���*��tK��? �~Wl��f���$��P6���/<8ؽ	���=�=i�#�Yʠi�'��?��zt!3�f��X��鵓����}K��0qgbk}ӱ��+�V�<^#�����[lIG��#n�b#�����ר�b�}���
��K�P�׹9�/	�l4�+#���l����e���O�xE��� "dEzﰫ�����UN���Xg�����~l^�<- ��f5:�w��-��HF!���x~��>�De�@m��_�t��h�G�x�ȡ�~�gð�E�	=I�1 ը�SkƋ��ܹ��j�W`���S�~��Ԧ�>��w2Ό�*`6���R�"��mI�����������%h���/Wbd�]�Rz���c>�o:��1I��Gv�ZiN䏫�N�q=�/�Q���#�+�M4��I��<m;�L�kw2�m�̰�^xx�����Ps��]��z�]g�Af�Z�
'��R�n#|]1ʉ�W��-�)_��`�^c��d�Z�H�"��5q���|kB�Y��d`�s�-׸>B��Bv�Q�M6����r���1 \+�UB����3�D'������;�|K#,�Qju��`���.�Q��9�d�I��'��� �n �����k��dhI�8T�@[�v�H��Ή��4 =`������6l�	U|.�W�R���S�䅐8��W�ތ����&7i�x{F������ך#z8/�m=��j"G�I$�9I;ن�>m���@�Ï�&]�����ն�dJ�s#�k���.5�'zd�7�a��3��a}���S���_o�W�\YLsL�/a/˫���rL;�\��}M��9�Ig�
�\�1<
V�\�v)�H4��sʗ��xٌ������M��G�C)p�"(U���u������7�&-{��6Be�����U�A�ld���M*Zh?���s�䤛�~Xֵ�k\E-�餁�뎶���I����rN0��⦶$�2{��)�25��"
ްC��0���?��_���ND�w����߾�ܡ�Y��\Ѥ�hv !e��[�'��z 1�Ќ��+MBi`��v�*Y����z������^��}c0�����:�������q�I��:���Z㘧�� ̬�~��F�k����s�z4�e��|z�w�٠�(F��d���4�u5�[��}�)�o~V嚸��q1z~h����leԳKVN4�Z�rݛS莒]2�!�Tx�}���K 5����!��$��-&�BT}=�^���R{�=� ��W��8�C"c(�̤�
�g��:A��p7�O�c���)���s@���r�JΗE���o}ؕ8� OBB6��<�2m�&jD~G�����1�G�~���S�1�G^�r{ٝ��K��&?䒒Xk�#� ����*���\�:Q}�5Pgg�:(=4���N��ԅ;$9=d�2%v+U���~�u�S�+zH��P�N]m(�����yISjU���^8��7�Ӄ�:"�D KZ@N����I4�������a�e��K>_�����:c=zK"�!�/ԏJۂ�m���	��שZ,�|��	B`�#�S�[��ýh2����-��ɟ�bŲ!�X7�� ����Rf�7�q*��A	T�Ձ�A@=Z�ؚ�������1զX3k44�RN���*�ƛ*�zd�Z8�Ա�{T����b�`�\����kM�z�]tq���FɞS�I^��/����O>Kʏc(I�]��[h<= eO�&���C���+�	a�,��G��>��Uk��*�%�B`�1����`��fVdc�D�A�:���B�xa���y�5kˤ��+@� ����i$ղ	zt���g�k���K��! ���8�i|��+���6'�o���W�of��Dw!��$�bO�����iHEC��˨A�s��"P�gU(�"{�۸5�-jnmgj�0��C]��@(�	���$��3~H��)�Ϗ���Layd�)L{��?�z��1%���v�K���+Ѻ���Y}Uܑ���@��-��/f��1�4 �Fұ�敡�4ݏ:n�zP�슻��� ��F�́A"(����I� ������m�dv&	:/��:���@�0g�5�n�G69��$��D&w�l�w�c�Юk�֮&\�heL���T����������/n(��2�pT�q�Gy(�@H7��,SL�19�Jɒ)���m?�vh�^�8"/ώ؇�unk{��l�Dդ�
}���VC_��P��+�n��d	�E�9�>4"��VM�$?SG�qL�F7�i�ҋ�:3�ώ�B�f����Z�;E�9�/C<_� l,cl<-�V�R9e�9��2|�Z � �����3~舥��I��%i.D�ׁ@H�%E_Ex��O�ƭ�j��q��۳÷�M��g28z����%I�*������C�)��3��Ga�:�.ß>�$Hi�-���Ư ��Z��9b׽j?$�2赔������-��3N*bALƴm4��N'6
ƴ`��N�8��T��,�����ݕ��J�rq�c�o��eghQuS�GJ�$��x%�o�����������3���FH+�-dCjV��J�	WNED�1Η���0�D��e����,~V��������A)�����\0��3�:zDWb���w� �sc)Ȼ.�&;qz ���sr�91uE�'�s-q�҂����ݼf�i{鷦�(���2�r)���w�uf�
��Y�@��[���T޺�*��D�蔔�jG]�TW�Ǫ1��޷?Q��L"��ka-x�����$T%4��h��?��y��R.�[F���R�&C��>���s��E�o���䤸kI��PJ%@�2������m��AF�9nb���!H���"�z3�Ŧ���Jf)�s��ǣ#��+p����,)�a�~���
 t��Z�\��s����0z�\F�������)6���t8`��h��<��6�qG���,�Ft26��G=���+in�k����Do՘j\�I�.�cQ�7	��Mk�dB� D�g�����K���S~�y��>ă]���ܛN�5f�,�^ŚG[���Dt�����v�׫F����ȟ��8�����L�&BW�l�M�.�ѝSkc�d}	� X!�K�;o�!�B�a���9ܾ���c��tt�	��U�v��U�1&w�� ���V.���������NX�K��&�|W5�	$s+[�fch��(��F�C!TQ^>��5���1gЄ~�
625�����tE��z�+IW��W�����^��!�׫e6�G2�?T, �������|��"�X"�d���D�(g�ڴ?lmo&����=��|�/s�d��:�)~ͷ?cR��v%4U�*47�_��<�W�BkW�E�k@�~���nuu�?���@R��
 Q`1*��j�����YJ&���-Qs�����~GG!�P�!���Ha�}��bs�ܟhȻ�(?%�����nI����c��c�,zȁ�C��qMsY��diFt?�4ᅻ7I{:m�i+��B�$J�fBpTN�Q��٧J"���*�������,g��$Cmy>��vN��ZR�7A���Er��L������a�����7�"=���n��6�����*Rq��'[�/�)g�@K���GU_ք ���k������������h�.�kO�H��!��pPP
[t��\��%��9I�i�8fU�J��!~^�{�&`-/�����A:��5��I��6U�WW�����h
P�.��W��^*�g(�����*%ZEu�n,�����81�jSl{��c���52�6~ˆH�Xm ���Է�LƘrgv��������ŉ�7��y!�����_d?�<�쀵1���B6��C��i@��g��-��)�=~�U��KcQ%��`���*��G������L��O�RI�o��74����٠��A\ɦ�̿(��&�]�}6(��T�H��0��>�pptDi*��T�C����UV�����Wk/��L焕~x���y�d���%���_�~-��fy[�Uyp��C�; �Qɜ�x��ǁ[��97)��Y������5Eh�+:�j8�n+:�Z!�<�J�h�����;o����~����A����d�5p������Y��&�ݡ����ϡ��֎��;�_ŨGݎi����iJ����vq�b�뼍���&}�390|]G�U����,����<��I�f
oGMzm�������;��A�c�!�xԽ�~����Y�H��>M�T���*yP�H�w�s��q�K��F���@-@���ڐMuԙ	�Yb�3_Ϭx�!�V�ZqXd�'#�Na8J3̾��d	u��k���AuhX:b"�WfY�`W��`�zg>7�1l"��O����������{�͇���Q�)�u��[�M��Ǐ��r�I����A4&c�|��@u�hE��̢�E<r�ꭾ�u �A n(�$�����vb����(������]�|Ǘ��ޝ����BkS�K�W����S`�'�Zn����V���ƹ ��$�����і�j�Pf<#�g84������X�,�����'w=}�l��V�(ϫ�
~,*t���`�V5�V*�$�ȌF.��!Y����Q�Z��2�.��x�P�!�!��MZ�ǉ�{��tΡc(���3Q�Q��Z��@�K����t2:+��m"s4P�W�#��]W�-,zCR�@��جrQ�(�և�c��о�]�Bgd�	�h���E �=��_]v�h�������r�[�*�pnY��vi�����;
�^�𭄹	1��8=,R ���t�@X��̤&$K���e���R̄]�]�Æ-�.���cj����Bݒ��}`x����Я-��lj�R�]Җ��W�I
�=[l+���d�h�m�#d�
��ȱ�GoU�H���E��, ���\�J��	}���\��0Z�FF#�RI�x��^���7R�v8h�'B&��!˸
B��/�5a�A���R4��t>2�ar��i媏��9ԏ5z����n�5�s�GQ����;�S9(	I3Ċ+��A�ķ�-u� ��u��r���qʰ`�D⃰�NY56J�B���N�df���L$;R�^b�_��`<��I��H��GQ� خ;M��؆��j�^��ɫY3Y?t��W�ӥֈ! p�A*7�zP����Fz�_C)�k������^�C�19L��J4C�{����X�!C�a{�m�Չͻ�e�Č�{��J�mj��'�*��٢9��U�E4��
��m7Zpd���ґ��RV�D����NnCL�z���\���z �K}�-�ᔑ)�� �@D��0�r����!������=;\+w��E�ܶ�W�TZH4W�bq�r��E5,�H��Eԑׇ��Z�K�B�/�=��P����0ݾՕ���6�q*���#=V�Ƌ������dX��)�4y
'&|�}\c�Z���!c�0F��þ}�I�FPX�{u����k� �NVa�^ׁ]Ңs��/1�J��NB7�T;ȏHx:�N��Y��7R��~�0<t%%BI�*�s��V:�r'���'��mW<x����tB99L�#�A�]�=��[!�^1�R9���-�I�݃�zp��x��qV�M��ģ�੧�@.m���@�B/�ɜ��HD���J�nPSV��p��.#�fX�7���$"��JX*0i��&�@[�Nӹ�M�+R�N�7���K衳�dh��� Ma7	����x����/�S�#qN_�^K��X�@���t�J.H)�̬�*^"�*�	���Mp��GP�{K�Ƅ�����i���Co,B��������">��Y��%��v��HKF�E� �ň�Ƕ��U}���P�0E,�]�u8��@��w��
�Ŭм[�X�i�i�( ���"�� ��oU��jӾΪ� حu`o�]�K@�k�+J�F&D�ŀ���sں�jq/I�J	N<�bԥ����y�c%�hf ��B<T*:�3����q�2*�n`17�V_t�IT*�"S�U�Sv��|�5ɲ`��SN[˙x3<h�K�88`�2���Y��{�q�"C�\�n	E�o=A1R2`�똮��>o���b�9!�C*裵�@�ݑY�����a�3�w�8g!���:]T�3š���M���A�n�7^.�KSSB�1��4��@���[�%A�Mr�-�����~�嬘�&�-G���U�L٨u�M1�;��9֘`}Z
]H!��lD��(��z���	,'�lYK2��G�*6��J�Z9�w4��ئ+��CN.;D�R�����0�b��kH;i��� ��q�n����썄ƻ|��% ��K[���&��ǩ��	,~���ە���.�9�� A�����腹j=w ���!M�)�ٳ���`-d�̝�kU<uxz}��/����Գ��|������k�L45���҄�m=�%�rԔ�����3�g<��Td�������J�S�:�gds�XD����w�*�ƞ�g*{ӝ"�Q��6d��z;gFբ.�3�]�0�>������H��[�blgqv�|.��Q�������M�	I1��}~�7���ӵ����*�j��K����� mJ���MV�����A�P'a���7��tVXݑk�21l�%�޲��s�99�z-��v�F��!�����˧�x�9��}+Ӎ�UTC,��~�qO/�|����TՓ���ds�c��9ز^{�h��╀�/椣R����7��j�?u��o^(z�E�C����D�K ��ހ�ub�_h���Ƃ�`1x�����4B�8��;.A�����9� ��\�D�\��_�bT�mSrE��T$� �h���[�][3ƨ���E�%oTR�I��CQ�f��A<Hu����xV�C1��H��P��e&ʣr�}eYRI��}/Er���eR(��p&����Mlܯ��86eS��P�``/�b�=ڲ�=Z|pcw�AO�~,�|�/V�]Py�M���Jg̫���H����7	/<'�)� 6H��$�;�E;��b�m��1?yp��=����q���#������N�?a�ROY������C�_���ޤ )�"�܅�����"cy�I(Q.�jT��^9�������4��rL�E��;�ؙ�����X����+H!l��_Aҕ]��8�2j�����3�i��"Û��e�.�[�$U�ë2�gH�%����3�i]��P�j�t�GbR�ߵ�$�8U���Ndg()��4���	�m3̹���������Q��L��;���Kz��{e�J�u����Nc�`�7`R|W�-F9�w��eZ�4Q|��\=m�&�a���b,2`x|��X��+��ag���b��,�I�$V��Qѽ���6�T����ՙ���� ����>� y�Gt(H��G�vq��1��p�D�Ԋ4	B+?۳=X���,/�P}����D �;�A��DB��;���fQ;�-���Q��nyD�({
I���]��q�x�RD�&�G�I�^���|G^��6R-�U��8Q��
�t+�f���'�J�
�	��;.��ӲdU� L�][��ԋx��A�DT���h����Sun����0�5�S:���"Y�2������D�e!}c��&��pY�3w	.<6��jjq�uQ�G_�3��� �_� �~�n~v��]���|K1�R*ߦ��x1y�yjV����2��ז1�9%��0���F[;.�iϓ* � ��y�JK���Q��b��~�����/�ڹe��vs��I�l��O�O�a��>�}�uG�_�����2B��B�Qd9<�FV]e���j�e4@�����[ȴ�R�?�7a���,7ܢ �ݓ����?����2��b�y�"Z��$�Ε�B�"�B�5g�7�f a�\�R������u- b;T��A���C�lfn��f�ԃ��iuO	3\D�Q��%�
-��L�ez-�'jo+�p�/E;��5�a���S������w./S�ܶ#A4�%������ܴ�l�����0/hd�Q>�IQ�o�z٬�wx<n�q��w��c^4`��r7�7����=�2E�#�h�O��6�V(^��G�8�n(o�{�'3�3(����^`��1%?�`&��,+�����>UF*��F���Љ����sKVbXV6�X�X�N�wl�X�V�Q�QI�oN�-Cl�TdƏh�m���,:�P�`ኊ:-�I�8G�a�ؐ�tzB����U���s!�~M��(b7�t.
��KD	�E0WX2|���i���Wd�<i_�f皽��t�Q9���?���PXEن*&]/J8J��k$��J����&������>�� Q�p��SR �y+G?~��{<������x������$��l2Rү�G�DC�����@qcK��]ݖD�EZrW�
�WXFף��nC��K��������S�e1�P�@�;~d��m��+�g��UB m@�F����L�q�S�S�(d!�X�hת�q�{�霬�㹎Q��=fCKx8R�.Ƴ7Yz�yV�}�݁MS�x1mm�$W�_���"Y�V�z��	�m����=������F����+�rJ�k�I������g*)���0�������,���G{���I����(V��֔��|WN>��Qȓu��x:��L9+`��Ү��:�l?L�|��T�c,�cI�X:`�����p�pL� (�����Ġ����45�ޫ������l)s� �D^?��%1�PA�bs�t�f(b���U��wOָ���ܐRM,�6�H� ��tp xZ�;�V��f/�O-�6�L {��m���R�_��%lՙg��`%�؅���p�%��4�2�m��<���/2u(gm>�oeG�)mm���v<�1�X��DYt���w<B������|���Vo��3��@K˔o�[�
�&��w�I�<z%��#����y�]'���3U Ua�M-#�X��#Q`�z�ƣ����pD7�lQ�r�:H�/V0d�2/Hv/�S/�q	w��)s� ��?F��p|��-��29���!�� ߲��;j�U&(�Z��D���',n��Za�f�9�ݫ�0х�O%�������MlE6�&�M���+��~�[v�#���h=; "[�
��n���1�2��]T� �g5��B$��l�,y��6��H�Z�o���+KK� ^�d'�dC�a��ʣ2����B�f6���
Y4��1����̋<AV/�ؒt���V�R�
'vU����g�W�V}ʶ�t��%��lkۺ'm
��/���4I��\�����.:�c�BB�~0��q��,Ec�,�x��˱�p�1�����BZ`�?H���g;�Ҹ�/X�!&Y������ZX���zL�)l*�#�3�z�Q)S��MP�iR��3��
��}��	��L�|bx�u�UAA�U��|n�T�ρ����^�<���*�+%����!N:�Q��������b����y�D^]?��ȹܷ��}(�w��a��S~�yp�/��-��~-�6ԜH�G�[y�h��zsk��f�~�һb�r���eQk_8Z��+�K�/�H�ӣ.�x���*cxB���x��x���t�rʔ�`K�ц �Y��I���K�B�Wcs��
Xx�8�?�"U����x��`9��n��6�F�/&���1 F.���X�4M(P�V3�P�
��xg�;��@A���q�ּ�E:%CE�[��y6��H#J��m�}�b�D�Є�d��D}���+��͢�q��h{�LȪW�V�pu�kK)�ƧB�l����8�%�E��܆�~{n�:Pr������g�L�ܬ͉�-�Y==~f
�:ܘ�nE�������`� �9�EA#�8)%�)�>t�o�C_��(���=���<���F�8̒������ِ��-��0�!���
;�?�P���Ҳ�HBC�n�`k30HT�ྍ��6���Ȃq�����[�U6�����"HM.�� �ƭB�u7Q���'O-�/�@��7("<x7ԟb��}���J׮ͮ��O���`L���g[%�K�x8,>>����}��S��p��3R�S���� ;핥�-JV*�Ν�Y���������;ɻ����e�Y���Xaf�t��!��AhJ�Cռ�]f���^��ʷ�������'���,
�]��w�h�L@��.[��<Sh��L��ZLcF�������A�r�	`�|�/�8���'tp�$�@%��kMd��a���|(�KS^��|����qO
�K/�P�� �-`��;���K�V�\:�w"�=e�?4�j��Q8h��)Ul�cD��)/FY�I�E66�(H�r��4��*���*a��������`��	�W�Q��f��6�Ӹ��n<������<ZX������2P��t�V��yuI������E�)���
�Y�іa:��=��T��d���ꑼ��-��G�dîe�t���cU}�d	�I������"v���[#]QH�i��� F ��:�j/Ȩ��>S�rΖv�êG���_;�u�Ν#Y��}7;��#yN~�Z0�	��2(�@�Lդgҫ�˫��o��iԤ�&ښ8���"A�T<ezr^E��+��f��؛��Y����M�ד�����e�����JL6�>ա=���|��Bw������?����F��Z>���#Yܬ2$S���/�ÒXp\a��;g;��B�����B�����t�V<}��fK�&0��.ӤeuQ�U��;ڮ����p���3��h��+wY�D� �7Q�j����������g;�J,���B��S� @M���j��Z��Mog��W��f��Q	
�O'R��a�I�s�^4�jl�����mXz��[}Ԑ��b@~��}�RJ" ʯ��(�F���W����܎^�"c'r���`GC��,��|��.���ըAxʗ��������%�2�J9���~\�4��r����F1�+\=H�D~o�bh݇�$��$� ��ݷ�� g���,��D�e��>������?����0$���O��o:�*A�rN��z67������q�X�9>˄������U�sJ�d�vc��	Ig�ɢNPv��2Xd.�3/��u$���o�5굲��K���v ����~��;�Q�>��`���|�o��<��Xr5{�&���.��%0g|ض@�����hS�h�n����0%:����48�-E4E�S'Ed G�J!�d�
iu�c��i`:ǀ���]�D�s���(��^�Ӓ����ED}��)�=R��g��x��_x}3dK1�	ߠ��gXE����� �I��)��[�54-0X�dN"\��M �%x5����E8���Q{1�յ0R��:~�\�h!hͣ?M�Ws/��gD�g=řUbj�l�֛�U:�X�)F��q���_�Z��y�RL_�r�y�&�f���נ6&�3�$���s�:�:ҋ��.�H�k�xb2����e�?*��ں\�-�w}~���D��&~�F9 ur����a��
ˏ�/3��C8k��0�.��=�߮�$�8}��%�A��:!) �f��F�������Z�����^I���o��D�^&l���hǺϿV�K�!/m��KE�~�1tM���⡷�V�8FD�P��,���1�(ب^Z���sR����D��k���H�%}����~�O<��T�`��	�2��yv~J�`n���p:yON�������F8� (9�2�C��/������O�ZcӻQh5���"�(~�F�j6´	m���O��z{�Z��}�h�Q?�o�m�F�����>�C6D\�����%@���77���/O������֟,B{l�]*�t��@���F��ͨax*�
ޡ� z��e(�"q��1���e���FD���R!Z���	I� i�q�d�e_�k�%��E��m���^Beնω���M�9��ju'ʱ�����g�b�U���]B��>��r�p4����Z|;G~$"���S�x���S��n޷�H����$/{7��2߷�p�	���7lK��.��sN<��Kb4Z�4���"0�l��.���ޑ����%c��O�+f�� ��*5��/(~��&'���g7�|6���?m�$�����[�8S<�.AT� 2�z�q���g%1ev�m&�#j� ʓ�[k���(�J����e*�;.%2�
��_yx�Z��|�+Ll�����SpH����J��)�7Q�\T�N��D����p�~��I]E*5��o�zcS��
�W=��)��y�q�`�o���087�EV�D�U�w<���f#Č�h��� �LfFs����b�t��Gn�x�B�!��.`��� OI��:k�d6O���x֓�4�3�A��ٱ#�j�<7� ���7�����dw������D�5��l��n��s!�
u� x[x�L�پ������eK��ig��y�. ߐM�����z굖����OEe+�&~[Ҫ>m��ny�u�G/Tg+�o��lm�C�B��4뺿-��v��H��v�9��)��ŕ���N�>���K4i�X��+��4��h��Ծ)�����~�5�"Cr��WY�XWN��;-6t�Nb$���M�F~��ځP�E�}����I��2���Y��#�FP)��s#�����_i/g?��^ o���
@�̨������w�L�,p��+�ΣK�S��V�~��]npFw<	�ԋ�1�~�'��c��ňBŴ����C��O+ă�l�	���Q�i|�Qc�JD�7^�L�n�ђ�!�򟍰��Qr���{P;��?
XM�� +*`��'g�.�8X��Gp/5�x'���%�d�|�	X'����]x��H �S �(N��d�D���7EGl"�K�xȁ`b�E����#�P(7�5e�@�2p�|=_QA����K=�Z��!�v�O��f�)���_*���8wJ~Jp`n*08��-���W�q/�0�z��L��Ya�D��̈́��]�  ����a�Î1�cӮ�	~�E������{�[i���B=a?���>��]������2ޥ���ꔌ�y=��)�>�v,������V��t_�`�)S�$-�F�\��-�3�H���C���c��-���m|�$߰gD��ɉ]�>�("��9���d|H�Td�-&�lI��:������N[����#�	�g�Y(��p .��cYp��<��;��g3�F�:d�Ƀ�a��n~��,�o�B���G�>L�q��:�)!Z"�a��<���x'�/�ӳ����g�����1��w�:j�nPK�/8�
�s)6��`7:4��O�t����S)%�~e������"y5��N�����!�bε�j���'*f�M�{D�0�'����5���S=yD�,ŀẅ�=��g%GN�h1�&�^V��UH�ݮt�����_Ԛ�a���<1��;j�o�S�&W& *�>�cW��&�z���tU���
-�i��
���]�V4��.'�ib���m䫎t�J��K ���A���;�8wڀY0O��+jk�=Y�|�:�Nl������Nm�t��2��/���	lY� ��>��+KJ�����$^Bb~�v�f�U�O�T^#��a�!$��2F��K
�G��k��]�ٛ�5֍DA��±����9ւ�~�u�t	���絴3�z�D:{��<"j��
]B���+>#.w}W�*C�-WZu��)т�M|#"Vx�h��J��QIZ�����������s#/{�,��,�g��pZ�W�
Sj�P�f�;B�'��7-�W:�z5���3��l{{L��x����5�� ���U�u����l&oCI��a��]3�u��A}�V'�GC�u N���W!54��.�4�̈C?�#�e�J~.E}�<��n��R.9�U=?����B�8Kà�2J�v�UO�F�`7�����X�$�7b�d^�9[�bVOD�a+��X��CV�CK��R9Y�N���<Jl]���R�%��������T꧖�/gtK�6o�l��1�ͶF�2�Ӌ��Jx�'�c�%�5 ՅT��"�؎W��i.�p���X�=f�$�t~rS���Q���(�V��$l�|[ۣ�� n� :F>Zjћ�ZY8�4��0���|ȴ,(8���z�.�@���Z�LΘ�V��^��rV�=��P'�:�E�Y���pFg!=g�C�::�S5��<���Q�D:ݷ���
�H��Z� ��E��)��N#��ⓏLAʎv�e,�؁@�g"\�m�`fQ���{HК��OV���n�p%�b9�ˁ��~��f�{Oƫ씕��{=�.�7�U�~"9M�?{��pO�Zی��AF����*�k����!�u"QN6���N�a!�HeF��j�#���y�^y�Q{�[s@�k�
	��~5�H0C����H��*��fr��:W��9�2 sӚ��gJ��:���p��Va�����y�կN_�@:95��W�zt8y�{2E��./ڈ�w�b`�c��`��T�;�6�����]1�g�H^6��1�^�eW:ې�.�����F.a�-���O�
#),g\�p�7�����EJG�׮:t�Lř���FR%c�S.�z0�dT'Ҩ�`��{}�:��5)O��_!-#Z�_�͜tp�k���(�r'N5�&[�e�(�+ڤw�t.����$���SN�<��U�tJ-5/�_��jP��l1r#�����}�t�G�p�2c4���)���y��|\�u����8���%)�w���<�x[./d�.	HP�`_7��ߧc�����tŠ�aj��GG��ZNSw��U;��C�E��R�`R��-ڠ{g۠�Q�D6����jt�AT���x��,��!u���~�q�Mq���)���DL���s[2��.�����#��rzbO(sq���nX�"r�Rt.͘�Wuh�E�r�J��d��,�v���o���fҴI�5��qp�U�G�8�&��� NL�]ҋu�uD�j�h}�|��/��!SM�k(�,7G�r�9J������@
΂�v���o�h��?s����(sI�����Y<��Ϙ�V(Y6[��yMS�P��# �Z6��	ȸY��>���);�P�� }��a7��.)���In/�a�%���h?��G����3�����u^<1�C���j�3A��ܸ ��W�Gr�(�.�� ��o���kDO�ky�t��JD�C}��3�D��=S�y��X{:5/��w�o��Z�NCC�E��<0��JA^ޫ�6Y�4q�b�3�8��hh������=�#�]:�|mHP̀��l�<�\V�	']�-9!à~U�Wrn���	n��!f���������Wx^f��Bmd���@�}=��� r��%��ͼ�b��t��W}ÂW��4 >"��B24�gP0akG���a���ȑ/u����6t)i�Y��t�15�ԩ�׭\"� ���[����h���-e�V��*f��V5R�c����5S�/l mFG�b{g�Ex�tU-?�N�����ޠDg2�.�1�gxm)/#D�f�Z�/ۋZ�z�L^����v��m�6)g2D��Y0��8l��*�C�i�7��L�is;<l~S�gh�[ϰ�w/��>=�o�����}ؚ���Lƚ��h�7�IƼ)�2i�6 x��8��f�Iڕ��(S��[�+��M�Z�޻�ך�h��~�e4�޹��� g����Q�"��]?���4J#�+��ρ�Bޅ��@?'W]d�4Q�"�p̓U�.8E�ab͑�x�;&�����ܢO�;���{�״"^�%�Mg�n���T�m�p�rO�bם���3V��jT7�i���@��׌I�!y�!�z?pJ�30�Kѷ�m�� �	��R"���m|��Ϩ����	<[`��;-�d�.]�����bdU��s�C�G?�Y+^}[(��7�U�뢛>���~8ߊ1��g}o�b��[e�#k�b��7A
��p�,��L���L2È���!�t~jߟ_��5g�#�^]S#[|���B��S��?<�g���\#�a�@6�v�]��0��ْN��k��e��H3����G]Dam�C�&Q�+��T&8���W4R��ȱZ����N6��`D%(3{q�/c�8�gu�8J8-����*�l�4gx�_T_{Y�N�n�ӝ�&�gc����4�C/mB?��aB�v�H�u[�� QY���D���y�*˧��~��*�y���v�h:�JC��yoHA	��A=�R�]$�WC�u%BVyRp�p{�G��奇�6X�(&E�%e�ś9�A�l�_��vƒ_�v����jH�}�!M���cvQ���l4�=C5�fY����U�Fe�y	������(�'Xy9�Mgf׉jF���%�����T�u�oPg�``%����4�Y�l������QsR�>�^Կ(
m-GcL��뜝��lw����ނS�w���dB�Ӱ���6cO��MhJ�i��n��>�9����P��٩�1�w�ʢ��C���������=���HP��g�ق��nTs��&��a�������$8ۜ��=<��W�(B�g�6�=Co'��+����{)YÝz]�H )���2����H���YV��W���G`�}I�Xf��H߬�9-n'��U�*�vs��Y3�!�(�J��k2,>=�pڞ��zX��C�&xP�Q��nb�a�Ò��ޅ��kL|���,nҚ#���ҩO����S���i�ވ퀃�;���%�IU��p[����-�g>�Ztl{[F����Z۩�qP��j/�)�ގUQ���&�����b˂Y���=�$\y)��E����4l�AÓN�].|� �F��?�笻�?���,�q����p1x��ӆ�mOmNh�Ws��u.�L�aĬ�!�d>6L�&�u�B3-���sJ}y]��Ӌ�9�{p�3}�c�]	<��//�����@��{�P�A���:>�I���㎗6�>�����C�"2�!����Q��.n#Ra>�G3bC��_��E`c��a���@Y��$LwA�ݠ���aU���&�F`d@n"Xʲ�s�#7S��+ܞ%ǫ'��N��pP������TV{�~U �A�#���x�=lLE�C��G��J���1��!�ZFc��kEy���?�Ɣ�U�����@:r�5��iA�P���33A��-�7+�r0u[P36��Ū
uiy��fl"�3��g]W7#��[��C̹̙�4��Ɂ��d��>���R�w�wlL�ͱ�-H�xv
�PV��ea]'�u���Hч�W;�ҾS6�2eE�)�JVcɚA	PԴOf�D�Z5�7����������d�0`��!d�*1��5p6���X<c{t�7���$s����0�8�q&�*S�{=&������$�
gz�������oPJyɑGRu�y��xH��c&�*y���z��؟3"��1܊}�"7$R冁*R[D�8�C2Љ�w��1	��p��h��~O��������'xM��0{c)����%��?�	��o���Q<O��A��`�x��+ݓWD�k��?|D��m\�L�;~����*[Q��f���o���x{H��WyQ�H����=?Ҏ5 ������ #�
�@?������n���a-L����--��#z�h��k�	j����x-G
<gMf���N ��(��7)SŴ�ǭfTR\�lMs�A"���������Zb�R�[�]���'�E	" �[
n�3��ّ�J�q��q_��@��h�z�bK�Mr���؉�}�ў}���<挗��SQ��ԤU�֒�JQ��]�c���>��if+��/#��Vc;�~�.E�'����VtBg�|B���?A'01���䲯��4�n�՗3d��9��%x�)��q�*I��i�{:=2Ɓ����{n�)R�l��d�%�*;y/Se��>�
)���`�",�
u������<%8P��"h&��Eo�%���`�@�5���Q^54WS�)�  �7�]�H����[U���9�#���Y�nUD�KrR�=��$}�p�Sh˾�r-�mb��s�����R^���5���=.���%؅K�pl�!���*}�#O:����-�� ����6�V"���Xt ,Y\&��0d����9�4ڐd�Y�z)�2]��1����K|�x��܈EJ��4���Wc�=�p��G�"�!p�D�T��R�9��8Ɩ���u9��v5�P/����yĈ�P$8���x]���,����\���L�}�T�z�)��0���@�+Z�RӃ� �\�
Z�j�	��J��|>r�l���`(X�뤭[��lu���Cx��J�/��������ё��T�2�V${Ӗ���v��[@^�UޜV ǟ�>�-���|n�0 "4�dw@h��]Ҭ�F�uL�d���g`�^��쩖SL�J[Xg��!�u������O�h��1���J~��)�}4%e��ʫf��	�]�F-+� +:����0��:I��}�$���������J�����,I&t���v�������`�F�h���f�$u���0��g&B5*�r��]�͐�M�$[��tϐ�/�<Mp$�bw�r��"��_��`��B���J+�Fw�
Z�-���x��	��[���7N\&�E;W����͘b��a���G}���/-3��nP���]�����	Ř�fd��������D��H�3�>�3�+`�PD58	� ��%�]%>��YL�oy�@����)$E��-hn�2v��8b�MIdKe����ޡ0�!f��B5E���J`��������j�����wӊ�Nᮆ�H��u%�O�"�_ͫ��}O4���.��y�Z�x����"�*͚��?N��=�O3-�)>��tV���0�0��ˎ)��^��O��έ�}ѿ;^Qi,��c�;�
O�h�ɒ�I�ֹO��wFeܩsd6�3f�}`M��L�%�vR�ڼf�*a���f�+C��+nr�N����"n1<�rL��'�������*J�X���Ņ�&�*Σ}��,�~�!(��G?v�/F.�ՏQ�6������J	��������[����:9�@@�9q�r���4΄�Y<Qa	=���or��ث����*Q�j�gd�4}ʍ`h�=~*�Z���fz� :��|�����ۉuT���mE�1��u��E�	��%�4+�ш�X�+m[�XR�}'H��G{��z=Xm��N�����ia
�Õ*�^�&�ab���x焩+��"i%6�KC*���@qGs�n�B���t�(����ՂM�wP�q1Ú�J���,~@#���L�KOZ�����9��0b�����ꯒgJ4�H�B2�y�F~�۽���ԥG�$=�@S�ӊ�`�Y���++"�&��N�U�Jp,H��2^0�����ơ�u�C:d��h �V����$���s�l5�k ��|'�D�6��Re#J3ޫV�NI�F������]'��(ڳܣ�rio�������-�6N�_I�.X/�!lj!7��D�w�{�<ޛ᪩6�����e��'��j�z�Pt��Y����]�Y��B�&���x��o����[a,��n�e�;������6��B>Ԡ"�c�`[)#R��"��Q�r��Ӳ�k�q���~���M9�}��Ĩ��-��xf�}z���7܏W� #p�[O ��iH����ݜ�2�vF�����ޑ̨_�-�Xl��� 4"�x�}�+�V(ƤWH�B�ᲁ
X�'���_ ۉ.�H��E�	�Z-]ƻ�9p�!%qW��eqQ������A�3�h�:\���/�������G��6*e����[r���'1'�55�ÌQN�� XRC�G8�d��(���x���Pv#h5c��P>gX�6� ����Y�a'MګN�d�E�+�)@�n)ŁW�)�0{2^���a�B`�����?n$�"�K�sY9.P�K��3�R7>Nʊ��l��J�4I^�'k,���S�꤯%��5_��֡�u���H�Ý}cC9��e�V� �@���
M�(�ͳ���q�"C�Vx�*���%R�zlW�6z�V�<,���rL�v���h�{�%��C!���t��Ӳ�c_�Ƿ�?TM����)y�l/r4,DdqƮr	�En�ˆk��ñc��uݸ���ǅ胗��v�[����4C�@\����W� ��� n��P��y ߝH�Z.��^2��_�@�ӲΚĲ�:x�{�ī���@���sٽ��� �)7�i���*]���)���_��"CZ���`�P��`N��U�.g�������'���GԌ9�@�Y���&>.�u�f�}Lbl ^�:����&����O/k�,�p��dT�6H9%1�����OO�8}ߤ�����T�kt���"��gn�2�O~��з=��6���YgP9�cD�
_��e I���B�Fw%�u@������E�۰|�<������[��@����\~D	��Yc�3ʹ��s�d��7A)�X����OC�d?F]P�	����-������d�|�
��rt4�U�^��y�~8�|t"�8Sȓ��9MO��U.����+48	ǟ���8bRR3SAp꼊=E��*dRo�8<�/�,B4���i9<��፪=z��Ih���T��Tȳ�A���.N�kR.�0A�}�o޽���N�S1V�l��P�h-�ZIw���[�t�4�d� e���p������qr���/ҪܖV����xH]�晉6�	@!b��`i\���s���� �_m@W\g0�%���t:#j��n*�g��C�V���]PN�*I-�=yj�%p~V����+�l[����+'���ma֍vH�;Y`�Ǒ�)�-O"��\�濙NPi�ܾ�=��$��k�L�fB�f�輰��!dT��$���4|,Hs[����	V�=��ŭ��72p�d��ơ��hsP�3�AH��<\��&AdF$s2�|>Ă��{�ս�p�a�,�"K�5�8��@E��\*,<vs�JK7�>��<�v�֞(�aRZ�v���~�\��1N��``��d&����6Esk3�����Dn����k3��k��)Z�9��M��C"��Av7�s���GN�)z��"�8@N`��/�G������Gy��OP���v��_s8]#躑� %\�6L�\��O�����F�"j}s�Ȣ�9ń�ȡO�c�?�?Fu���K�H�n7��Pm����Y"U��|�x�9 ��Ê{u���T�m��.��hhި�o����|�����ǡ�@*�04� E�_�Y ű>���S�dË@˩�S:G�(�7�1��I�����q6�=��n��������U�>o}���2��y a����O���Ѷ�����r�Tu4�uHul�\�j���1�?�`�zuq�#G&�7E EwB��1�e��)U���������o5g����ѩ���z��.�I�pb�8I"!�d�h���z$^|�|���D ������o�<���_&=`o�L��-^���m���O���j� ����%&?��	� ��E�nןR�7_������y�tg��K*�G!*!�SKZ��֚{��q�m�-�.q��/9�*��`��o�5�kq���=E �_�TF�N�&5/��+�&�_����=�I�R��%�LP�=k�����9:G�eD{VM`aZ�:9Q�'׌V�y}?�d}���Ҍ��_ɐ4�]�����%�ц�;3�w�H]���{��?�;rrƘAǁBp�+��{�VkZ���С~Z�t���%`A���\���ܐ�Do�M%��.Ǵh/	tGi�f\��Ю��!;FlO�1�%�#I�O>�鄭jX:I�4R���B��r�Y�OS�Mځ�w:�����������DѴ��	����Z�O�^�~�޲;��<�@X��D�'�ؚ�7,(�X�l���˶ȯ����kFj ��Q��