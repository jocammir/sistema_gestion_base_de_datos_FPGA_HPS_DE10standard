��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0����_���3���eĭ)|u��XXp�qPb�.��Zp�KC4��:�-y��y�Q}��B�+6Z��yF��; s���I��4+��.D������az;�7��2�{��6��}�,K3�өLʱ�Q�|H��pZ��|�Z��c�<��`�\Li2!oCX,��Y�QV~kL����+k��A+1s�>�pf�����/Q��i��x��֑��Q���u��OU���I+ޞ��@hmghK.�P��9�@�|W@�3Y�8���A{21�I�j���(h� �h�F[���f�u��.T�s�s�Dƽ�f�#�t�V�y��,�^?���}Wrc�	�9Pac�H�4�T6����p�M���}��K 2�N�"v	`��%�%�J�6��6\��`PF��%���/q��q;Q_K�T��-��	��Bq|Pq��)d[o�~��RwN%�#��.x�l��ld�"
�.S2O�7��G���$J���s�:fͭ,��K�M��	�%s�lc�D�	� �{9[i�,#�RS����a�D�����`�F�˪C�T+����%�Ś�4$Nϡ���Q��]%?���q^@�>a,���B����_��6�猴� h�����]M5ޗ�K��0K&��LE�Qm{�	�aV��R����u����(D����o)\o�����7��#&w�o�H�P/<Ú����?��[�a��~J�F��o��j8�V-!���q��k��\q���ʰKh������teZl�,u({��n{���фƕn��m�P����4��"1��"�t�i[�vrȕMeT,|Y�4WP��m�Z��1K��Rj��-O�ql��<�A-�K�P�&{��G�����T��o��DͿ���
&C�,,�?Bee��D[���Q�K�<L��.Ǎ����=|�ܜ�P.�9���~�Ih=���+�"�>�����ǳ��v�H�S��ϧR�Å��Y��/���Ľȫ�7]��R��9�Z�\�Vj~��g؈�\  �kn��.8&�������7��/���W�#K�k�t��;�w��*�� Qe۹�.����Y_��}�!l��2<`"��B�=���3�+�$�\%�'��49Ţ蕭��zh?���>��ݾJS*�h�L�A��Դ��;Ղxճ��>d�s��k�6��Ɖ��\�U�՝T�z`b�څJ��B�TW��WQ�LN���x�l| ���dR�=K��JwB�n�=�y�����G��v�����;XLҲ��y�ۓ�-��p��F�廀�X����b�PpS���w��uY-����3쿮�1J�M�ず}��Vd�'o�o�DU������e ���(�B~�m���D��X��oO�j���CC(O=^��k6���[�%ѷwI����[�z�Hv<o-�èO9V��� R^�3>��<�󃣋4�LE�AE��!��_b�0V�������v�j����z�)�f�M�ȯ:b��QiC�C/�K��r!'Y����o�wpp�v'�g� @e��D�?���m�/�����f^b���c�b�v[�Gh�cX�ac�|��x8�7HN��Z��0� K ��jU"]�>�_p��EQ0N+N���pz �<5�������(Gs�c~U5X'7֒@�R��P��5�ұG8�1���ߞm6���XE\� 2�{���g��35��b�o�1����o��!߯a���z�ĥ�ń4i}��Ԇy�N��G�"��ȇk�$��5g�7!!z���B3����O����k����+���s��;-���ه�9�N�1�YP7��/̬pP1ό�t<Vř���+^� ~�.Ėh-}?��T5}�M�;�V��P!]