��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��Nڭ�	�����B�#Z���?�4�j��0�ΐz�A�y�[��I4�fB���_Ɛ���-����B���M'~��k,���'zf���]A�� -̭���ҧ���D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T��P�]��h�� �x��ϝ�BQ�H��B#0P�s7�D�l�������Tct�0��{meMR�p�R5��.�6�F����&H+W:��G�]'���c.�����ɝ�5�����2���5����TG���9V?�zu���s�{u6Ֆ�ɽ1��0Sp�O��l�����-N3����[�3F|H�Nr!��.ҺE���7a³?���^&P?�j�]��[5P�9W{@mKe�󀽳u GӰ�^VB�ZiJ"ӟ�µhv���Ռ��ɠ&��֝��М6T��!�1�tU>��b*:bJ���y���"f����xq6�)�J$`Ņ_l����5qƙ����j���4(E�`���4�0^^ߎɰ�|d<K�6~β&�6,�'|�9n)R�~���j�d�8$��n��M:��i���߈e��-��''!�U]@ͷ7����xmd������Z��2#�U��Z?��;E+?�1�Ĕ�*6Y���Z���f9��޾�>�n������[[��D��}G�I�J:�#�.K
m��J�>��(7_��Adt,�H�6����2�U�-mH>�״����M�P��x��3޾���8�<�d��|בlq,.�ڇ��ţ�/�����Eo8%��KUl�^gUb�j������Й���}Ǡ�)S�T� 	z��O8�������&���K2����vyD�$�t�0�����f��P	�;Xbj��	�~VM����D_[�{+Um�[[�y��U��t���b�E-����eN1&�q3۩Q����t#��N�~;7��Q�b'W?��!�Ϛ���U���t��({�(�7�����n�ox�dE��Yr���莨i�5Q���w�U뙈-���K}4�E�0��	q���F�k�6v����6X>��*�_����|*�v��(�zcY>ϟ0��x�V����4>s��?"\���9 ���+>A�Kȹ�[�,���������ހ{r�&@��$�_�d"<B�ޭ���}���?��Qc��I���R��g�;�U�n�c�k�E>
�K�
Y^\��;�f�1r]PK.�< ��Z_6<}���3ǹ�Y�`ۦ���&�j��I�݅�x�3��*�`8~��c��6�%η
���Ox	g}���b~���a�_^�6�Uz�5���Ԟ�eo��鏉�<��c�Q/!X�	���k=j%����J��t���S�VO����<�;��$��*�+�g^+֦���H�[�Цz�l��IlE�$���S�̍����U�7p8O�>�u=Rg��� 權gG�A q�{��8��IT���n+.�YA��o���0���ߕ+/߈�]��G�Е�K��U�'c��L	e�r�j��*R@K�[����`�py��'r�e���ʜ����7l���������aѾ���X�DV���rҿ���������4-�����Z�O��lu��ޗ��^���K�̴(�%�m3e�ΛVC�a�M��1�Շ�e~.�JTw1�^�atڕ,*E��du�&0�Q����+�%FӿRȗeUʴN�3T� �u4��\�O�G��3Sq��	�r��F��5QoL S�M���`J�K#��t���1���x<PV!��^��g�K�4�n������ʴ;���%ڔ���W6Xca?�zY5`�����tzJ=e�M	M�Z��`H���'�� ���\�����Ϝ"�SQ�B�����;�zԙ3��P񕩻U	"l�O�a����(��"�D�zu� �%t](kj}I��z\��ll�H���d���8:�y��??3ye:f��j)}�Wk�SH88��B��}���6�h>�Y�/��7���vG�h���o#2�� l�ylއ��礀�N4#&�� � O�
L+��]����)��':=a�<ß�u1��GcIꢂ�%(ר�\��F@����|)�dD��`�\]�}S{��(���&���i�%��ZpIQ6Xe��xk�|0��`��ץX��.{������3�bώ�]�#RҐ�W�]!X����\�z����l�f�û���W��H�B?(@pJ����{�:��8{��Y���
��}�lׁ�nH��l|#<I�YH�6ɳ��({�+&a�yx��g�+��w��Q�r�c ��6g3S��q0�M�%G�韗���)�4�"-�I���4ψ�5ס�}�y_�#�y��7#Nk(�R��[e�X��(Kuڦ2Ogv�ߞ����~챳����h�
4�g�B��]���V#�_�8�����iޛ� �mEr 5&���M�V*5Ai�W#�w��a�4��S1�nڃ�Z!YĨU�:�Ȼ���j���ܐJ�F29�����ټ#b�iU�#|^"�5_?�VY�jKE��`�}(W��������e�H��F*����d79�3��s���g�\�h�X ڤgl���L{L���������ZjV�c�f�,k,���8xQ3
f���e��~�۱�GB�ߺ�c�����f�tw@��L3IKq��� �}�MV�]Pҕ:
��vo?�H�N�<d��:��.�L���o�|��J1���~�E� ��(�4����!��� ��EE2{Q$���ݦ�"���P��+Swx�)-�������b�2@��ع��8��>/1g�ٔ+cCQ��AHX_���$&a?N�?��';Ԟ.Icr��S�]��R�HT~�����ٵ#Y������ygg��4ކ,*�H�����-`ٱ>�i���O�l{TV�fn|<l��]�%�	|3�;�Rv-����9��q��U��	���K 5���Jlrz^� Oi����?Cred�STq�IU\��D�3�H�"v�3�\� �y��!�<�_�mB%�P������9���΢X(��U��t+pF��k�]#�C2O����q��D��%����i�
7��º��Y�	k|�������Q)��廲<0mP��ڹ5��aQ��҉8}����[����/v�ܪlV֖޿@fe�ƭi�A
 �FVU�.@�����|�`���lh��a0�~Pe��f;O����&+?4��ٛ&���w9���� aܽ}43�'�BwvA_Pl|%��2�#�G�&3�i�ܐ\��+�*'upg�\��.bj�j���
�_7h�������^B�!k��h�~D���U�`�N��!6-��cx�Ö*��aRu��2�i��u(�;8+@�ǝS���1�	�8hM��L?W�z9����x��Դ�!`Z&tG��v�DLn����%7O]7��h��q�b��u�Zۼ��3N���a�e%�~����99���� �]0�Z5N��ݷ��t͓ot��̬n�!���>���#�K���2�
���ކ���R=��uO�.=i\0V��-���NC:/Z\�����I�$��_RSi=��U˒��ޫc���}_!Ud��ne�O���-�i���]C�Ȏ��a�G��噏1v�T��~m�!IW�°������I������'�����~���1|ܛ'��/v,U_����J�U+Z
�v�'�R$�#ĥ��d:���_�^�LF"���bSM��\����2M
���m��L�H�'�w28;{ i���"�f���z5�U3a>"�N.�E]���F¡3�H8�+Q���)��r�ѡEsp��&f�ܣ��v9��|H���|�p���˙��F�3�b���4�>a�7[b�my��&|T�X|Jnit��.-���M^�E��Gj_���$˥��Uٺp�C�� ����Y����H�|��&	�ѥQl�v�s�Fw��,E�l١գ�3Q�#��	����Ǡ@�0˱�)��t�a_mv���~�0x�B|�0� 6���à[�Ӗ�"�םHP>�� kFz�+8��Β��=��ᮘȆzI�Ko�4�Ez��~����P�qpQ�'@sl��O,�>	s�d�K�y<��P�4����+٨�e�nm���ʀ}����|�Q��j�H�gm��?C�k�IY�g�1Q�:�"��ߩ�b�l5Kv�'��c.��72S�GE҃k�͘Nbم�n�M�� .wauP��p���^0>��J[���)zt�)#���;ou2!g;}���w�jo!���QgbC>r�=+��s��Y����&E��GC�+=���#��w����ᵒ(�%O�G��/�Cs���VD����7����Ȥ
����ݥ�L�]��`O�l��}�*� ���FR�hCN�^+c��@���q�]�)�K?�b�h"�����a��a��[��Q�#n	��'k���[���U��*nI�$���gv�X)r�O������h��a�Q�����#,�ͅ�;}x�O'#� �.@�*��$�Rc���b"|U�]�K�3�:�*2�F�QT�,������
���`��K,��m���c®��Z�B���� �����:ielj��m������=��r~�e�����v�O�� �(m,O��4PK��9�jǛ��5�B�_*��d4�P����3jBgG�/�8~���H�P��(ۋ�� �Л��_<l���Fe'�(q��E}z��[�'�y�ř��>1	���\)�I�iB_��잣���*А�tS�n�cGH9�|4����J���7��t�e�L`�I����@�ƶ�"�2��N�ۃ�8X֨�ŴI hN��B��>��^]����{2��Y���P���dm���eEh�Ƌb	J�\P��e�ÿ��cǽ���EWk���O���IJ��ɼ�J��E��ABi��5���O�l3E���X��>[R��Sꑎ���G^�Ĺ0��>�T�R�\^�h��xc�r�m��F
`�ՙr�iE�`��2�Ay��k�{u���s��Ǉ���#=]/0x(��O�0��!��1*��Z@[����.�+X!a�>�(9�A�΍�ݾ_�OI$��E���<�¢�g�>\���J��L��3�z0�R� ���
��<!_���[�K�ԗ���=o4��,	FK������ �%����׼t®cѦ�>o��dW �qb�%M�o#
@(1EH�2O��[����>�@t4���I�`�'��"���D%��~V�_�ʡ�����_�f���o�WJ���>�}�2?���I���,��0�g^�nyI���~��_�W�=�dA'�T�W�u\�n�V�Q�b���꠆:9T�7�?��Fe{���>��ԣr~��)ť�?C�[�j3��䢻��o�Sj;��=DJ�M�y������y��k��D�zn���˰?���j�;Y��o'�՘�\�ʱ�2S�V�v�*N�?6P��id���1`����:�_W��;B�LoE��P
�"��4��Ѧ;��% 	s4Ǫ��7�5� MWS��uIaw���u�c�\��Gg�v`�a���hQe�
&�27��<��:?�\�0�Q�b���]��m�ı���V4N/�D�O�ْ�ʾ���KY����Rぴ��m�Ώ~�q,�S��L6	��r�ل�w��C(��Q��M�V�hs���ڧ�s�R4V��mK����/�.�s�,(|�&_�(��L��g��D�����na8�xRa�AN�b����:��cř?�kr�{wd���O��t��,�b�`�]�I�<_fl�F�dW�� hQO���$����6�x���$�l�OA-NX�gc��YJZ��������P�[Q�|�rF$�}s�6���iw2�)���,�@ �A��ڽ��E��x��]$%�ǗK�b5d�"q��^#����\'��/I+�XT/�/b����tm!Fa$;Qt,�ۇ)�1QCm��<GP����@"�Ȳ��MR0�1��	|FM�2V�sY�S��R5S��>��b�6@I��O�v����4���W�=o���{V�t�8-�<�]z+�<~�@�T�.�`Jg}*PM�zB2�������3�Ͻ��]]S1/������ᥒ���H9#E�j��
V��>��l��Q�;�/� ^�ׇa�� ZT9$�*�8��nK�q�Q�@�}q�ˈ��"������@��~T^���\����<+g6�F6	u3��o5��O%L'r�������q{�3G��piK윿Q���z�6�������@]���&w���m���6�E.�g�/��� q�9�գ�Z*\>dl5�4��^�p�t���/�[a�#k���hhP��|b���u�z�|�`�0�������ϩt�S&V�tx7%����8��P�Z�&w���,�D�d �̧+�l�~~1�ʉ^X;v�-�68�	/��ef]��B<���H��{K��.�E�H���B�ә�� �˖o�!*{��P\?�Qُûy@�"7�p�ci9�(ɧ2�v�S�R{!��_0��7�h�a�0���X�4�%�RG;�;�֘�Z��#��1�M��ؔ�F9u�ǚ����M�t��R�)NDf[��x��1�Zƽk��
& �E�#ݴ��s ˕:	 J_J.�/(�*Ԑߕ�����u���8{����İ#������G�u�]�����JVF:yF�j.�[EDۨ0�,� ��1�T� T8t��l�
��� �=���6 ԝ�d��V�w��<~m�\FF4�"�ᗇ[�:�Sb
,I��F-�����7��ޭH��z+����x�qy����}3#F���+%�OT^���y/:���,�TuyQ��Ӡ�p���bRei�_�T|��(_QԬ�r��֬\���+L1�:�(k�I{� � ����m@+k��A=X�������9I>Ru�����im�}z��H��}��eF:�ܚ�0���P}X���ReW�8��`44W�C�&0۫|%ZS8؛��S���/�̝�lr<f'� �i�s��>��Om��M̰��%��;��ٻ����D�����/V[�7��]hwuFC�(�x�#޻�.ϤG�M�B���=��2H�����@�#���Ch�_�J�d�x ����E�9�&r��	������K\�N���fu/�)��ؖ��Y��=?��%�6�A*������H����. �z�E��i��0;��i�n�DN����֙f��T��Ɓ�'*�k��
�z�*v���v��4
۴�/}�WC��U� t�{�)���H����C|���,P��؆���������7�G��25�Zs@��1g�$�X�����A�)�h�U�*Zة�̘y��il,A{���B	e,�ͼ�zz�о��Lb�I�'#��D�;)/o�;��e۽d�&b�#�E�\�flK���0��m'e�h��;ߑ��R���=Lh�	}��R�C�h�0<VɃ�IF�\����#٬]/9&$~w(Jю�f3�M�}�&q���̄�䲒����Yi�$����J��K/��=���5��M�06���3�J�UrȬ�����<S��N�{%����G��6�ь�&�c����'�oXb�����,4�j^���`���r��(��a줢Y� ���XO��jj�c�
Z�;�౐� S���^��mG��3��s�y����ƙ*��g�2��FbT���%C��GU���jJ�h4��s�(7�l�����mr���E�z�~G��S뿿�s-��_0rxqI;�ϫ��6c����N������U׬[ ���rv�{�ee=N� �@/!ܯ�(��1��~u���&���""L#�X��][�1���Ђ��HM�ާ�P=���rnDo�3�?��ŰU�N�b�6K�W�T���Dp���SB퇴�l�z�d(�rT�x5��l9�+���!�Ż�8
�ͨ����)ϵ�����j�e�J>5#��j6!��(�<!k��9+W���.~����`�N��E��W��n��5��p��R*ޣ�>�h��nzH�%�b$!�G��5_p,��F��)�֩	H���.x��ݻ���V�8n���W	����%�	��\�ݎ��̤�"[��o{�u�.�h���y����"M
�Oa���"�+ �gЧs���+�٬9�4� �?��v��s�'�W���-w<�6�%��u!%��S�7O6K�cx�ŧVD􃢗w���Ό*?>�m���)�ʘ'��}�/��0B��9A����~��Eٳ�V�
�A�2��5�㺕�\�p���ش�Z��É�Z(�	t]� ���[p7	(��7�4���Q��3�a���.��v�J�$ti>��
0�y�1�����p�)�l�o~t���s ��N�=��G~�0]�&s��}��'��?7��3�_ǭ/�V�[�5W�66?��(�@����"
�|��	ʛ�7�o	����O6vl<�7����ZZ	v
u=��EO^m��2�y�~�����莗���7J=v�� �rE����Ì>��Ð�`d��O��_ӏ�پ�t�R�ԣ%��kh�xMPog�f�P�̫�j�(��,Y�I~�us,�Y���<ס��GDs����N����#e���Z��]�1��+�t�B���!�'��x�E�Υ��e@cv�A	렩L���L��N�n�����/�5tX;_�T+��u�@d����Vj��5�TQa��G�������l�9�C���>�P���֪A4�P�p�
�(��7����=���RW���&/���d%�3i�o��ٶe>XF��|�-���e��Ji�C>JH��{���8�#�8(�h����P��q�P����K�y%)	�w���Z7a<ާV��tt�k՝c�*��QU�j�����)�˳r��/`�V)��׍嵯�������؊�3�8���aA�� ��\1噉p��?޶ab~RR9��t�q������M����U^����^
��P<p�9��ƨ��"tl�/z`�{�zY|����V��B.Ʌv�5����t��B� �̇T3I�X�s��r���`O�m��^g4R���Q����۸5�T�'��dx!��E��������l���P);l���������x�_+^�]a��$<��[�N���i}�;S�QE���ї��H�q�K�2 N^hY�r�;��K&��1�J�����M��:��ᡴ�[_E�s�!p�Y�X^k5_�[��P�m���c�x6��)w�V�٬�3�Y�W�6�J�+52xww^f�H��z�g���&����*�����1��c��XI_�L<�c��������bx�ݦ���rGt���J꟟��9�Dcn-�nD��ѭ�;�����?$�be�*��2��炨���0*�����s4"x����?!,���f��{�Nh�]���B��A+i3�
p��'i�y��$M�eC���h���O�RkAgt�n
�'��sv���%�\��魍�=p�D�o��E9��瀊j�{V�h�J�>�vH����:˂��A�I�1'�GZ{w`�e����O�סGC���b�cl�u��E�$'��}Қ�5i�ءR����e��p��Bi�� G����Z�]�:3�;W^">SN���Q�[t�\J��Vv�jE�@����P9�����w(0%񀺐�2c�L�[��(��9!ѳRŋrĲc!���iZ�xd#�������̚�SB��_�!6�y���= 5���2!�����=x9@���fN�����{�L)�t��t�ρ�eE��,m�T��D&YE���ñ)�X��f)�<f~���:���7�,p�A����c^��'\�����nɸ�DJ} k�U�>= ��A:�	�����D�"����OϢ=��q`�C^|S�Ƹ�_ _z�j�>�O���Rs�X,l��<}꫅�󋳉��T�$n{�K~cd�l7���z��46��T�v��#�e�y <�]��Y�H"�č�
*�gh��|/Ok�޳ ��j'\]����νc&s����#{:8�&(|#g�f=UM�I�����Pn�P��1�6A����ȶ�&:��z��;��X��`��2�q^#��p��m$d��@/��a�_�t�K�����#+'�D3���`2p�3!�^���c?�W�7q�
op���#�A��M|��a�c�	�2*�.���xfy����걫^=�6��d�6)'��2>�@}�f*AP�v����g�K�]$<s��4YFs�@��I�`��b*�0[V�Ũ�c��6|�4Lt~qTz;'�ĕ	�֘Bű3�S�|�X�]%�`w.9�	F7%Y���4����޸@��f�{��Ԣ�ԯ��W���	4�%��N� ɼ�M!:gM������)<�L������%����/;��s�`����B�c6C;>aG��h�Krx8!��s��M��`����g^#���K��f�<m�w�8U	�e��0t5w����Pt����/-��}G����0hN�33b
�{�t�D8��k!��3��!�ΝH�.W��%��V��e��Pr�ٯX\	u
BY5�9z������1]>�f�~Q�sb$�Ŗ'^�{,vu+���ls��;����d#+	:���rޛ���ϐH?�9�V�ʩN��i��/ᥓ�90f?�%Ǐ��^�f�U���ڌ���)��]��B|X��ȐS��g���ό���P�(8�$N�_�X�~������&)��8᭙#QB֛}��v�Z�ș�O$w�Sv�r����$���L�M��ߣ�A�M�*�N}_&S`�ųJ��$-
XU��ڼ�ы�?"���{�,�r��Iե��dK��B����Qj��v����VLK���TZ�=F����靌�+n;������\lω�=(]�z�8�ܠ���%5�Ɔ��\ �M�Q�#Z��{���<]��P��C�nT�Ga	^}��xV��'��`�Z�DeV� ]�o�f	��.s�a��׮a���U����d��.��80^�o�We��
�r�.����`����y[�G�I�*t����}a�w�!M���nX(��g&V��`�l6W@x��ꬻ��������D�3}���0�ՂeǖDC���r����H;W��յ~bXM��,M�u�����ٺJ�H'3����:I��#���?"#.�f�gB�c�kO!D��pΰݍ�P༬F�³��67�U�D;R�|�_�s�(��Ά�����	y�H��2z�NE�\������\k�pN8��g�uE��?���v�"i�ݕ(�	a0��d��Q���:Y�Aֻ~uU�� �k����X8֪~w�CL�)s��-��ױ�n6[XțI���kK���U+/�k'|����#8~F����No�W��������
���sz�7t���y+�hL�P�ى���n9�#]n�wA��{&���Y�����E^np�u�m��{ X�)_ې8=9w��ϧ}<�s#r�nn-wA.�d�]D��j�.o~<�A�H5�%(�ԡ��{;3��|�XL)�4������\W�%�����t��Rc�\_��	/`(���BWG�6�Hԍ��8�$9��?_qk�b��!�s7$���x�A�� ��j���A)��t����5>qX�,1�DL1��W)8��mSŷ{Y=��9�²��a�	>���xI��I����,:_�S�[�+��z7�����AT�%�l�f�uf�`���zJ��]8��$����`E�h�c�]�f��`�W�v���҈S�:?{%T0�N��}I�\aoǚj;��o�Ew����O�p߳"��i�ﹸk�͔6���:ܽ�n~�q���>+`�\��/����z�;��0^�����4�����<ܱ���a�9����w]�]&�1��O��b{��u$a8���ٷ��9͍�,��4/����zą 0{�����&�t8x����Z3��-�8���`Wҗ��FX��sA��p�.��҃��=�t���*���4�7k�a��I���I�!�������O}�²Ȥ�;~�����*W�����l@&�7��ۉ���}Qo�`TgB6[�үZ�cp�w>�*u?�	y�^h�P�������ԗQ��MDʀ��TWʆp���t= ����FL���<&p(���n�%���0�l�D"_q/E���6m���!�Jcd��b�4���^@Y��2�$�dl�FO�/q^y���PH��h����A��b��ȿ�z���X�.��,��j�x�����rA�3��@!xB�n��A7q�7襴f�i�0�Eg�`jE5��.!�8X�yuIZ�$@���4��m6�ueZ:F�M�GӘ��g� ��l�� s��M�`���p<~Hݧ��$�uH�Q��/=�宷w�s\�r��b�yv�_�f���ؠ'x|�g}t�4A�)|�t��;쭀�%d�b�ٔ[�t�����$�!��,�}�i��G�A��D!��?�Y0+��HSs�)����	�XVv���Xv���W�G��q����ҐJ+�nBF$T��#��P�B6��7I3gÀq���iݎ�ۗ�^&q�:`����+��Dmk,��.%is%U�.��4 ,���d+(��V���8	`6� "�����ȂS� |�+��|��o{���V�7>fuw��~��l�f~�D^^c�nID��eQ�P���(�l���ؚ*غ!�S���v>H$�x�)Q��:��`J��V9��#e�{/����s2P7�˧jU��e�ԪA�A�~6��@G�d�z�.��wH�+ڜG��|�CzH�+�-/�L,�ߜ�<��ɵ�e��m-�;��Wv��Zζ!��ș�2\��K*�oMwL@H�%�6�x���g;05�#�D�m��s�9Bq���`���r�'L���ʸ�͹W�Bb����Є"b%�mrv��x��e�TfE�
#���6��gl+~�y�G�>@*��$�zP��z����
j�_��٧�2�yI$�� j��r������P�L�\?��x/�:�]�."�bmW߼�{7� �|�);'lYԦ.��V�	o��bQ�Nk�#�%C��s��j��)V�
�y�-oS�+��+e���MS�2���.�VT��(k��@b��
$���6#�ÿT����E�E�����+�e�����<QF����n	�R�:Wi6�gM���H�GX0�[��>�����������nD(Aֻcs.s�|ǎ�PD���%�V	��g$���硯;������بe2���>�����hD��AV�U�dDuY&��3���N±𲰏��<9�4R�G�EL
S�0iw�8��eM�����u/�A?+{l¢8����(�6�ߖ�Jv�8�d����dsWgQ[�7Z��.Ր��8D�Q7�M�l,g��"%Ӿ����0��ξ>8K��hIV���\=�*�ٻpi�m%�s��,�%��ٝf ���Ř���㧎�9��蔳��K������!�gEihG}D޿e �r��H��,l��y���C�r_�����qS+pt�c#�G�D�_�)W�U�<[FtM���N���icu��O�w�j���t��367��~��u *��	̠���g#̭d9%�62�c���ȴ_��s�5��,#���KtJ���?�����ZTf}�tі���;䛓�.b��b>Y�s�L��z�%��^q}�(��/{a�)�sF�ָT�1���ٕ5��u�ZI����5`K�@���|�zEz&��A�I�É������vd7LP#�Ol�)��oP��z>�ި�O��4e�=ە��P��`X"��֬���e�|�s���)�/�~t�{�:05��%ג�r9�I0:�d��̍y�v����#NG��턜�,�3�	l��[��s�c�A}���	�9����QI��ı�8\/��k8�r�&�H���f�D�v^�on���O-ժ���k����UI�r��VJ�F�n���Ҹ�t+CY*JO�Di��d�o��`լ�d/9��I�0��o2��c���5��j�Icc����q�}9�F�(�Os�~��6tR��xpI�1�e<+�������)s�$?p�X���R���:�רIPZI��������N��������#`���}tGF���K�o6�������,%=\Ssj5�V�r�PQ!�;��qp���/x���1o VI]I�~.��ZQ�0E@�t�a��t�����<���v$���f�|��%�$�L���B���еf�kd�Ֆ޿A���@�^�.�i�������^��5(�c����2�[L�&^���#,e0V�5,ʗ*6��۩���9\`���<n7����NE�)��6}�`Fw�@'a\G!ݯ�����h�3���^�K������:i� ��c�	���9�P���*�FN��9R8��k���}��ٌ�"r�ʴ'��B��=�����G�o	�fד|N��΃��#lD3߱%��B6Ūʗ)[�}�+���l6��5*�6��E���-y�R6�ۘե)z)�~1�,�1�0���xO:(4�}�D�:+�����E��D��VmE�Ĉ�%�Y�R�����	Ca���;>����՘�Dj���}�=8�����X�ث1X?bS5��FBkz�7��v>�&N9����(�	�+�a���[�U�sg.�f�w-��4ՌݍmFǽ��ż�
F�~���Ȗk@�r����
=e�M�-�x�\2K�$4���j�2�g-`�Sb|�Y?��Z�Ļ���� �+�1�6�gX|]���u��	1*^�Xp��OP�S"x��V�V����C3��A��:�L��� �dh�M��I���9}&��҈	�&��z�3��FJ�]�B:����?e_u��Ň��e�7�N���@{TU.��	O*&����-����2�*H֧$���เn�ƅ �����X���=������C����j�8�]�����P�D{Esi^q>
����CP���Kg֔��&�|ci*�,�Xh%��t�"eT:�+K�:�
�#���f��=W��tw� 
�ŝ�Kt죯�$ӭ��:;hT5�k��ԛ��|�V��G]����������(�êN�ڡ]+."��z� G�O�5�Ɯ�N~v��0�q.���G�3�
oGϢ��>q��#(�:���B�.�0��M�,���|���q!@��9��%���zt$���/��u���]�u{Jo#�e�u�-����~�]���T�[sӥ�Rs��-��`�3���aV�r{=���Y��m�¦�_��jDXiZN�W&����y	"�/-� �l���"x�ܭ��7����3����z�y��#G����&��<�,� ���s�`.����BL� S�b�!��0 �kՍץ��h�.��a����Ɇ�S!S�hi�Tu�9��f��G!U4���>6	��X��Rz�\��l�Uܱ��j\�m��o����X��}�#�X���`c�ے�V�̺��!c���i]R�|������nϬQ�v07��+WS�Wb���RN�YY!�ȑ��aOVnP�!y��+�kMU��V����������O��<T�s`��:��C��d_(+�f�Ǝ$x��� �����ԢdWs�?"*'�a��#��)ߎ`��-�G�a���!�1Z{�%�,D���i���\&D5e�0�)N-�hXu�����xo�I89��Q2A����ˢ"Z|���jy�>$���������QWPx��1^]*���a�c��
���Y��׈��i�_�D�KY�0Q :`b������x���u8:��l��zE�2��+�>��9���x��>DB�4^^]�˯�@<��w��3���W�T��(��7wH<S�6�cc2�"���Ir�����v
B��:3lv��a�/AX��}�s���V_LÅBCq��,�Ȧx�� �U�4�Q	Q�׽C%��,)\5ޚ�a���������-\O�P�=K�D6K�R��#�~�^0׈n��f�d~��71�j%ul&Y�`�U<Fh���?>O�(?4��A�5b| ���9�v�oCqJ?�J����hN�\���컂:�%�ҹ�;�K������׳ࠄ(SƱ�O�n��	�TXz�K����~��S�}�n��.���2b�[3q��VfV����f�V�ͬ�����q �*\[X���P?[�8� ����Crn�1�~�)o�y���w�]��>�6����EV������U��K��,�/����{�6B���6b�ڋQi�����f��®3���2>R��Z8���2߾������`u$�����_\������F?X]�vL.w�V��i���;堽i"�-V�?8���1m�@��.�-d.'G#˜�;Ѩ�ߎ�e��69��Z�G�R���{�H�t��_��y�+3¡�C����7�C���������ǲ�T��ZE�+�g�*G��2P��l2���:dg��綐0x�Mi�m�<�&m����B�	�KKd3�12R��ub��"m�P���}���s�r-�E~u����'�j�1�Ш�cC-
վ�%o���'5W叚�D�x�eԴ����QQҴf'�=JƳD��<�=�MA�0^�݀�b�xk/���N��%�1R��{O�ĦM�
�/T?z%���Q���ڲ��Qʓ���6����J�{W��Vd u�L�_�����-{E9��+�.��a��68���Z��M��lW}\�� �G]}����-d}�2۷/�s�v\@�����^M�|����fuw����Q�ٱC�A�3�EM�?�g��E��K9^1r�D��Z�$5D1V`-�%�����>1"{Q��N���k�J�􄜿�M�{��-Kg� -�Hg?|e��G�ȟ�15� V�A$ò�	ω�)cY�'b1�F�˚��>-�l����Ek0�k�M�$��%�DR�,��'a/����Q�jz��b���e��hb'�5;Nf�b@x�FJ� _�ԋ-UC�l����5�c�8���㻣���e%�g��AH�;IVM-�Ѕ�>2�L)H?�a�Gҁc�;��M�iy1+Tc<H9�к\9�ԁc+Z|Fq2b����9#�'$0xt+��X3�
���$]?�5�6��ư�ZfUz����A�on�!ֲSLw澌����_:�<��u�(����1��aܞ�
����ށKl�n�!}�_�ߘQ⓹`.�����g�hn?��ш[��h��!��]<��t��A}��F���:/��2t;��T��^])���ׂ�}z^�>(}�&���}JwWx��^Uͯ���}�֝�f���+�ڬ/'�J��n6:��\��V`����]7X������3D����I��Z<�_N����������v�@%vhy(�����"�X�i��z��}f���}���5�c+p�e����0��Z���1;0�1+#chŶ�Gi�J��u(�a��4��cɰO��0��_�Nyj�.P�:��v z��H�A>����+й{���J���ۏ���e6��>���@�C�pG�ھG�S��;_a_�G*��M�0M��(�M�G��j�-�J���H�N�A$��S�����2q��V(��6���c�5��h����e
c��{��z��=���@�s���������jn�|.��;~�n�x�X&�/h��ٚ?T=3�P߁z �0j�#�g�>�2��0�il����|`wC����?�U��+۾0Ps�W� \$�tu�����G�{\Ǻ��z�����_����ڋ� �+��B�uT(	m&���8��[��A]~%a�=C�~h��J��Bw��أ~u�h6��H�K�MFs�sD��o��M�T��.�Lb*JW`��A��6�l��Wd̀{�QiD��J���Y��"�	�l�z��$����r�P�]>U�1O�c7��jTO��|ݓ�������Qq�Zi�Y�p���ϢA�\޼&�l7�~ ��+���ëi}\�Y�Q���4c�.�c�LD����2��/�6�0O�\D��d��N�kA�΋M��O�0R�a^LM�+嫉�	���u�jA�X[��g��sl��i�����@�J���/5#ϼ5yZh�`M�-n�s�8�\���[+�9�s{������j��o1��k�`7�?p�J�"��_BP����^{�����T�*�mQ�
�D<�0��jT#4�2Cj+���I]�&��$D�9\��'�%i:Bj�L�2ĈR�i@?�wg(��p�Xj��4ZJ�]����b�4}_�V�1�Y¦�<�hocn�>gm��{3P\O���ɻ��h���y�I�w��$~N�Y%��h� �C��t�޲��uS���6H�������7�H��9��/�Uo�������vJ��_I����p�R��S��������OBn��U���%�U��w�o�R � ����J!������O��K�3 9lt���n�����IM����{	H�{)3˶�.�u��É���h�J#�le����&A�!QT#!�}����jZ��qy���F��Du�`�2��d���'Xq�� ��㺠�TC��1ʎ���-V򰹝������鹆-E�x��BG:�pQ��X��H�}��]CvIh�,������m��K�87�WcB�t;���#��oΆ�����ex��`�UߣW[���s�b��8+�xO�W��}�&5�O3�3�j*ڤ�łv;g98>;y��H'�E�A�啚V���*�d]w_ى�j�������t_U\�KQ8���jS�R��6��W����@�C��1f�DD�'s��Dk��7��#�(��GfM��^0�f�������y�{]��
�;/\˶�����w=&���3#k�i��y��n"u�Gf��E��b3�8�T�J��'��On��>5_ �uq�Q�3MR@�=�w�����'*T�1���@ެ�9	o�}Q/�����/,L?��r��GK�Ѻ⪯#ޔ��Xx��T"0�gx���DǮ��!�i�*uw{Y��*��P���,^e6#H袹]���|6��l��M7�i�>N��jT�m�}6�`}%����ݕ��Y��ڬ�F�4o]��Ou�Ԝv�sK��E���6gЮ��.�qP��m���n��W�"bu���m�f��W�B	f�Yю+�eh�K��|��mr�WB���!D�b N�X;��!w*�aNy�f���02�1��8�?�c�۠���4m�ш��>�ǓxS�S�Q��Ԋ����Q���7��z.����*rP�>�Nf�~�m��GrZ�6�C�e�e@=k���{1�1�lZK��{[*�j/���s�˵*4i�_j-���6��и'�P�e�Tn��O��+hݙI��`Ԗ-$��٨ZA>��͟��6J��c ]��7������t�,[��P:q2QZ�xf�*�q#��=��N��`������ɚ�W���懗�og�RѴb�
鼃�ir'3�9�+����$��ީ�e�[��f���~�ϙ����:�Ƹ���E�ѿ��ʡ�ǘ�I���,�o^l&ԫoz4��"a���� ]����$��Թ�w[D1E�<���x�E�4S��ڪ3�;�A��a��Z%�ĝ(%:�	�4�E�eP���T�$ad���Ꮓ�F�V�uB=��*]O��q�i�����{�0�pR�U*s�|{h�O�!��Ad���D��mٛ/6�\��7ur��o���> 0�]^".հ�v��C��X�#6�ۆj�AB�9�l� �h�"HjqDc�+6&�u���G�
�vj��N[���$�)ۜ�1�v<��U�>�}��ES*GԥԀ}8F�s���0',�>V�����!Zt�(���:�ùɣG<�߼�4]4MC�G ��g�(�*��Tҕ���+Jl����,PĘ��}�UxaOʨGfx����a�f�&�/k��xt�fSj��pk���]30��9�O��eώW�ԙd���%�E;k��6���+̀_1�T������I��l8���IF:t��l���3S��j��ZeZ�E��7��R�`$b��R�n@��W��DA+�\���� ��a�/���+�
t��?]�	���a�jv��]J��El�]'�v[���ٹ��:ƭ����B�e��G�����qu�!���(�G�;�Y|C��@+<j���	�1�%> ���r����4���-P��o�
��W��\Ge��LA��|3eZ��@�\#E�S �H�́��!ď�&fQsId�M�D3��$oF^K"Zkv����]�C� ��w��e�o� �^����%;���b����W$ `m�)��ǩ9�mb��[���S��͗R�*�6�����͌���������(qogm׺Kj���㧪Y}ʵ��&AMԮ�3i�q*R<7)��}G~�v�.[L�=�>mQY���f��ݓ�L�z8�A"�.�ɂ���9�*Ѽ��8!��'�����[���9uQ�5�/%�����ÁD#b7�ȹ���se_U�I�jo7�g�c��Q�S+%ͣ_�ɍ/����|�7^��`7����B����V���Ǝ\��G��,�s]A@5�M�L��&b' ��_���Ywy����eO������u�?]�`��)j������zj��y��E
#���yG��<�pR�/�	������5��e�]�ˈ�B/蹎A��
�˨Ř���34�]PF�DS�1#LFq*���rM\��a�(�nCh�>�FK���,H�z>oE5Վ<)�qd����=ˆs��c��`X/�&'X-ʟ5�c��	a�������v5Gbe�P�vN�)X��(wJ���������j�х.�>�#2V%kT�j~�qK`��M��r��Z�֛p<sDtT��'bC�?KfJ~D=<V{Oy�ʀ���Ām}�x�/���1�y�G����f; p�Q�:NP�M![��{6�`�����k,l���#s�<�\#�[5��cCI$A1	�����'H������� ���%�U|�(�K�S"���x�������'��w�9�ߣH��F�*�Y�D1�w��������N��H�-�vEE���wo�ֳwCi��=k$k3�2�iS#��@;�y�2�>z �6:�y��M� t1��ゐ�a���<]	�����i���R��Ug}��w�L�s�mՐ~H���1ҊcT���h ��I)RA$�^���N�fAT~�8�?uuY�a�B/5�Vsۀc�k�ƴ�T4[w�Ia9	���wj)���<B
_-]U����JC�}x����亂M)N\A�=�,D�ɸ�o�"H�*��+�(�4vj#�8�u+Tq�~��'a7�)BK�k:��.C�;l���x���ERQ��OB���}6-�ZӰMS�W�� �$ߠ��$�0"��TU<��a��#Q��~���Vfm6Mq�)Ы!>�������M�랡ֳl��|V<0�D���sF_#�ykkM>L6��@�`FH%=_���I���t���Z�+�<��Rڵ�p�|����3J�'�5�j(Qq6����'�ߥ��p*��e�d�84��m��:; 2�;���'��_U�Cr�Ļ����aڸ��]��0p��:�)�k�K��th��ֽ�!�����snR >g6�J��k-�p`a=W~���ü�G_�B�K��tbKy^'���o�!HJ���Wp�����	%���`�ΊD��j ~ѿ���@�����6Qn���\���4Ң] �q֘��pz� JQݪ�a��agR����[�K*�i0��� �+�Qu�b�-�/>�;~Q����߶��Իi��)O]����5:>,vQ� `h�j�兘�?	��Z��s�̺K7��A��<��=��OA��M�����a!g�\��<�C���ZK׬����y 7��{}.�^�\��<���u9S��Z60D^��b8'�=�k ʑ�z~���~؋�S���w}�
��O�����'<���R�o@5�\���K�F(;�����{s��-k	j]O�N��Uh�-G�AI릆"�{��8�*^���k�![��4Ni2,�suv��%��_�oP�:�����|�&?m't_v���E��E�Sg�~,:Z�y䊶�+���[`{����rY�W�n���"/ɸ��b�4B�YO��6����|�Ck��A�1*�������rEUH*��X��Q���@3`�	$�?\�� ��O.ܓ��	�<����2��N�^E⡦<a��������MS3���V7�!��vG������#+i�5a,k ��p,� h4ʿp�`�\�A�/�����{`��%kB�F6h���mI��v���_�kr�12�z�n�t�(�}�.Qo�XC!��v���2�V��V���^}�]�]�t����.�5P/XgNN�7�$d������0���e&�77���d�u D��&O�X2z2� ��f1W$���%D@�&Mϐ��MJ��J��ڃ�Dp��oS��;�ͥI�t�?{d0�G# ���[��T@&f�����o�6� ��vG �Fe�r$����V��n־��h�X���ܜx@���8�������k��y�VG��VhɁX��2�*�	R�3q"�tX��^9���}i�N�ۣ�C�Von?��\h�o?e� ��pS���O�T���YWy���k����(/z�,^�:_jI�Q�U�Y�-Ю�,ڛ�٠{]�&F�|�#=q� �+��`$Gv�h���z�6���q�ӛ���)�iֹ�<s�����:�Ya�ߘ���`�Б�]�d�1�epc~�־�=�7q����8<�����Ckfd�*�:���v���w���ۻv�#���mN)��8�d�F�c�>�
$����לZ.�"��b���]�����=��|��W���?fZXDe��Y���˫�9p�%�����jA�`uf�槡0;"�c��g�1�����ΝsV�F�q�a�8��x���]��t���"��x2�m�Y_L�x L?Q�ɪ�6��� �[�N�ʕX�W�@�b5���������{��o;wG�a �4��Ψ�2��m7�R�{�>/"H_ـ�^��
��(U켞 �6ǃU0�˲RO<�v�����@��;��=ýC����Q�3:Ϫ/��s?[��j�]��L��X?��?��?��}sO�>l�T�5�n����. �ߗR�}������KK���Xv��;k��q�^��_��qǳ�1�m A�D��l�3�*t��IM�ꨆK�w�@V��~�j��J�Ww
����
�}<G�-Y�w�+D���}gV�9aE]�'=C�q�~"�_V4���ٟW�"�����C��'d�<��^� ���H��9VEg�_���3[=�F��`�Ȣ�8�y�G]��n�4O{~ט�WHҨ|g� 򥼗<ERW7��r��s|�s��DXS�<)QKU��Kg8�9��ع�6dįWLT�[���r�#a���W�;^�p�O����c?=GN�rX�zT~}�rXebO����bx=�W����ub��.F^Oљ-��CM|I�,y�O�o�˻z[�L�D�e��^�k��sN� �7���>!�K�#ݕ�.�]�%�`�6�_��Yƣ�vP)}=���f�8<қEh�3�r�Y��1�|;4�a;o	I�-��	�d����4�GV�����ⴅ�X*������k� ��!/�K�.!��CsW��bo�:I��Hyj!E\R�"�u���@�e�gd��b�b��ݮ��I�a��E?���	�ڿ��^�k�	6K&+&Mc���7̊�k��w�[P_��������Y�Qf�h��_�"]�(U����W�r�"�|�>�:7�L@�Ƥ�˿2��m�:ۈ
k��:-H�mI�W
�eu�Z+������/ :���s)�Σ��g�_j~$q$��/t��<a��8a�j�p.���O�{���ڟ�9-����
�9��	g�"�,Cs�-���c\cN����\Tzd���6���X�E���d�0�}���n���G�]�_o�֔�O�Uļ��^��\	]W��x�YJ��H����P��hDD�������0��gY6+�L���������[�����Ė�&ڄ�'S���?M�����3ӲU&��h��:���b��9�#k�����K>�X�P�kF=��������0�fN�E��'�{x�-o�8Xk m�IW��0����Wp0�qjj�Q�w�)�ز���r>���
���P�/(;B	)�1��Á0ި@�UY�f���|��{�,��"�aX��w9�I�ٵ~)������