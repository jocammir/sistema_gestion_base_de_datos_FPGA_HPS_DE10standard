��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��Nڭ�	�����B�#Z���?�4�j��0�ΐz�A�y�[��I4�fB���_Ɛ���-����B���M'~��k,���'zf���]A�� -̭���ҧ���D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T����	�i�q�f����}dV�KE���y���Z�^����U�Y�!�	�4��氳h��HϹ�S�-�À!����:x(+(��զ>��@�̋��,~�d��j@r6@�eЪ�b���>/|�J�C<�$�MFBz���"{'� ZsKy��� ;?��J���Oܧ+=g��2�
�>k�
��o�(�E��g'\�M*�Q��3	�ó�6&��^��vIt���|���j�M���7�8+��m
C~��G�h���_��bmzȩuAU+g���l_�f�D$օn����_�����OE81����u��\D'��%×��ȏ]g��G�9Cv�,[���`Gn��m6��z )������fx�/7<��1��o�0�?S�� �)|���yk9����Z:R�'p:$t �wz�S#�Ļ>���F����&�K�5�����F�=I9j��#�0,%ŵ���\�b(��J	G����-�A)[x�֚V� �XP�d&ܿ�*��4�
��������W�+�o���A�8������@/|J�+�)h��X��Y���w/BmvbI�ٚ:#Z���3�+'�f��\���f�A�༼������C�5�%B�CcA�|`e�׶��^d�<7�Y��E�ٍT�J��@,ި�?#��Ԣz!4��l3" �f���;1r�^|Q���u����M>�
���=��Ȥ�J�	9�Ѻ���c�����d$X���,2�HNE�P��@��ŧ��
�~�ć�ڷQt�H�Ӛր�>��[�Cd�Pq��W��B��s��B���l���]5.Я0q��2u8z]��w�"Q1�P��<�L"�#j>�rr�uq�J���0�?ƣ�%����h܀-c���"�G�5؆������Y�����q3>T�l2Z�t����m��=5�_>�����$�UF_���(��F��TL-�F��?�%����^fPt���;3�jg����ջ�l��7�~V|$ddJ�������xqwX������yvݢWr�&��\<�P{*I�G\��1���wWi�P�(�%���@�JB�T�"��4���ԥ�e�/�=f���ɏ�g�%�<�;ȑ�E#,�
��{g(L;c�,���n]�W��.���Г��4���� ����fK�Y�F�/8Eq��_G�~���w�s�8U��6'��h�A4�E4�����v���aw43p>f���7�������::F�7���>�4c����#H�W�F�W��&3oK�g�ό��LCHa�3YC�����"��N�W0K�8�zV����р��Z�z��k�U��0�Bk�ܰ�܋�%�=��`W���6! ���jV��+'�T-��Ƹȋ$Rs�z����ǫ�!�Е�+C�H���|����Y�D��O��Ğ}��-%5��㘚��b[K�ux��-��N�&���}&c@
��[ ��N
ƕ'(%F��o�`;�za#��%������9o[���;ۯcBe�(�<_��W�_"�3��4#}�. ��,"�g(�/�΁iM�b��W�5�2���!�~�]�w��=�z�}�h��8� �ו�J�+�+�s�( �`pZ�OA-�ӛB�|�I'��h����N_�os���u�E�������BH\���`�o�O������VϳV�c�(+��A��	9_�"zgy�xv��`����� �#�fx���en�vMZU֯rθ_��P ��m���=��N�SzP�$�!��n��ѡ��V�] X��H���'>�����N��J���|��/�z���Th֧4ej�Y��AHs�}�ʖW��4����BPA�JҴ��ų��"��4�J�`c���>�7xl�7��];����`{�|��(`@��8v 1�\!:�@қ{W�-h���y�0�D�P�o�R�ӄ�+i��h(�?ͪX����:,�g˘�BD[��b"c+< �EE�ʀCxI�-x�Wۥ� �ܙ��1��U'r��n�%߶�D��9��l�|��^���F���M�����1��1y �?��/,��LP�{���x}c�����ypf5wµ$�!|�l��JJ���ɮ��%���k�.�_����S���{z��x��)��M1��˒���mG���{���+z�:q�G�0U���|��b�1��^ʴm�����hN'"����@Re���l-���PQ?�N8��l�T�/�#�W�d�Ɏ���Pp2���į�4�f���	�)�<�&�$����:_k>�[XJl-���A��#���\NQ�F�����I�	�'<���-}�<X!Kگ?����x�-����a�v,��4�8���i�i��� ��'9ՋRu"����)S|i*R��A��JJ2�-1�\">Yv��4��̏� 9�R�7��@���p�)>���j�v�@9�$�����S�I�W���5����A�X�ԇ�p��0y��@@\��3��Oo���6�i(�+O-�AC�a=R�,%�ew��x��@���f���J%`���{�ܔ�3�L�=-�ڰF%s��T�RZ��S'�V'�d�)�D�)`m��j�A��Bh(��蓒���	�	��ښe���e���4����<y:)�c�����
������6����M�L�V�e3�d��t����<~��בN�ήm\QGp��2���TR=^��H)h����� ��o:�F>���(YX�j�ML�ט���/j�#Q�$��jP����t܉�)���l2�:���u����A��ꐟ��:M���e��WH�u��9;�~��������zٸ@�Pa���,F��䞚,�#��̡1�1ɘ��@�n�Q�D�D���S�*Tl��o9�=�1oaܖ7X�a(Q9��d��C�+ ��8� ���AF�߃������2J�@��+¶��d)b��gM X%%�����Ҙ�<.C\������+�,z(� >߃D�_�m�'i��{���f#�,U"ͨ�b����q����uN3b�:�|��7W;�]�4�M��=��G&�r��+��4��W�)W��Iʆj����9�^�q;fE�b�� [k!ʫJڱ%ߑ�� �z�lR��$_��լB�B�����5�c�*���KOy�ō�V��BJ¢^�Յ�t���?����BKI�%�p�����kY�u�*`����fղ����.���4N���r���*�˥a@2G3�_�)�c�G�xq�C���y�w��������6���\�~ۙ�g��R#Y9%�J/ՙ[�Q`Tq�(�nc2�R�ax�x���Eyʭ#�U��E������P�Nٚ*���0s�T�Vz��	��8�,�0�3ZD/]�7���mGu����[�7�!UVE��AL7��&;��d3��3�1a���Ah�6��71�	����
�q��2����=���M
�js��v�55�H��x{��8N�PKi�zy�5��i9���38v&�K"f^���]�~5�oJH��������k1pp�\,\X@���p���v=�����*r�<�<z��9 �Rlx�y�>R������6�O�}��7Mb9w�o��sh���:�E��"r#�֐%�+V%y���,Wl��{^JjQ�ٗ�O�;Lh��I-si�<Ӵ���hm��,��Q��f���|%kSl i�5M�TF_J������!�Y���mȷ��ȯm�����,6�{)M,�l�V�*N#Β���;�����*Em��A�,T9h�y�+Xu��0!�s\fQcmҊ,���׀O�?^��W2�P�΢T�_V�[v����*���8�i׀bxL[�7�`��-y*A)��t�O����܌�6w�g�H�#�qM��|B��q@U��70����F,�wBtB�u�mL���Q����$p�cW���E�O�T2����%px����M�^�;��� A�Z�
��5��Ib+��ro�v���`>pp�P�����Y��\��^�)�c���֌�u�/�����dĊ�RF��c�V�AѸ�瓴M,)'�G�M�q)���'����_��#�Ժu.v_�w�� �j:�Y3)2ul�v�\>�K�F#ᷟVH�����M0XG��~7�}Y+��~`�Oɉֱ3|Ҭ���b������-ym�����T2:y���TQ�R�V&�vfr�[b��pg�?٘����,�,�w�b��a���۳={l�1�E���*�b� 7<�Of��#wVƬ@��D���Hf/�� ��R���"�[�ȱ)�0��b�⡒��~��Nm�����͗] QS���ȭ���Ny/�߉���"�O�Z�|Ct)�q�O���ˡxG�A!ٿ/g�д��]�Ɂ`��Z���k,]��R��ݐ�l�y+x-�T�V��E\8�0�^d�z:g�
BT~���hy�Jy��J��+�f,_D	m٪(t7>��KZzBE�ח�m��A�.7�˝�Mo�x�_�.>�nO�����K��p�7�[��{"������R+^n*��L:c4�=8������!w�
�� 
G0�FRS7�F\���4d�W�N������q;��d#O�5M��ִ�n"���x<�w3�����h�[����pW�*/嫈�S�t6�'Ч٥`.2�s���ϕR��ma(�@٩MV{���J��ad�d��t)o��!O��{�t��Ql,����z6�����0Vn����� �C��D=��8;L7)S�ƕ���裛:J� o9R �(=�r-+��#X)�dE�"�����oOdm��|ũv$˴S�Xj˘�p	�b+84ʾB)є_��~�r�[�Y&A�O���^ ���X�Cx4�����l@�3�~�褫s{Xkf��0�)E;1��
�x(�j�x��o���}-�I�����@�~����N��ֳ�p��c�:^���Q=�#�I*�}TH�W�}��G-��Cs�Ky�b/+�+ƃ\ �o��2�)A_�W�ý�f�%F::�/vu�8q���2�<f}��v0
�Vw1�?� Z�9��L����p�;��%@�.��|<��;]p�2�M{�@]���GAח Ҷ�%2�~��q��[hX�NT+_�Yj�8G����.�f*��
Y�Q�����HK��7��XdҮBQru�}�pNZ�o���~�"�^�4h a���&�c��W�]�_�pT�"�܅S����ܱ|m�~����B8U��/KJwi	��A?�7l�����y�W��A��Y���	G��
_����B4 ��
X?z����5�?E��eĘ��s�%��>����!�|�BD@�����@���H���"ֻM��%)��_n�`j�`�<����l
}+V-��r%�譐Ոޭz$��h��f{.j:]Cݵ�(�ן�tp�Z�Cr���N ��}���4���B�v�F�@�Ƥ���*h�mE����� ͆<��ӱQ�&�0��n���jA�U��x+�4�WțpkF�����0o�h�烨�,6��lQ��l2�z�y�Nn�i��<�����j~=<7j	7���$z���H,+� ��H��� Y�n0��0�0���G Rx72��R�%�h=�y�j�C�	VQcϡi�8��R�@)0=|�$ֿ_[�ŒV�	jAey��zfD���5�QV�DY�y��י�O��v�C~Ԣ��7M�%��f�Zdi>�4v(��.��h[��~6��|�������<:�r0#?��`~k�N�-�^Q�o�C�#�$4=�u*�a_����� jۭ199a���=kh��&} ����耥$i`7��Ab8JK�.�o3a��8c�W:�/xa�p}��Z�κ�k���h���|ꛧ�x��,�\]=��/FUV�ds����dڵ��V���O&�=@�P]@;ʴ��X�4C���cw�l�e�4�.��G"x���&�@OlG�Ll[�E��@(۶�@�̟���|J v\	p�9�u5��[ PĦ`V��Y< ��w��T`~�p.*��"D��'���	wo1j�쯹���`k������[���wB��҇\BآAII?���"fж}Q[��_��ۘA��|��^A�p����+y�pҡ���j��bi
��x�����:�t0d��FA�A#Z�s<Ko���/��㝷5��&h]�Y�d	�<5�p�=���Nm�b��l| S��Gb�; ���Լ�S�����ڮVUo�����\��)�B�0��c�.����jk���Ǘ���K��Df�JbF�X^d�i�.���K� 1��^YF��2/�8�S�����!K+�c�4A��xԚ��K�y����R_-��@I�&.!Ng�_؟��u�>��/� �˃�!���c�B��NQ��V2��yZA�濾���8n�t��Ø��4J���ǞɂX9&�ȥ?�-���<Yl}��8�ha�]�
IaT.�B�\�j9mrRd?XVd8w��;?��3=��:�=�45>~0K_�Q��c��9EmGtw��nz��3խ�5���_�l FEr}���g&�����:���j���O�,�����p؎n8�x�r�\�c��5ֺ���=�@�q�v�W�0��
��Y�Ƿ2Qn�@��	4��]� �I�		&pڷ�ܔr�@A�x�zA��4�,�䔕�;%��b.J!t	W-)e(Gb���5R�,,�?S,�Ğ�+Y��@�ށ��(�2�A�/7B�T��`8R���$-EL���#W�+�5�>5�恩|��+H����fu񙭏�h,|d�)���%YW�y��yOъ:�yF7�3���+$���ۏ�-$3�&<�}�����Aa��3�Sf��{�_xzc��K�?�{�r�`|�������]�ةL:�eA��{��S�[�y��-:X�+�gXsgDb�#F"�F��#�����dd� �X��7Ӌ�¾n�O0���-��@�"Bs�]Ե\�]$�V��r�sU��CY�$��B.�ߑ�r޶:�F�v��&�y�\1��WP���g?g�s���-���	 ���-���b�Vߒz�i�]'; �Ć��p$���e_�0՟�8��,=�쩠	��d,�*OP�o�Pi��]A'o�eH�3մ��������/;z�T�'�Z+h8��8�#��� �u<�L�٭��Z��#�B��WAˇO���F*�ɴ3*��b��g�&��G�U�[-���2ٓ虉���\;�G�����==M�	ȇM����Wa|����/E��o�曙�k���%@1����Š��=3�27�u�?}I�[�i^[�~�|�)���^T�@�F��[̆ͧ����P5���]gY.í	h��.P@M���tF3)5���:�U�^=�+
�?<�[m�L�����_��8��G�G`�jv{p��� �0���J�����;>�OQ�v9E�4�w8�k_�i��Ty������~�[o��]�j|�л*M8Ȗ7�q��@��0j��Q�2�n�9Va�j�nz�W����R�E{�R`��q#����_Q�ר|o����*�\w$Π5<��hT�r09��~� �Fv��:A�I���_���l����1u)��?���z����e�x04���Si��k0$��LN���U�Fy���Z��)��}�%�ek��и�զkj�g�%�j�h1�,�HR��Q"�X�����(�lu��?��>����<͊n��b֝yW���<J5��X�Ka�EE2]���շ$r��l��������`1�k�EOF���ޛ�.�ih�p�������3z�3Ƒ�qw{)��<x%3��"P 5\�i���z/���
56r����$�o^�*
W$sa�n�w�����m"����E����-gkQ��H�ͬ�&^��f���AwƯ�-�w*/V�bo�J:��'[�����D�^%?�S�ڴފJKb��(rIA�`"AB	c�-��Z'vT<��F�|@�,�M6"����,=�� �y`O m�b��)��������pc��!�b��6o�6*ƺ���X8�@�T#U,�8ZsL��UŻڪ�L�ӿq���������h��>B��*"����8�0��NQ�<���s4^91�S�Zx���~^N��:О��:$�š���1R��Q��\���&���L"�|�0R��3O�� ��[��zݎ��Wr3p�']�n�g_�]�꣹w7���zsFN�v�om��>�����SK���^�Q�E�2�\��O
��N��$�UϪ��}(��;?5��}Wu�e�e}_�N��k֠5�kA1ٳh�,OA[���/|�J�\��Hf�V�-�۰MK�G���0���Jq�;3�������RWuVZ1�U�vH��:T���������>��5ի/?P�6�GW�\����mz&r�'c�W�z��]������WE�Qxq�&a��2�T��.q�E2*`*�,�i�Γm�	��R]z�#I6���}[�Z:n�3�����N6��zM
��!JWG1��z�����!o����or�z����hbk��w|��q*��C�S"5����]�$�*��X�N3xBphm��\�2z�"�B���Oԛ����b�����ҥ�>��g}������rAT:�E"�N�VB
_�\�/�� 4�I��5**	�@H[���[nާ�ϸ)��S���vWwR�*D�z�7��4�X�
wX�"w����.y}x�?�L����Ė3r�8<?�hҢRX�y����Zx^����F�tvyg6�^��Bh���~��)�~1���)��s�����d�t�|��n�������0��gU)��r^�|-��P���!H��Ri�sr��H6T�������ɠV}��ێV�XS���>�:��q�\:`o~�W�&�.�O<m�#��r��P�V�ѷ�[�p��7�h�$�͟���	g�������_�!E�T�Շ���E7 d����%vR�R6Zl���{F��|��ez�c9�{�C�bpO��Ĕ�I��푋�#3��)R���K���?7�+:��$�c��"۲����:��ý@���mD�V�Բے�l���2�0�g
���.깖��~��Q���T2v���<�$?6�}�b[��),hn��@�[Z{��Tk[�$��j�D/AzL�ǈD��/K�ux꺄�ҩ.*Y��C�zDC2�t1�J��N���?A��f_jұd`�e�,^כ���cbbHQ�бW&��x���hL�f3@?F��sp�3�B�j�R�-�wucK\p({�,�� =h��^u��׫Y�'�,�G/���ƚ���G_�� ��IDm\ʨ���>��l>�]���>��L�����cb���A���Ʋ�h�'�� �{�{�����B��E�|aa����k*8�����"��|M����C��|ؼ�-R{�1+-���@��zr}fl���j���A�1���u޾�*�8^�MÚ	G8��ѷ5232��'��_ֈ`�ɏ7�I�ʗ�I9�a�2'���_i��w�oU�D�ǟ��U�u�T��Wyc�߾��>M��z���o<�b�r���4*���t4��)a�[E�0�A�Ux�L���}C��c(y��]5�S����(�"�}�~L�,�:՟^b�?�m�#=�?�t�s3�� �V�O�����Z>�b�\����5��Y����>��9f�Ǣ�Y~��o���Sbjک�H7�%�ZRu䈯o��>����4M�r����67�?S8��D����~��t*�@�{����:�M<����rH��vZ�R����y�A�J�<g�+-U�%0e�~�9���LI3S��~f��#��hd�o���8�$�ց�'���)��+NW����R��7^��[�n��#���=����PI��:���sU/L�F��z4���[�NЗ��Ȓ���k��� ��9��u�gnh��9r;&b���7�2��f����M��$�YC����vv�=d�nRB#,`	K1�D6�#��#~�E�"�z�Ns"y�G�%"$�Me�ZX����Z�3�薑S��LȂN˴D�gtPL���U~��d�*��sW�C�)[���࿓�3�E�TxxA2�^#����`j�=����?۳l����$?<�z_߼�4�6x�� *DT��ơ>Η!�I��i&��I͵��J�rY)�W&^��y�]��ϗ�`���k�9~�\\���kN�PP����&}%Wwt4��	����4���D<b���BB��A��pit���0�̲�鱰��s�$��x�)�vz �u�`���N�Px˃�bP�q=�ZB<l��:���02�P*�!	��$�7�a2�`��v��lؘ-Ϗ���..���Y�-�jW��N�bp�ñ�vYo�4���!�����oh�<tA��OL��ai�M�TŦ�8�]OP�:�1�э%�>�m[���w��{#76[	(D�P���f c�M(�R�k ���d�t����>�:�������Ǽ�'��bl��+Fd@�I�2�R�|��� Yh���]�6��yt ?ˇ�ӌUd�N/�m�F�W��`�����/���V����8`u���Nf��k��&�[B�����済h��֮���I3��5�g���?�ځ��`��c��CBӁbF�l"���.2�Kf7�	��v�UhKW.o!�悓7(RmD�T��|T�%����Ȝ�ř�-_�i������n_:�yIŇ�+0�Oin%o<�g���ܻ@�wڲY���t?��h]�,Xm�if���Q'�+�"���n$���4�IC	$4���k�u?��m���q"g�xp� >�TF ���3aB�K�v�ၟc��R���� ����f_�n��=�`��M��Cr�ۘx.�iJ����LPL:���?�"��kOWv�����5��p��]�l�ﮭ����Qv��B�F&�4��)9_�ySB�+�\ϳ21 (<��̹Q�[:	^N_z�i��t"���t�V�g,«�f�$�;�@H�fL�0�����8rl���,Y�}�t��;q+5�O��}//Z3��)���fs5�(/�[ک�s�/s�"�����D��/z�]m�">���u�󱕂L8�팠��}T���l���󤔦,U=E-���6�m��rU?�q�@��0��ݸ�nT�\�#`7�2���i��Տ=��l��Y�2�9;@(�`�Ub��v��(�)v���0��	�z�ı��9����;��m�>�$�xX��(-}�,�F ��۷�=$ȋ�8��i;�Y��U�x d�:t+��(���t���U�]ǆ�j%�,�I�T�efEh���R�k8��AS�����ҥ�ޭ��Fov�l�u�II��s�I7��O[����ȕ�W����o�2����2�oB�����>	���*��uzn�]e�	�7����Bv�eڛ�m?�dɹ�9��S�bPB�!5����Ajof�ݏD��U��^Db��FrU�qұ0���)}��%�Fl����&ȃ�g��wҜVT_Lo?a�y�2���@������\�9I#*�S	�~�V5>�z�7��׽uw������Ϛ�����T�#u`����*IV���,�"[�(�0ygn,�l�F1��������*����/o�t��u�L�n��Hf��3q�z |iu4Q����/�Ձ����C��(�-P�Fg�
��,|ŲՇl�߯�tь���]��
��Ŭu��/P2�]8�.�3$N���e0^�n���Py_*�ԭ.1�o�dL�����a�<�99/W��*W�	�bP;;,�ߊ��n���c���}�$hqqk�y;e\�$����Q�E�]V/em��V��w0�u��sw�)6^(��9�4n��A'!����PP�w�%! ��U�"��īa�vnLI���B�Jn�*�4���U-��Q��W�C��}�N������F�F]dȮU$z���ˈp�"�Q�XD�uot'�3t'���K�&�o8�!��>PgZ� k�G^{6�.�J��3�ݸ����]:,X�E]��P�)��
$���
 1F�����5+�Ώ^���[t.����|��GC�"gI78��d�E�	�m����)z��8��%w�8�l'��^��eZ��L3�3tw�*���q��I�ջ4�1�Y8��|��w�����y�h�7Y��>����4?�M�V����3����/D��mm�؅�$�Et�ck=��<v�^L�5R�X�u��  K�%�]�L���@��ZV8+�{���1J���+�!�W �������1!�T��%�>�G��e�Uf�r��4�W�����H9�G�`,�ڵ��\�Jka}�����(9D4�VMt��ӅI�`�%�F�Z�س����Z�����x���횃�����*���Ӗ�!�-i#�ɋߣu���\ʴSɭ������A�0ȹ%h _�8�d��}j�°b���H��2����*KA�������65il�a	����rzPO�B0sA�!���\9fi���ͨ[e���/��xSő�iL�0J��e�L�3�Y"��~p����D��q�C0yS�+����8Z�?�R��Kl�]��X��t��N8s?�B��Yk�<��>(r!���:�.I�K��{���#x�N��׶�W~�$ߴ��ۉ��M�z�Q��������������93WĪ��w�/"nV��I����Q�`]q����p�H��|�}A�&�V���惩�>���?��bU����8���d�U��)4���{P9Al�a�R�Q"$�$��4��0+T���p%�+����n�^�^]��ǵd�-�n���h��I�쫾�'��������͂R�:�v��[����#��@��-�\��D�U�A�b�n�&|Ċ4��\B�.� K����r{T~��3��������B����N#ͩ�z09����tpY�5��pk�MgZ?9uC�v�3NvV���`����M�⁩�M��4�n0��O���^���U����0鬒D� ��G�[��AR!�]^|�	k��q��}�q������i�^B$�p�˺�k�KD9ߡ]^�'����ؐ��]e)(^���%d(N��SqV٦�-�d��%P�o���KC������δM�?�Q]��o2@f^4����$rZ�k�ޞm���YZq����<ɺ����p�GV�R�W�LW�S��'^�uy!K�8	(^U�ɧ�SiE$<���s�ใ�'{�*P&h�`���xo�=
� n@<b  �\5L^�*��!�3|D�n\Gɻ���g�3��<���:�.-����z�����M��३�����/�{���ݵ��u��!ޏ+����":��\8R݁^&SK�p8�6�@̎�M�d�/1(��}>L���a',�񟯻_�T��`�|��g��D)���o!F{#��S��~/�WcX�i��{��
�A��V�Q�����DdV�������<`�߶����-j2x��d�b��2�A`�cjf��s�Ӧ����~�=^hsu�OĐj}X﷘�C�����!��������'x9��j[lð&1W5D�<�V��IC}(� ��\]�K��)b���ʆ�-Nl��A Y�i?0����9��"��)Iշ�����n�j��1�hb�5����5a����px6~[\!)[5!�[<�3���z�R ���Y�Ǆ��p���U�]��]�Y���~��`KwIؼRR��=��娶&�!�O9����<#DV=��c��$��U1i�
�Ly�ah�|E��m�	�bl�O/�<�#9"c�,��	9!�w�P�P�kPrh/�H��̮vX�#קz+�b�J�yn��+v��q�`�#_�%�9�Eg�/���t*X 
M�B�R�2X!�㙀�܅La|U�
O��𱹡�0�c�7>��&_%����������P�OC�6�"�Z� F`�fZ[�fLYJ4p�-�x��f�-f��R	c�a�����F���fg�è��AbS_X���RFte O嫫c����6��wH~���e䔌ӢQ���n;�A��ǁ$���3@�k���/ M�-E�����,�fkhgN���\�s��A�R� ��!d\��9���6��h�a����|�	�v�%�oK��8O�:��`���H\�R��H_���!E^Jn9�tQ[�,H����<����d9�P��l��e���%9�3�oy��������#�?������A�������y�1myv��w!&>�l�]�B�}�8�� ���#�s���ߧJj�-<C$j��������C,9���"Ys/d7΅WNۑ�Ej���%��]`n�䭪��V�7m���8�ܗ����dCd(O.u[���<EF�]5n-����Z�
�/D�2%`�J1C[Bv�h����^�	J�XR��X~i�Ɂ��n<���{��fE�c�:+%���T��dM�N���I]��C��Nȇ��~���j�5Y��>�fJb��˗�J��^ƐZ���t���L�+�֠��m�}��7VDx����K�g\$ry�����53�Cd�oo����M�f;2��Iq����>��!"��D���]H ]���lvD֦��>�^;����`��䑸 Fu��nC��+�vg���C��XZ���6rz�g!�p��Ÿ�I%)" �h�"�8mR�z���_�y��#$�N��|/=Q�'~F���8�� �;ð��TQ���^�<\�b��a���#a�� .�C�8��odK��>�Me� W��������W��L)�W����f�b�����rY�%���qE��� k�[����4��[]�(���9fl�mY+�q�����#��y,�g_F����
��+m��f�˗6�a����J���91�+8� ��\�+B�����]�|:GNX�'i�^r�����9�����n��M�D�y�;�2M�鈷}>U#�X�ٟ`D�I�X3��j��s&<���M����J*
ka�ƽ��XbQ�lV�td/Ћ7�<��LR�[���O��&Qu�4f��kI�&&����O��R�cr�YÇ�d�Z�'�Ke�^b-;��(n�\�}�*�SuDFȵ4sP�'j9 �ǥ2=�-�QHC��e�?3����<-x�Q���F���`m	��>P0s��LIJ�a]�$�|��=&:R?�0cRя��i�_y��N]�y��cm�5~K�F�t_�VC���UI�I�'0H~-�� Ën��|�t��燒>��	�7r2�7�����M)x���e���u����Q�:���,
�nᡬO}�����y��)�3;�;�bv�����a��D�͕�0���
{����*΁� waj��Y�/!��+��Q�Џ��R	~�����8��=�G��S�܅��*M��~Yq�= ������A]M%d��4��ܽ�1P͖N�IZ}�m�Կ�{Z�\��d2�-��+˙���NBys�;��M�~��'��3�M�AmFF
�@��G���w���o���RJ+���nh!u����II�V�eub_�G�fe����y@ؐg��gv�#ѵ�*1״2�ߊB���W��?��07>����=s��as0ˑ�*6v(�?z�t�� �u�h�%fq� ���km �i�%D������9�A{�F��1�>.<�]�ٍ�g�Xŷ�����}dZ65$;�������)*�ն����ۥ~;F�Iv$3���.�} ]�H<�(oE���أ�)b�X�R�>R���l��l�i&�r�I���j�h�<��ڗ�Y�͜�s�rcx�K��q�|�|T�g~�!��O����o���:p1h5�H��Ye�fv���������(� ��m��%�Զ�٣�"в{q��{��˫L����!_��W
���,�f�z���,l�w�N���Py� +� Z�����{e8���@��S�g�E�2��κ���߼�\El����=�g����0�������׹�S�����L������S�3�fxL��Y�u���W��R��²ˍ�7�,s-]ӿ����-�I�A�8~)|f�%%/�U�>��*9���RVk�Qy��E$aB�c�O�'�B���Kk�k5a�����vH���� ��X�g|�h�Ê�jG�(�����Ѡǔ�OF`����d&��OQ�W̱���Vg��]9�����b^�ىj�X(�W��Gs�hFam�L���ZE:� ����S9�O����?qJ`qzIx9������JB̠����u}Th���z�R�+l1Pٵ �^�4����rzһK]����Q ;ű�6l�1�s1(�K��x����l�ʆh�W%
0��E�j�	�����1������{���!��<����� ��� T.�]'U�>)�iD`2�8�[��}4�s�h&ʏ��iJKFC�
J���������g�4Ubk�q\o�o�ᴩl���&�l CT�U�%o���9)�4^�=l
k��$o"1�~�xQV�4�ߍĨ��.ք�k�AR4M*{�lQ��OG������.��u�n�����H��^���)
 ��W�n�_v�Xf[���k�}>���d�/n���ԗz�W��?hb��=�x���8b��1�M^$r��ۼV��� @A.�WhLXJ��<ܕ���xc�!$�t�e"vB�;۴�j)6&T��z+�w/@�<A�ߗ(��SlL�6��[��[{�З^�cXgN
�I�I\�����({$ '��l�[���Weuc<������Z��R��]zz������:G�ߥ͗��c��\�����3]lpE���(#����%5�L	��qG`����C4z`����fx�%���{V���y~�����-�L�k;t}����5��U�'<�v���D���vߟ�L����~a��,"�qy\��+F4� ��:�ʝ���b���!�b�fD�Mh�!WXq��t��*Z<���3f��� q7�Q��ud���:�K��hh�=���uJ;1�b���Ǩ4%M����zӜ��N�Τ��h0;��:�C�^p��y�b	���;_�m��u��ĦxϖuSlh+��c ZgH�g.y�VO�L��J�B�j��� '�Tm��;P������10yEޖ�!O�&$µI�:qh��;����2) �aT�=Y�j�vic;~B!x*t;Ky5�~N�yAc��r����ӕ�Co�����C�f��5��jʨ=?�WW}�����e�|����^�8��_F���ų;�b|���Q���x���du�᩾�_�B�-l��AW٘By�@{������*%^��ܦݢ�Ya#8�s����0�ع�|MY%�|����԰�Q�X��M>�'?���v�ߜ�bj@��h���W�X�s2!Hc���1�P��V*�,�[z����=���^.��WR��<XjyIb:{t_�1�󷰕u-�Ʋ�KX�O�c14�6|��fLc*�c3_t�_i�ACں���_�R�]h�aI4��q�8�a�n$r��^w*�m��sO�Y=��ם<����o�@ÈȮX�Y#}�^vг���])?���PWp�6�S(MBHGgO�4�Ck!"�T
�J���W�� ȖG�+���UIr��F�6G��$�\�V����"��(}��+���
u���\�R	�ߏw��f/_�(2&��qc�F�mB|��,����1���Oqf;5I`l��7��g�A�T����3m]��!�`I���#1��t�)a��l�M�f�, �tG
oaW�懨��t"�w�eӲP#o����z�L�]���s�h,i��.S�rֿ�C#�X�)b�,P�����]�dgww"_wz��XY�;��!��Y�ׄ�|���{�Hw�DwZ*)�P֌���1"�� �ޅ�KKVL�)����:�a���ڃu;V����<F4��rg�%��W����p+���U�3���7�?�'a<�n6��=}~��K�␃��؋7K�'n=�Σɔ��ph�����Ye#i�DImq/�E8�RA)�_߭\��e�����]�rB6{���	�����"|��{]q���1K�sw+��oɨ�1�Q�
Л]�fqϿjD(1�L�+��z��R<��զ�K����`.hэ�s�����xq�Z�m������J��۳�h](goͱ��l �l�G0�yz�Hs��W-HW�Jy򎙄T=��Q�< 5L��;���l�h_V����O �<��Q˃v&e�e��'���7I:�|����)�V^�s�#*��Iw�"�7���׺��O膽�ق�o�Dqb����>,�����&���{��=�TM3b�ڸ�	+��8�5�a-�o�L��z|��9/V�$�Ž	@�^B4��Cpw-��-�O.�
��?{ �Ξh?#71����վ9�t�M����y���zS�����)f�n�������6�����-7���溷��Z�5�m��ec>،]�D^x��)A벤�����%4t��U@�X�����]�v)&�:@�S�r����=�8�K��0�BM�̺qP�hjO�g��ʬ�}ШXu��$���!3�~�v�lo��6��䶣�+��bs��1B�m.b�b�����vf6�.�X��%g���&���{&�����g�tJܹ�u�~�&$"�����a�f��BF���{��=�h�@,�@�i���g�3*8YO�0;���M�j�7 �� "#r����.��3��X���zU	q�Pj+�qk�ǒ6��x�fZ]q�
��HCGM��R�^#�X�q���'�l=IA�R;��2�*)���1&8>��ݑdR���j=�w[i���;2����ѫ��Α=A�S-W}O'�~SԠ����D���g5��*2YPxǲ͝����Y�Z��x�5�a�;T�Q��J�`�\e����׃=N��������X�7�u¡���o���#���Q�$
s�"�д�P��t~��Ñ�����}�?!6RR �-��l��N]����U���9��; �;;�N��%�4���z��4$k1�Vg2SOZ�3�76X�K*$X�����P"LʘK�t)2ԽcH�~0��2ݜ���ŜM���m�������k����'���_��s,�	{q�Q�Q�#�*���ղّ��|��%Q�J��X��\�"A s�`�
PܡhWv�c��Zǳ�il�����u0��T;h����yt�q�������7!aL$R3����uۄA�;[gc��L� 0բ �ĪC0!w�!=���4�����9���>>5�ϧ
�lʪ�	��7�����J�4�&[��?�QD�I���4���Z�+��NE�^�E&�0�.ޡ��v:,Ǒs+�Ӄ�[l�%�'�yA������_#���r�1=
�F���v��G&МP�Η��D����bz�m�O<Ԁ���:3�3�}�&b����ȁ�E�!]�͑���>Ӱi�rT�Xz/ߟ^�T)�"��g#�����;�"�yK��f�K�w�v�M�N!���p�,1K�VO� �Q��<Nӗ�2���	0���<	�L����j�NZ�`�P0IWA�2� �*�=��Ù��BVsS����49i�?.T����Z��'�&����$�R�ӛ�*q+e�$����Y;�:R�N�6�a���k8��2ytq3Oʂc1�hO�{��/��G:D��z�t��1*T���-O2�,%�]ﹴ��ddf��֙0S�`#3�c���=����]h���KO�y�{�S�� �U��P��(�F���/�j��dp��������M�Fh�lifZa>՗Y�Jm�7c��
��j�Q�1���$� �y>	�Fh�%P��D��޾�R�Ik�cR��h�����꒹�rj`���X �\
���@T�4t}�; ��u>��e�@�|���H��
]u���"��?1�I����L�%=��D�##Gs��b,-;&j��B�vFI_Y`��g	���n�>�5�n��$��*g��!�& ń�N�*�.���E����-�����u��� \m^�k�5�M�Sgl9ڏ�tG�S�1Ω?��I��.�������Gn���DC��Xx|��\�Ȫmi�D8�kJ��I�> ����a�^g��X;L˥7�^�,9R?�>zr�6�1�GEC1��}ŞO`*�V@}/��j�&u�&	�@af�Y�K緘���W�/Or�p\njd�hGFS�r6�q@�ʛ�,�YcAC�ۛ���#j�9E�+�SޗS44�=�ю�8t.;0�Z�r�3&i�(�h:]Z����`��զ٢ ���<��\k��;�q�A0i��"�Hۍ-#�p ��rJ$�A��Inn���|$�d�*ℼ���[��M�ge0x�NI�5��q���VYcr B�I�1G@Ë���||N&�o]e�����ڶEv��?a��m�8�Q+:��p�s�q��$ˈ�1�׮�	L
w�E���츍�b�����T�ꕞ�ax]���y�?��g���_a@�\�J�%^\�/��TI��؁Z��oo\R���Pkۊ�pˊ,.^J�m4�y�h��4S��`Ô�]�B�Y�~�0�K���f���K©�[>Hd-at�8a0�72�<�`d�ڭ8x|0m~�q�{t\��X3}�u|�~9 �A1$��]Ӻ�z��¸d/u~.���78�껛���F�e���`�Ƭ������Q��OG	sS{�l� �G���w�CIzU�-ҋBV�V݂�=�l<�cs5���j���^u�@�ڎ�`��P�R����E 4���l�mY
3������-��QxT�����ȡgw����'�C��Q�
aBI��%&�4�b�ھ��B�k�(��P�!�^욜����&]&N���q�/���e-w�'j�ފ;#V^hPy��/�ӂ�I}�p5r
�esC�|�y6nh������C�ϋڱ��i+�R��[���0; �j�$v*ˠ=X-{{�?�b��^�<,�^��� $1����P��K�O@�#��j�Jɳ�4_��(� N���2� ����xϾ&��K����YGW�{(��묝!@���bދ�X�/`ء��ji��@w�������.݂(��JW�_L�}�B��Ertl�oP_���)]5���js�wu�ϊ�P	d�3ۜ���t�����
��?M.߀[E}P�Mq ,�����<h ����/ak�)���hv��@�7�ɕ~"�������!�iu%~����$R��_V���^�N�)�Lt�r�^(:{̙[N�y��~��|S����BȦ5y1-yj�(F{��c(����*�P�k^�i/z�${��`�0s	���ÅQ�"�ߒ�Z�]����[� �����=��ug�ٝ=y
ҍ�A��q�ڲ�� ����A�l;�
�P
��nr���J�{�����~���o����t������^ت�t��)�0�s�C
�C�(���>�-��=j��mpts��cH�<<��Vb~�b=Z������$st��21ڸIN��]������r��r��r���ϱW|���d6���5
�~�W��,"O�-,��㽴�Ԑ����7�����0�k����y]�5n}�z.3��fv�-�rt�3q4[�j�j`"�@�S��t��0f#����'/M��az4�|Ç��H%��2� �'@�#> u�"�Bي�����(��R:t/P�h�}�♀���3]<��!���Z��2_8��~L��x���x♌��H�c��Yŏa�̕_��j�Q�pM��O�\��n�K�;��z�
B}��1�Ѧ�h���B_�����f��٥��x�ǰc�@��ngZ��J���CV�G}�xvl ���S
Q��Ҡu3�R�ȑ�<3����9Vk���Kє���D�k�-�$�1Y����zr�6�?J�{�FNT�F8�;%�|Ձ�"��84��K,���1~�Y[$�&7�N
=�gB�$j�pP�-b.^�+6U c��j��:�|L�!u�߄����寴e�V���6�{ض_��p_#:�D'ꕰa��\�ƗE���������ԨA��.��o��B������)e�,���3�>�� ������F���h��G��J0/�s��Z}n��nB��6�Bԝ��Oo�G��\B�u���ӓG�-�ݚ�g�B3�O� yo�ǂ+��@���ȭ�[e1j�B��X�V4V��f�n�A��`ζ/J�@�����WIWz�|��ø��@V<�*՛��߸;-)�����"iL(o'�M�����R
�F^P�GW12?Q��x2,�gEN35T{!n�:/xI�r,�
��m��j�7R�D�,�~�d��k�h�$5(��/�Tom1� +J�o�%L9�~��ܯ����#9�蟔Ġͦ	���o+ԙ��I��l}~��vB;6/���0���Q�S%6�D�O�D�`C��)W��Q���Djn<W��B ������!�K�-y'�P.������7*|Tx�x�Z��L��*�s
B0�l���oR��إ[��e�6}8����>(i��!�j��.� W�%� o$�Z��*��C�����+i�뽍�͕�yb�Y2��k�G4{,V���]�fT^���{���]g^$��Y8KT��B	3X�}�K4�}��]N�C0�g�T�	c|�R�{4�/V"oN#�Rp �r����C�UԚ!Ql�F��A�<�kQ;�Zr��[���U�Q2��ҥq�8ٴ)Ͳ\ι��9�o��"�>�A*+�4�K���͒��%�^��~_�	2B�C��5]=o�p�*�7�'W�_�-�`���3=��.�KҚ��u,�z�n�6� k����1�J���d#,�:5x��gx¥��PI�$�]�� K�+".i`C�%)d.-_�9,���~~2�Vн-o-F_p-��[�#�p�F~	��ِ�͎ZY���=v����mX������J^UrV��w:�jh��ݶ�%�\�>�b�BQ���Zς��0���p뮙�8s�|�@$C�dJe��*WX�+ۢ�ot�d�]�{S= �w���<��Mn�NhԼ��%�:�O����B���Y���-�Q��"�uB��q��w٦����9�_�����J�߲O��QcV����H���f���r��;T�&��-7��/zY�<��Dc39~��>]oL�h2�	�	ض�1�w'�e�� C䀠X[�fG3F�WF�EЄh�ܚ��i������e[d�������}�\�:�t,�c�YO	�%ne�s.sS�L��At�Ry��^�kݎ�6��Ӊ����L�|��u�߫�F.���G�Z��`�T}�uc������(���al�t}0 +��^����:psۛ/�1�� ��	z�a[��/6��������g�g	?Y�qL	1����t+V �c4��Y��Z 7~~�v��W霈���fO&CL�|�F�$�*lǛtɥ�(��4�;���k"�.��J�e4�o���0��w���:�e�2�-���O%V9hF9}
隀�Ckm1�#�F��·;N�<��+W<�V�ӊ���Aa�2�v�����ޝɦ]��F����"~B��Ӣf�~v��H�"���l\Ù,I�l�z�=(wt%#�i���(ȂB�Y�P�A_o��/3�4�<�cr���Œ��[(ktc���ۻ�n?���T�q��ܓZ灧�����zzd�I�ܲ�D+Yx��L�M������2��Ǥ�G����s#��&B,%�e��˻j���
���l,�e�� �/8v2-�� z�=U�K2���Ǜ�Zo���Q��S���{��E�������}�:4��~}��������L���01��IkĻ6�]D}��8���F�B�r�Eӧ_�� {��<v�����3m��'Ż�${Y���0ӿ=����7V)��CCk�elƤyi�|�5m�$��������v+�(FOIA��;p����K&G�UyڄK���:�H ,L9���N"Z̡T���^t�B��������v����)���:4�9���H�!j�h���Ajv�VJ:���z�P�����?�(2ʹ{������X�ů^R�0�k⹣X�{(��XQ����72����r֤�j�)�� ���!�����.��^Я���@�_0ף�����Y��!<o�RE�k��2��,�D�!���U��f�����M�+P�&�ۤYĥ����4�Q�X���l��C9!��S�GM� U�+�U��Z0�&���#4ۺg�#.>��w*����R�\�|�����i���,G��%�!� �.H���i-]�Ϝl�B�[<���m�"���wy������vu���m�I�w�*W��X.c��?��J�bz�u����R~�@~ �����z:�3��d���z�	���"�����;���J��r�i7 T/0�����׉��)��GA?D.���b�1L̟��L �#��'�u�2+�5�������LG
dk/y��(\�XⶶG�J7\�q�(�l&Ŧ��/y�AvŠ�S��1Ɓ�ۺ\Ϊe�����eb�'�]���(M�H�1��Z��Y�'��פ?�8���M��8%�Z���*�EB�:BC�@�? QXG�`.��Sc��{.A���.@��Tɥ����7�2( �~&����Q���y��/|�|���p��W�So�D���4��A�i�g����`� ����_�聉y�:��i6s��w���T|��&��vG�J��ثO���ӈ׵Ot����yآ�.ϬͿ��@s^b�5������A���??�z.��_l�
=�B�Y��t�mJkՔhD�g�fG�%�%d�A�����ހ��c��4�p��WrCwZluQ��v��q][�$L�KI�ow�j~�4lƐ1����k�Saj2�q��I���*�R�~[^�1��Q)��V��F&���ؼ.h0��<4z�I�wM��bV�h���~�t�j���-[�*�y�ۗmb^f�Ut���Q��Q��U%ڬ�]x��sH�Ο� ����俒��M�U/��(���z�Z,��y�f��,v��]��� mGͳ��:�MG��3N�ã�}��/�M����g���c|?��p���ᡆ�.�ܸn��r ���z���u�B�A���A4�}�LNBR�[Q,�+�l�n��S��+��I)FPr[K�
w����ƞg�����^b	]~���Z��Z�����ǘ�[�	w #�z�F
�g�$�b��V����W��]9��K0����N� a���6+�ͨuj��@rm���'�e�Q���kzA����S܌0��VB�~��+5m�,{/�q�3��S�%��ic̠GU��� ^P����WM��u�>��dd��hX/?��	'*�)�9������)�:������>�<����������z�<~C&�%G���Bވ� �g��D��%N��A5� n�)��e�HT5׊��12�2����ש�^.mv�-`L%��s��G+s ��.8T�f�<�����!-�aܡe~4p�s@Õd�yt�/#D���[pf��Ę����j�AxTL�G�Ԥ{K����A`�E���
��Z�j��;K7p��͍��O�Y��-I6�q9�0���+!�i}ҹ�����H������]#f�����S|��S�m-�4�%F��$;��8�p���	P�hX���\|}G�BL���D�Ѫ��t�W��6�C�N(����S�vy� ���k�*A���~)���V+g�����W2�w�B���53�Q�/��rm��ӳ勐�I1��s�O����kd9aH����]��^ X�$���V>Ӡ�Nb��o���QW��RCv�X,K��~�e4D��AbQ�	��1�2�a��I���4�=���ӂ^fa�@Y�Ǻd)/�JP�(��V'��Z������&���e���b�$�ǟ>�'@�������*���N�~n��.�mR)��Z�":���I��p�3�L��sq�a��Ӓ��hd�0�5
Cp�咚�I��#Z�T��d �X�F߃��W��G�+(ڹ�~���mڠ��"��y��R8`��d ������]�< �2R�� "�<��S5�S����!Hf��8�����<� D��;=�@rp-L�φ$H\u�Qa7�63�k��Cj��:�,Z�FD�`ɋ���PRЀ���x����u��.�=EE`9������#?滎�[�d�a���A\<~^	A��>�^^�ZO7�������R�5�o��p���-�V�G��s��S������b=�\�I��]��j���2�O��DT�p��~�@��~1>n����P�۷+tS��!e��%��4q�Dl����4)h�*h-��kKm�P��������L?_��9�Q�z/z^���0R�<��?��q���_k������}a^����H�4d]��rlۗ�\�j�@Y������W+��yP4���("��h��T����+w|OG��Ǒ`�OS'yA�4�>a����C9�7���v��by���N~B��^F�^����n/��� Qh����׸���y�9W�y�4������I�l:�������`���I�?�
�TD��
!��e��p�AG�\��ݪ򹟎��$�� '�
��a\>�'��h�c}�W�z�E�D����u.�b��aa,�~�+�v#$O�}NRu� ;�����.�  �����m�!�1e���)�f��A!&eQoO�vÅ�'�'��o���7�����Z�j�e8�۴��??;Z
k	�$�"0��"�P'�`�Vs<[�^0H��)�W��	c�1ާư��vꤙ�g(4�4H��Yaz���?���-
l�ꡥ4���l@��d��4{�ԍ���l�`��cK�h�+D �i���~�yAM'���qwfv$�Ӡ�&DT�kӝȭ�|�E�E7�����e�{��8���������mQ�Ş�<@��{�W@�q���}v�Զ��&�����-���k��i�B��ׄ�st�V��t��ʹaO9��J�)~QBF�N��E�~(j�9ϑmS������o��Ss��5.o�6|:���1�78�7��"��Q��Л����߼��l>ҘstEr#q�]��!~��U��D�"�=�%��,:JyI@2��S����(����b�Y�	<W��.�Ī }��iLN��VH�V�W�Iʲ(g�x���\u�l�`�6�ī���[���&���m��G�R���Ns�c�� h��E��<�};煨��L�T���>�_i��$V�f��lL4($��`#�ș��x�b/�9�q��A��N��e�fJU8B���I�8_Mc��̜�Z�ʍ�fj'�Y+��Q�+�\`���B����U��?��&�"e�l�pk��ʸvF��^m���s�tF�/4��Ѯ��j�)�Dn�6��~{�z���d�+�:)���^%'Ҥ�F-A�C
aӺ췧GJc,I8a���-�v4��HPKÿ���3J���cp���&.��kٰ��?�E�5�x�K�p�pq7�s�����u���[s��	Gɲ9q����ڈ�Ӄ�����u?P?��⻻MA��Ϫ�X�����4U��B����M�i�H������5U�B�|-�2`g�1��=>#B�ޙ)<ńCp��	k*�H � �Հ��씘��%|~����[mJ���w-����"V��v��U#9���������*J��S��R`��C�&���~����$o�я�qPvX15�b���AdD����6 ��J��Ŀ��K(�{��0�:�ue�H�S&@��S� �֥�È&�Nz4x��c-�*TO���?�����w�(� ������L֊�Y2O�Q#���|tJ�t/��q�P�Ny����ˡ�qj��ܪ�)_��S�j�	���a����D���6~��Գ���6��S���V
���Q}��� _�/W1����+���i�6�5�Ұ����y���k��3W��(ґ	�,B��� 
�i�3��+��g���g���S��Ws(�vl�@�/^�K���eW�G�"e����R�=����Qlp�;��VbKl 7��t%>�:Q2�I�3� ۴ p�z�]^Ke� %Ы�i��j /��lC�Q����_	q$�܁�ԯk����W<Xn�Aբ���b��n��0e���VNl��k>|�<�/R�xq�/�Zs�N4��z�i�����9�|):����u����A*�J*�"{�d�&��c�рQ�x��2]� �Ի
Kk�	��H�D�#�Ͷ`C&j78�������T9I��O5���gCS ����T�a�pt�X��_�w���ț,3�B3L_E4Y�"������'%G�,��1ı?���������TA?��($$�k$�K=.z��ډϡi�����)Z�O~ �9���/c����\�Y��;��7JK��%uY;=�Se�Oq�@18��]�`a��bc��?��eE���������;��(T�5�K7� OG;�ii�%�&�ʫ��[��H��xyu1��I�y�38iv���e��+9>�]݄&{�ղ��Z��?�l�g�L''�s�ْ���'M���}*��td]���ncG�w<ޑ�>H	���!4Y�?�;n�yM̢���B�h�s�#�(H��c��b^-���k�^@t:�us� 0j�AƢ,��h����T�,2��+�|���r��!���d�3������Α�����9 V��]�y���KY%����?�sJw��5���x?DP�	����t��{3���}��0а}���һ΅�8�.{��b��MV�e����D� {ږ8��=ɪE� ���6�^s��Zl���b��\;fF�4!��.
��p;�\0������7a��쐏��8�HWEt���F�������	#�&{.bv��_���F�p�4���󼪴��%���N�ѾB7p�߾ִ�"6.j~�7��Ƣ�{�'��8<:�Dc���z��H
T7X�&��ɯ�3���S��R^D����I:�4������b�#b�E!'���돝�\��LHv��SQ8��
��9}ʈ��Ya=9}ҽ�1��F�7q:.AMy^�3]Cf�]X���[�e�a��� �\1�o��t{w���z�,.c�H�Q�5�ƅ��
��E�0�p|�7������x>)�2�lPI�L�*����),�5�i�
���bϸX��
���Ғ;���Z�wrB��x
�%"S!�.!�VgqM�.c�	��B	�Np�A��r��;��K�iP���J��L̓��E���wݺ��|eV�'���_�F�mU���I�������_�+����=�x�U��.��8�}���v���R�l�j����^�D٬�Ko��c��9�a�`�B4v����R�"C0�n)��E�p�g��EM���~O�6he���lQG��Ky�@�r��ڲ���:��ј�ާ�S,8���S��T��/��J@A)���1��sgpvF�֞,/R<ۙۗ�
q!(�`�^V�jr��z'at��<��;�"���þd*���IC]�#xR͑0����k;�G�z\�ҟ�J�.L���YЬ���7���NT%%�~����l���lX�.�u�j"��+�1�r�`��[�TpF�&�)�Kt�6�6'�F�Y���1�F�բ�����^��r��	,@�ȿ�m�.5"�ˈ� L�_���(�独g=~^f�5����Mo4�yF���W���K����w~�Q�>��)�1�B��nH���j���5�x9��Pmă� \���f���Uʄ�.��\m�#�R��"�)���_��v�X2�o�젋��C��6&ў҅�@���Pg>�K{��{��?")���K2�o���M����s%r�)�(Ky�������.78I�%�&ީ���Q"y�]?�[���o�-�-aT�VK�>&��6bpъ��)�y����y���0��a�p�P;D�e�^`�dMY��B*<㉼V��_zkv2�M@�j��?$M'=�6d�^ �!�l�)��^�ݶ�읥�� U:c��k�y���mQ���?�u
�z�}�ۥ��s�ٮ�����ج1��K��l�_��ɲ�c�ed��d���o"Z\��c��/�ޮ���ʜzĄ�5N��_V�Dn���,4�� ����+���5a4�؀gf4~��J��7:e���t
�*�`$�ũx�t[y~/���5��п5�;ɰ��Li�{A��"�z��t\��@��F�氠J�=h)4����D򎖶���i��jl���3�Ǜ2WR�)��B�_���aH��f�J�Kn~�U��+I�-.�.��D��sir������y�<�WY�&�oI�J䋰������YBt�b�+�ǣ4�/���N�4S"�qTyc�o~����D��f �{�k�k���h��#Y3B����_e�F:f����sT�G�@���;���G;P'r�?�T�ł�p���"�#�O��2��gw��;���ItE��N�b���B^G��>�ˀ���z��=}=a3sAAiأ�Ҩu���&����]2n�����;I�X�I��?�����$~\�p4���'106��=��5�7���6\e�|���]გ{~]ʺ &�V�)��8_��u�
�I�qU2^f�M�Gאָ�m����t�nra�S�^'�G��e���}}�V����?5�bN�/AP]����m3,b�jW���|�ִJ����K!d�%>jT�?��رA�J٨MBΌ-<!��X�ã�H�8�����ɸL ~���hxk���7ru��ë��l��r�@J�NC�j������x3��
<��ɧ�t!o)͉�O�t�@<��0H�[�0��{�����>-%���-H�Ў��<���Xʵ�G��Dk-���/ڍ��rJ�+rw���)L,m[��3��<BVL� ��t@;ۉ�W������
f~�	��r?�sc��u���W�6̗nW�-��%�*y�y�p����))"��;���!'��άv��.ߤ�����D0�b4����ԞK�q��qw��[g/��ݷ[���hack>f!��+O�d�1��sUr�u|9i���V}�0��7ߚ^�a�� Y#"��Z�ɃO��z0.H�)��3t�R�G�Q���Ӹ֙����/��i/}ըEB�$g��;���VȢP�[�+�rn��	����D�0e�ݖ[$��L@����`�)���4�]�!�?�5�&��РjYd� �%��#?n�}�)%g v9������.$�x'ȰJ(�d�A��'��&������z���R� l2X�u�E�i�}C�`�U���� ���^S�6���`�`4�D�{[���B����v�mL���؅zW�%�	���pE�0�m��ۂ��7t^�:�t�J.�V*#}.���;]ܴ_?��6��X��Gcޟ�<c�՚h��}�1���`���=p��7V.��rW���H4���W	��*	�g��i@*�K�
] ����=��l�V�>[tc�_z(�z�Z�廁<E͆���^v[,�l�G#�vrIC:;�Kn*m�pƠ>���qv�%��2�rҳu(科��7�d��Bvr��B ����%�Ǝ}�c�V�X�<�	�,*�,�YDY�����q�:֊��	�QgH���[됊���+\$@���Ԣ�{��Y�R8����~�������@ "��7Ѓ�A�#�̂��zGAnn>ƶ�����Q�]�,wՅ��5D������*���m���n�8��ixϻpSw^R���P2�#�w�A���c��s��hă	E��1b�.I92d����(��n?j_�m^�2��g��J�7�3����է�	�i[(R���vb}��A�Ve]���Y��` M=��'Jz�[N�ɾMr�"���8��4���sE$ߑ����Z)J+�QÈH2&��Xd�D(���a�Q���l���� �J�Y���!�L��;�e*�t���j=�A�*U��,Shh7������+�Y�+P�z^߯�R,Oi�'�;�
�����v��Θ��	`r����D�P*��	Av;�s�cz�	!Y�^W�m���Ok��e����t�g�W���1�a��(0|�&4x&���`��h?T�]��b�	|i�4��,�ݷ5�}��Ea\&.��u����`Un�\��x ���\;ӎ0m��%f/&��̓��;Pj���׾�4���!}�Q�@7
M;�~�;0�=�n��#�v�}�UM��q��J�Y0�^b�B�w�=DƏ/���uݕ�S߰�`���O�L7i���1�;�P0�9t"�,���h3X0Ҭ��%%ʛϡjUS�����:"{ۯl�|4����-O�s�$�L��e�wb�����5E�eW��F�i&=4Wq_5J�����u�7��xV��o<�b��G�,٧I���b�j(�,r��;�����w��'ʠ>��sE?鲯<�Q���?���ݍ�8����2L�pE�E �C4TEP��m<:+�wuD28�Z:i��e<x�Kά��L��}(���m��5j��&�|�k���$�� ��h�%s�'͏J�����.q��gR�G9-T[w�>UU�x_.X��ǋƱ"D�ɛ�D�0�џ��ֿ�
��G%-9�Ӫ),�?�'�mlu�&��걛1Ll.�x�
n�D���Q)�7˵��g�L�Y�Rdr�sݛ��~/6��d�q��jd=��'���a�y8�/²�`4
oX��W�ܮ˩��׵�Ff}���� b�0�5##��M��Zۯ&�4�L:c�m$XMFYG�seV�twx������j�%��U�q_3��7�!��k$�y�������B��!��~�����t����աf���q"�ߛ#�p"u,v�1쎯=5��-V3v��~�ؓ�A4��_��>I�����:[�{"�D�We�b5=n���ϰ�]�=� Xi���	nM����������U˙=)R�%�[,z͊w�&�Y�&O2���R�ǂ�!��9G<��p~�d�i-R 1�  f��
.�٘U���ߓ�ĕ�M�4�����|���&�=������L]�fX�ߚ�Y�f(l��3�����(Θ�\�|�[���b:j��T}4�k��=��Z�n�B}N$h?��U̸��G�rr%�u��_o ml�E�.��/ZLC����ʍ����ɶ$��"�h�2��M���)��/�Њ9�`K�w+�]}k�"Y�������	K�s���@ο��p���:)�#�:2gj���>�GC%���~6�Y�懬"�IR롛}�����$�x8��Џ�=ކ�L��%U?%mh�U��ZZF.�.
�l�_���SǏ����D4s�X�	����e�	�Hɽ8�nz"�5l�Uo�$MF��K1�,��kb��SH�up��� ݌��;�f��ݟg�ۤ8�N�9�:L��񏊕������������$L��x$<�h�\��\�nI[�B��̌.�"ߕ9��Y|��ՎY�z[l��],i7�iBS�5;�:�c�>4�CaU�i�	��o�:'�n��If�_Y��8�ո}����C:e�β}��VR�݌:~�X�������E�vop���\�ռܫyx fm��F��Ԁ!�»G��<��֜�E��.�.�����X�G�Eb�ŀNq��<���+�P�pj��ya!�녟O.��6�5"*
Jg^��BàM�]�xO���1O]r�c`0>=��x�Z���O2����"���;�����a�)[���W�0AJ	�,H~�%�
���w'���>J�{��k��'�ΛE¿�h_㺗��kD��?�y�x���C��f��-Hp*n��kފ���#���׉d).�a�;��ϸt�:�5―�1�D>���2j���"�F�-:�(g*� �F9�b��.����H�����6�����Y)�9��qK`u�pqA�N�:v�1c��Ԏ�ŊH@�x�)�m�I�Q�H�k�!m�Mt�SP�y��`����tb�*��A8J���t�P˪Z���}>b���ڝ}�!=�*L��|�8J���t����}�L׊j�%e�(&��7����'+�8�f�K>o�I 0.w�L%�w��`߯ތ���$�b��Q� 3*]���^�X\�]qq�qml)XC#���@z��}�*�Xm3�����# K��ةz�|�%&�2 ĝ.�^٢�p�I�6�0�������A�W�S��-�>f7��AM�t���@ñ�����mHY�݉����#�&tT#��)�����}��J��h=�x����)2F��Gp��~$CDC �_��.��|儸s2ą9�%����/q0J��vq�dX}w/�M y�m�)���i�W�@�T#gϛ�21��*��D۔oA����VQ9m��R�kh�
��w^zd��1�Ļ�Q��O��f�51n��8�\��-��/���(�0X�T_=^݅���34&l�
�W4�q� ��~7��|���D/v�8Ђ0_Ƀ9��,.���Q�L`�����3=R���q�J���+a�����<м[��Y�A�C'�e&�ŲU㏗�	����v�+R���Z�a�e���B��v֫�#��tG9̞�P��5v,R�>��K���cAa�هrDLC�\���MJ������c��y8���>�5e��|�p�?�C5�^Z8�oг���N�
�΍a5�J�O+![�`��ð���1n�?��[���%�����bJ�O������+�=��jlAz^m��c����#~��w� �7�&s�b����+��ٷD�7��-"�*7�q�}�υ���Q�e5�g��J8��}J6���ZSO��\�x�����>	�ṔN!gzv
z�����a�y����"�ݳ�m��u�\��rCO5��;QY�M��IϚ&:k!�[Ջ����Ǒ��O��=���H.��X�M�D��I�w��kݲK�E�����ׁe=�ߕ�P"|��A�kJ��-p�����윚�?e�^O�0��dx�6��'��2��y�p�SU���57p��W�>��Z��<F�;rg�Q*O�߼l�D�Ѯ����k��#$G�Ŀ׽����탯n�ָ��K��Fx� ��d��K�;�	dV�&%U(�1�}a����~bѾ=���fQ�L��6(:�VC|����p.�,�,u�%�D�� #�1�1��=GE��S0�>�b�7T~����S>^z^У��,R�wl�!���}�U�E30�*&R��f)Jv&�?�!�*3�L�F�c��n5��T�G/�\�)¬����5z��6��{��)��p0�ra1��y��H�k���=����5 �$�Z�{*���=��ݸ��b�ًR����\��9ˎ�g"�5�-5����y�#YIZ%���v+�W����Ά/q�c��F�s�v�?w���e�TMf5{T�������
}�/����N�K�y 2kBJJ���YߦC���*�B����ۤ���%&�)M�,,������}<���|�QK���;o����]F]���)3Ъad���J�k��#���X���=�>�"�f6��4[�F��K�t �^��Ya�GBlm^�A�00�*J*x�>���|PA����W��]P[���ep�&��"=�߭�ބ��6����������gz9B�� ��*d�)q]��}$$>��|t�	�1$��8\�9����K���܋g`R����w��g+����B��w~Hg=1k�7WwsD},����cAK�E��UN�v]&}$�]'���S�E���'V�7��b��U8�;��8��5a��	�y���W(�^��aUGsV_\��y�v��^,�޻j�z��9��L�F��F������Dt�z���"Qý�#��J@�o��T�~�z��6�dpt�A4งû<È�?3����Ma���W�Ɩ��4��R9���<���t�ȸ���'�7�ƄNa�sM���������KD�R唵�6��P6���=���/��o�u����=�������"_��5z���\�Pp��f���D���T�]ͣ�.�`s�u	2�Q'��x�N��$�|h���z�Mܮ�x
��SI���6̤�c�͊I�^Ƥ�S�W��ֆm�*�xX5��{�m��+����i��[9�Rg����������^�vtn�$-�X���ֵd���E�s� �(��<�����O(^�M/� 쳣}�vO��%����>N]��2��n4<R@&�
��<k"��iA���8����5�n��dA�bzdE�F�JIװ2L���ǋ��+�N׭]�ۓʻ�ye6�@�.O3�MW\!� w�\��,a� �1qO=������6ezqb�zv���HL;Y~�[3�Yl�H��ކ����9~ȔL�U��#n�9�����-�`��w��]���>�'�r,���-�tG&�+���nG�b��47���[{5���������N�i�M-H�p��S��Ҙ h���p����"Z��Rt婗����Z)�aB�-l )�eT�	aMϺsyk��j���/t��_7h�X���>��e�S/綺2�LE��kꙟ���~�$�kxLy�'y 1����������E��`��,`�V���=���U  O6��P�2��=u����އX&���9�?~\��빦��`Ԑ�Cf@A����rvz��g��3o�{G-��\�~8�fd�Rm?�\���2R]��T�Thj���y���&F-���,y��[�E	� ؛de!��WIr۸���V�ʜ!POzj�1�(9j�h�b�oP��d�����c��7Ԩ`u�4MWH���g�}�ɼ�t�k=�"E�D��ҩ��Fx:$b���KQ���m�^�Ut���>��u��v ��,kXd����� m�h�Q��a��DA�$rQ,��l��L:d��*(�G��*5�>Mz Mã+	�n4�Es�DH�{����P��㰰�/}���kc��\N;1W����d�T�nL��閈�!�2TY�k�0)�|(�G��5�[����*�8@��׼8=k�/��J�(n����Nԏ 1ђQ���UOb!Cʄ6ۚ��k6{l��N:���M=��
-��qݸG�Z���k��m��B�Ɉ�;I����R�����0D�7�%���I;6X!��S�ǧ�QH�K�(�N-i�k��E�����3��Z�(�^>�I������b��u7��Z��f:b��'Lp�bVhoj�U#[&"�4;q�g��>戈k#
F����܈=�оx$�J$ܞ�Rjxy��{�B�#ͮ���P8��� ���k߄�ڄ��(��C϶v��٫�>d�2�s��h6�o�5E��j���1�r�/��ñ�	��� �d�������p&�8����F�&�Ǽc)���/]E�w#7�u��Gvkzf%����7}{!P�_P��F���Xv�~�ـ�Eu���&p�#���6-/ ��}�o�gJ��+kN�K�f�Ů�`�4&�p��A.�*���s�oR=M�&�#�}�& p�/�.�Ӓ�m`�Њ���C�R,����9����X)�I�z�S"��3C�SЅ�9?=l�PT����t/?��2ȃޱ�)��%6r'�o��)=W㫾R�|��ۈ+��5I��>�)����,J�V�$���v8��wE2
�Re766����$P�VDM��r�jN�RL�;\�T��O�K�G���-�p�_6͗wt��.�&Jj���O]=>.�<ѴD��E��K�K������C�*lҜow��H��(�� Fr�W�ɤ�^`�r�0z�7o��f��-k�W wM4ڕ�x��Hx��:��b��Z"��n�W��:�qg���>�bK� SL^�E3dk���J��U�Sw��eo�*h�8f���$6b�q��"!9O�'x�}O\H�����ؚ�[��JM�v�eR!�۪������m�٭���H�慛dG�傅n��]���i�e�瓎�B��a��v֎�2������;T�ʉ�Ͳ����ұ:��1�H~���#P��$�;My�]b{0���2��>��+�"���������(D%'V���ݾ�� %:�􅡜X�_p>��s�|N\�U��,���]M�bL����M�[I���s�P�zХt���b�A�Xt��~C�b?H�qKGM�|�H@������3Cy@�Y��[|����Z���G�w���[�*�]\����n9@UjbD��̥|�Z���D�\�mQ��g]v`H�+ @���34nۓy��P@��W�	Y�G�����YX�]h`k� �(�íIw+Q�.�z��C�fd�l�,Ft �w@)�N���Dà���=�:�#x8q� 
�f\�Q��I�t|�Ȃ
����K{tn���t�o�k��G��?�S��q�J���	�#p���5B�f	[ZIK\�+8�ґ{g�*��4q�|L׹y:?��z�8�+��^�f����!��w������nj�E�j5D���%����G��dP��f�"�W�|�� �Xq�ho����ϸ�K!شڏ���Uc0�%�����>	��D<��6�΍���&���mOY��ɽ��	���|�<�#���b8I�de|J�hl��;Eq���"�k�����P���Z2Vc�^G�Y�Y���3k�bA�>�$yH�hY�˯)�
BY�#K������1�������_���m'���=,��%��]�Ⱦ�!��픃��*z������?������ۧy.Ѧ��?ށ������/K�.g�h���j��2�>������Nɠ�R��d3�����!w�p��s ��z>�]�a�)��9���ܣ���Ч̗�v=Ѣi:9��Mi�~gJ���˃d��s�W�����l�|U�M&��؆�E��H�~�G��J37w��wm�z�!Ő��I#�.۞��b��񜕧K��II��@\HX�MT�|F�G4����ʠ �e&di"�c�QHOjy�H�#��jL�G��_9
����O��!`�u����>��0$�E^�jDM>5�d{ ��(к�Ԛ���� Q)#���i�u3o��Z���^�l�aOE2&��~���ACS⣑ĳ���a.{\���UR�V��2P��{���W���q*øo����^�bW��&C�Յ6���U�y-�ɸ����� ������j'�����#��{$)7REj�"��~���5IMe��kjݡC�@�٥J��c �!E�3ߏG'e��Y�����l�u�;PX�ڡ�ҟN�k ��� T�0�;��]��]%� ����:�h=#�X�n�/e6�r���bvL+�ֱ��wk�3�?��嬽����Δ�A�b��(��#h�H\�a����J�ס��0����渆A�<�7"��۬�r��)0C��P�41���@�@z��e_�t� O#Q;��-%�"-@��N��iB{����x���.�(�B����� ��ӳ�Д]҅��ʦ�sb:ռa�v�E�ݤNL���rC^�;����i��y�����B� �9��篺���A�.X,�G��,�Y&'f��q���?��EH��` ��\ON3G`U�D�*�'Sc"�f'8
�����39$��]Z���'���΍s��"b$�]I��s�^�f��-����AO��ޮ~��DT�i��h-4s���T��?<l�o�ZV�?,��N�)@5dIB�#r�>������P�]^m�/r���,��V�A���f���LR�,�Ӭ�.gJ�u�)�Hي��|Vv��!Mb�|�/����S1�'w%ˀ0B�=^Z����c#m�cD��{�w,!cZ)��e�7��N
S�1�啗k��~������9���"������n:)��J#��߯{��y<zbW�A��qV}��#���?�2_Z��5�V��M�xB.���J�z�^�8[Y�6���|α�� d�8oM�eW�+�TcӒ���!���j���#��50�c�_��'�8�����[p�,��E��<�-��M��!��&����(�t���x��a�;Є�_�e6�:@�XYܹ8,�9�L
�P����d�մ���])�J��>�V�8�A��T;�v�0-g�N�c��a��_�t��|H�N��uiB�o�7���a��U�~�.�a��=ރI���T Dс�t���X���e��txt�]S�[�!!s�1/BrEQ4��qRA,�*�����\�/?"1���D����w�/��A>&��f��~WuR�iCm��QL�W���Ր+��$U_����sO��ֵ��Z~p�޳[���]�f+nP��B`��b�E�Ї���3;�*Oo�^Ld�3��:��B�V�4g�b���<M���@�/�H��J�ƪ��v�ݠ��8D��W["�@�_�Ɨ���r�bP�n#���!��1c���ՊiI��\-�ֺ�|ٹ�p��=<U��Y3wrD4�!Q�D�oa-J����S.��PkOi�38R�$�-�O��>,��7�oi��W� ����RPc�-A���U�Zі��B#"�9���@�)hZ�;.�+��F� >���H��f�����b���<�����dx)|��~���I���[���������4������߅�Sm N��Z��wx��yO8����?���E� ��Ѱ�V�/æFT�т"T��g�����d`�_&,����Vy�_CĆC�����3���zP;-�"�[��61K�����������w6���FS�D����5�R<��b���N�V�=�N<I�#-w�Xѡ]�*�֍�5�-�*�1��}��蟠�2�#�o�o��d(M>sF�h�$\���ҷ�������էy����i�x��M���}�nj���eCX{���5�^}�k5�P	�ք����g�Z��K��DQ=�`�~1#�����;h��4q��������ԫ12iX�h�aE����=d�SbO� ~�z'�w���IF�xe4H{�B��RL����Q}�&.p�/:7�Y&�Gl���f��,�ePz�Mgܓt)O�y�yw3@h�Go=.�V�8�J�Z5��/�_�9�����km1a/(�;g����5y;�0�B}�^����<�jj=�0�܆���?p������E	:k�����x���D`<�<�."%��߹T�\��7��R �_����~%�TJtfk9�{D�����"5c�T��f͸���$��ь���__� ���*�u��}�$��>ڵ���U��<,�8��,��t8Q�C�YX~��	<��޺-�P0x|(6��Y��_�[���T��g��fm�>���\9A���j��/��¾��o�p��TS��S�I4���UG���&E��)	- Ҁ��T�0���.��F�9u*yqp���$ۊ_M�Fn_N�" <�6�<hr�B&��W��`�Rb4�;<�OtmQS�X������ʧc�$����޿l����y|�:�Y�/�-T�|�`Ӏ�/@E��C�qb���Yq%����W+p�LE���m9��p��=��6$59��#u8�RYXrP�gȠP2�HP^����=��u���B9J�QR���=���*�z��s�#�gm(�?a[�6���ⅺ|V�3V��h��#���U	�E�.ѬPs���n�Y8�1,MJ��5Je�D�G}���P�4�d�H���O_"�C��)F`)�#Z�Ho)}�Q����~��~P��6:��BY����Q�˒�\,V��=ѕ�g_�uz���;�g`�"d5���C����6��y�h���u:#"��$�?b���	�1�Pzv����YB)�;4��ˇ�*iK��*YȂ�YhJ���C��H{�E��i�i�z��ӄ'>���2IvȈ<9��.�z����׉�ǥ._���4Z઺���%F�v�Ѳ���i��M��k?I����PR���<�>��'/�����e1X�1��	�i�ʻ8F��IH���cC�zA]�꫙��n��'��?�@�(/72�p�w_^/�-u_O�$-�C�����oQ��h���1|��(�)�I��Hb�`Mg��S��_���L"���}-��1ء����'�����#�]G�c��w�Zҁ�>tچ��A�g-Ę��"F��~��f�V0b�q��2�Ej�{������j�L��쉶�6G��#��	r�����?MFC@q��ʋ���S������#��V���'��Ak�%��#&��n���������Y�e&�@�����+�~��&ժ���8�V4��{��e,�ȖPa��d0�&ڕ����_>��UX��m[E]I�'�Ё��N$�`ڇD����>	n>�� %w+��E�%+�3j#8{$�t0�������J��O���Z�֙��V���2#��j(t>� x��͙�<���xq;bfe�>�P���UŘa��LHNI�˛͏��1+���)^�[Do�������;�T���ht��\�R�L �C06Qjc� .�AF����%)p$p�h�@��C��:v#��-~k�O[�+Or��<�d8JmQ��q�s�"
_}�t�
����2�/���0��-�X��9�^	�A��Ԙ���J�+'�FJ�^er���`������/j�������(EE@;1�מg��SM&��Ҩ<�D;�A�<�y3��(yz
���-;Ykl/��π��	ꏭ���=RN�6���2
�^�L�����l�-�fI1l�n�>I����??a�Z�-7��c�	�@B^�7�	��G]����!��_��T�3v���T���Q�P��A1�C�J��/�V1�����u�mt9	u{N���h�I�3}��7���	�(?q��yeՉt�{�c�.�0�9�4�x�����X���?v[`.l�$&�w>Jb��k�rs�n9N+����P�� �e�����}�	���w[{�F���H�v����A>��"��@H(���n����qgb֚�j�97�a��d
e��/m�tH"K�U(%*q��[A.�V���
��V�[� \�p�زz�����@���P�H�Z��8�?�{+���f��Q%���tv��QdE�N��Ad��A7�	R�
�j�`����v&��&���z��8`�;T�]�T'�Z�b��@�\7���e��S���`�d�hp��z?	���hT�~�>/V,a�ii ���V`vK��\�lµ�b8��AӖE��j�<�;nH�A�����߳��Ɋ��:,Z���P^R��Xe���zю��'@�1i}~��bEO�O���[M>��"������3��rQ���@�׾�QVGc��x�>��H"���-7����.�_��J�L [�#�G5D|�` sNV1��P�7��d�ךqy8��,�Qv{'�������ծǄ���te���b"�˹�|;Q>Q�����26�ōq���*�ۍ��L\3. 	`C1m"���Wŋ�V�[��c��jP;���<;���;.���ݔ�H?h�	:�����0[�(FI�p�i�FpEJg@�7Kf�WbF�/�`��͹���
&�/bi��
�{tYJ�xdA���Q��2`Q@��S;c���X��!1�mdd$���z�f�in���px)fϞ�Q"w�}���Q]3���&�]��{�:82�ҖO�i@s�f1�:Ӈo�S��
�h�]�Ȟ�fh�<7�16����%��,C�~s7zU�Ub�o|X�.�.��c�>~2�&G��b��K�Dg@�5�<�ͽ�9����)v2$���8�d��R�r�k
� D$��(���d�='�	��q���n��[�|Fm����X�B,d�y&�M�s� 3��8�A�Z��P��8�QT�/D0�p���>x���1�<,�xTFObv-x/��l�Ͻ��>�
��/v�c�
��O�Xu�D[�8�hR��BT���fM߽�B��ANd%��J�m ����0v�U�Zs��D�u�W��hۆ�?crf��i��.�� \�۰��zA�P5�1�� dwއ�{����iq�Ё-\}�2�ӧUҼ�T��C��F����)�!�J��-W��-Q��������^K�鍸-1�ND�zX�c�y��Ѭ�ƯME�%WL_֌�*q������p�ȅ�[4�Q�ko���2��f�	z�h�jN���o�+����z�bH���`���������9�ډ���=��Ѯ�����Ϡ;+ڞ�����F��u��=:9���u��a�Y��(����7�~W���{���:��B�0؞�������'����5�{�q�S:���, �.J�ā�����&S<�-;�q����)���ባ��d����"��sw�9a4�xʛ6��lX���7�vf�ʛ�ș���H�M`��B���EK����e-|��
4IoJ�:�73 ��m��"��DX��Y�4��ɟQu��9�x�K&�KjJ
0k?	�1�2e&5����},?��nD�iC�T/��+)�!���{�=럄��Ø�4+g�Yc%5uлn��!_����!Zlw�D���%�Psh,H�h�Ȁg��A����M�ݽ����6�?)g���2[��.���&P�x�o�i�#���2�7-���r��uR���T�>#B=йMַh�%���ǸCm�+�Y�zC��rU�'@�4�B&$�"�\�e����(I�=t~k;Ìi8�J�� {؇_GrX\ч��7�Y�u�n��)Jk��u�}K�ҿKGJ"�E����Dn�$�iG2�LT�A�/��3��צ7����t�2������b ��4��}�4%q�%#��k9�Ŵ�ķ��O�S!Yh�b��Z�ܝ��h�j
�]X���wsNv�rY�N��4���T��%$����7���<��B�f^���
He��T�L+㞡�0|�� 	��H=�*���"�_◵
�������S4+��p��KM�$թ��Ik�h�	ɢو��@���es'qS��]i�j=ω�8�Ǘ����7�k�vN��@�{��8�Q�<�ml�Fd��5w�6��H�&�dH��flЪ�ԅ�~�2���V	;�;(s���띱�`P�&�7��O�tP��{�݄ ��o�g�d�8u2�p]�*�	�h�.�+��>d/������fK�o�z�6˴���(?Y�Ϭ�M^��x���H"|��XU�9��B��J��@i�J�h�}�I�7���^�GnV�9f�MmJ�ԅ�	$ه�~���>�
s�kk���v���-ܸPf?7u��1�ت�SӨr���=A�ܮ�b��e'��X����{s�Ip�fP��lUşy�T*���'�܍��`L�}7�n��
�y�Ľ})�"yi��$�Z���-�V`�h�m���6�O�2VԱ�,�q��B&Ǵ[�Cϫ��ܺ����_�\K�ݥj_�aY$�j���d.�\�h��p&�vý%V�j<"̓�3�̱�G��|mਁ)��&6�	.�щ��a��$�����r	�����&�3K��G��С�?�=� �Д�u��#>���#m�v���$II�(�1�5�~�(ݿz�Nn���!－�!Y�_=�����UD)��E���_�u�b�_�-�h��x�CdS���쏃�l��*���L�\w�pZS�~R��O���M�Q_i4��C�wU9������d�730���q�]�dh<�~�,�ڠ��t�Y�\�L���	��}O#��y�N�p�S ��}W�@5^�����UlltlA�܊����;L��r.����u��,x�A��,I����4��b�se���$>�����ɝ4[�*{����d_���K싶8ټH�	6t�@ϕ��#n��k↌פD�	1��z�A�Z}���^����!�70w�0�5
�P�/��o�������tJ�#����u ͡3�/Q��.���,����ٛ����Vw.{�k<����e^�Ϧ>%0"�;��d5.���-�4x��jy�w;gL��w�K����}��L
tC�F�8��Q|��"��HQTw�xY5-QNI�[&owTS�hj�~&�CEMR�([*���Y�FۄP}�WH�5�6����C���Ϋز+�%��W��:r�I�a�sW�4��Ͼ�q/aݾ0]Y����Z�2BV��KA��/����"�v	�5���&�5w��j	�-T�"̳?%{>��b*r�/?�a-0�#����
��������`'i3[�?h�箁x�bC�#���3TeNTp��[�Ҵ?�0yQ�{�(��T��Ɍ��r ۚ���A���Λ�[io�M}؁�*� )Gy�P�z���)�0|�}�M>I����C�a,6�[�l6i�xa����F������s�+�!#(;C�w��,�ȹ�$H_դ�&�Mj�l������c�jz1T���uCĒ>^3��kp�H+�*�a�N�x&}�e��v���<�{+Z@
&���(�NZ�P
]�}�e��!8k9Pb��)��T���O����x�ɵ@5CRI�Ij�B(*l���}h����5I��{�>�-e�7�&�j`�D�A�:ʧ&��؏�>�D[�9I~��m.wM�Q���R}.���3��O��獠����'�U����b����p�L�ƨ]�_�Ip�C�0_���x�6Զ�Թ}s��=����F7,�C��Ω]�N&��Bh���Q�-����ʻ���Q��
�/����J���倖�#����r�"ȶ�?: �'p������1�;����J(F����1="�lJz�U�$���q��N-"6,�Ճ,M3D�H/���8�_M��oKr}M��
�/��q�g��8m�� �x0�de�'h��,������)�%�s��%�r�/%��8xB�􂨥	2Q�m�Ob�r}F��}��<��}:3>mp�Z�P�^ý�IƖ���)�W��`�`w���\K��V��0\�P�{�yԏ�dc�ǣgH�+"��[�I�����g:7Xn;�����CO��Nka�y��o��]
�L>!�s�6�ʉ�S����'o��x!u� �%Y#ww%��I�rǾ��GC�YE�Y���s@g�*�B�/ɚ@�vIy!��)����x����*��p��_���	pR�I�:�N��P�6ʎIcǬ5Y���Y���[i��V
��0�:�?����-I��.sZH݇I+-^v�@n9���[$���?;Zl[#��8����Ȅ�;��������0�)�?��.�m���  G�(��XT,�|y�J��(��_�]�0\2t��"�� �پPTh"]���ҺA��������l��Ҋ���Q%�PP�hҩ1��z�2���ה*�ʑ��}�>�H(����g��YCX�H�G�>�1�$�����y/3|	<��.A��P1�Y	�H��č(�tޚ����to�l_!�[��`�ʋ�K{�;�6w��qR<�m$��b�"��.2�Ѯ��g���dh;%�i р�ۘyٟ�ɾO���ۻ;'F߬LP��%7�GjQ��72�X9�c̓ž	�8�<�-�<z��?B7ɶW���u�(�L��:��k���c�+�n*�N(�<���2*����&te��'���7�&Kl���g���Iv�����G7���`���>P��z����@�%�z�
����T��;��I��A�=�Og|j`zؚ;b�M��o�3�D�D��D���x]�W2�e�#|%;L}|(� �#�q��i��R�s�u3�ߍp�Rm9ǟ01k���V��]	�ݾQ��ބ���k2����0]+�w���^ �%�ue3I��ö�$�k��,˷�s��7C ũ���ff*��WFk�,a��#�A�J��� ӄ�
�m��i��*F9\X����^��
gl�o�7���۝�et qW+7(���=T�V/���[��x96����=���P�i����lm-�I���u)�i��\;=���T6(Ԛi���N��}R����6C2ބ��f�ے�B�؏�ui����W��F�[�N��J�r�,f��ݐq���.����k�9�{Ϙ<���f�R!���,!����o��ۓ?�g�柇�����^#�r�w��-��s&�&G�
{@��	X�^���Y��Yk7��D��C	V! Pq�Z�]�2�_a(�G��-;���r�DipdSYU�ɍ����J�ׁ��z���V�[c�t�zA�Վ)l9��-m�a ���ZJ6�߿��[���7�ϸa.SY���
^"�Jg�o�G�9=3�vw���='��V�,�M
�ίAT��֔��O`L�[sd�8�/�;٩�_��D���㉳�}P,��ٸ�\�?�p�Ɯ�`0�\��.�G�IJ��
�QW	�IfT̵��>n��5g�c,��넢�\�N(e**����<f#-��Pon��W� ����Zs#A���l�p�(�³Tȃ��
i7~{�zZ۲*'�8�r���8�9w�^�,�����س�6�%��/y��,V�_�8Du�1@�_�hR\��c(ۺ�ٌ��wN"U=\i0O�s��3��1ʕq��=k8�F:hv+}�G�D<���<ˎ���myp�V9'�|���;�l��A4{��jO:.(F/|H���=͜6Z�� �qbb��6�w1%[bP>����ߣxp��P6@S����zPDZÜ�^Ԣ)(k{���/7�#�·����ez�CŬRJ8E�!]"T
����?h&$�}�a@�-Cv
2�׿'Wz�cW&*˓WϺ�p	#?��>[s��%�)z5v/�����ָ��k�E��)r�B(O��q��hv&؊�U�'��׿�����n����+�r��'�0d>��.(_pW�]:�}�ӕ����R�*8W"��U�Syڻ��M7p%>��t�[��@�h���%�@dp�v�4��`x����
H�x��O4�o�6dey��T����{��sʩ]���"Lز뢉�p�܋���	] WY%�X�
&R'�S��^iL��eo�ա�n�P�������t�t+y���nȯc>5N�N:��5=)�R�H��v�a����V�-"H�ڦ��y�$��$���J�x��>PQ�L?�����H��"8v�_� �֎ԬR���+S�ma����ù �-*zQ��)�a�BR�G@tFR:|��~@�n���g������4�(�ol|S�{i�FP	&.�7d���X/Z`!S2	�7N��6�0ǔ�g���5����hQ�ϱ1�8��s�?$�X�����������Z�s�^ 
E��:<L_dt��I���/��
�鐠�Ơ�^,̪�XG��2|(OzS�7���Kƌ�Va�e�$wqF�$����6>��v?����,>��69��8��?�Ӭ�� o�e �����~O�g�˕�𞝳��rb5b�)��g����GM�r�z���=�#h��O���=�\����;��4��qQ;�5�E_W1T�:a����S�o ����1�κ��Ft����o£�ܫg�TO����#˝ݽe�����=�qaW�M/�j�1�+yO�%WG(db��8�m���!Ƭ�(*��<�8z����AÛ�s��D}������V���g��~���L
�gzu֭�1F��<����JW]b3Ae�6`�~�C*�DB��Y��d�?O��%UlO^ ^n�PI�;�I�[�d[- ��Ac`$�r��P%�#Z(J��X9�;��I�X8�����z�~]Yʁ�$t�w��o5T?O���q�n�"6pD�0��X�5L`�́$g!���kw���!��!����YE0��h�wl.��� ��\�x�ᶔ	���D�8@�����,��F�X��+�{�J�����.��"�C��_�X�ַ;��TzƐ� u���6J92�Z����̈́�7	��%���Q�g�DK�+DJѨ��y_������������"o�ɝ&���ϱ�hM}6M���C#��V%���?9K�*����]��I>��Q�n"R����aK����}�t�����]�ʲ1MC��O#�'7���]�B�읚�+��/r+1�k���[u��-��7}������pR�u���3.��{�擿�U�ػ-(�W��c	��q��/�ߧg���ЙwU�o~�
j���	��_n��dg@��b{�WzET����I��2a�Ա�_bq�qwN��FLabe���*ֿ� c�ޱEp�	����㘦�=r���yY K��� Ѥ�t}��,���H��@��4���3Y>���\����~�:-��n< _��x�n�n�jqpo��$Ͷ:R;����^e���dQ�0����?���97xK"To�P$;kNo��v������9�e��hV(�F�w3��)¾
���i7�V��U��5��1<i��3��-╫5�%��3�77잺�� !&2�h�����o;ԋ���,7�s s���Dv�x��(����Œ���ݮS%h�� T'n�u���F�[Ӗi�ɋ���c�ph�|�b�����e͔�4�vb����`{(ɋ������8�����0��q�.!�S��4V��\��7��:��l~N�w�����R� ~������4��B�w��Kvd��b�sD0YI�=Ҥ�E�c��,ؠ������0�Ģ��A&~$'2�a�q�ˆx�RX��=������>y�G�J^�g_��P��~�lx��jf�����zz)&V3���I[�g����s�����1�X�R�D`�YO�w�`#<9y�4 H�/_��|:��Q1K������3pJ��X|C!r?<G��Zsz0(�[*��(�_�k�[�(��l쬏/��� �r)����ڔ�_��w!�4¼�VDaeX[�w���yc�r��ks{b��3%rQl���=c��:�eN����+(���Q˼���������QK|c:���^�A�S��5�H0\}R��`ē�vm���j�4��`Y����7/���|t���+�[*8:a����d�:� �P-��g!�����W���#v̕�C8VD�#q�wGҩmȈ��H��6_c&��jǅy�s�\�䫽2:qe:'V�x��'�1�BW �X��)0�����J�'M�R�uRaK�-M�f����nB��-��.j�:x��$V� �r){�<Qw�z���t�~n�J���|Ҕ ���>�J���\X�������H*X��h�� �i��Gipg��3Ӈ����6l��Z�D��m�IS�Cst�g�xZ�,�-��l������<J����R����xn�/!)�����Cd�iC�<wR�@`#�
�gL�L5Au ��ș|7�����E�v����h(�?K�r��lP6A����JO��v�x���l7@@�	�*����H�k�1|L�s*D��_�\��A��ý�9I����^'z���|��NѦ��Z�T���$�4���=�YWF�.� ��e�t,��*$%:\4Ъ��G��9����5��0�ͽ.��>���A*�Ur�-!��6�� ���[��$˄�g�'V�iDMC{#������3�!X�4T��Dc0�eH�q%�Z���lg�bO#��x"� �.����Q�U��_mV�-!cI��ApQX�� ~���JVah��9�����;8�
�y�xY.7�t��d⒘^X\<�me��衚��4���i���z4/�;^!@��CP��M-_*��춟��ߪ����)�:�	ʥ�3�s�rvթC��s|,�9��aĭB��{X�zO>�Z����������X|i���l����@*ۉ�,F[��oA//>���g�(Լ|k�/�(�&R��|�SN�0뺋l�����WQΐ	��v��������#lH���&���@��7N���ׅpe�<�%bGݕ"<�����6��ۼ�DI�*��~��'l�z�5��"t��U}����O��vl쫑�*����;,�e[/&[Q^Ԗ/*���Fv���rtw�+�zH��P�G�S���
�k}��| 1�Q����{sk+(�w�ա���ڵ:
3"@՞�s��K�Z>PUw��q�>�d�2��"@����3��S��ΏD�^T\!|:�l }�z�z�BJ�Ԯ�P;�3S&(�2���,�#��|)aWY[D�a�z�u��zP�叮0#o���1�τp�&B4�6�2!lL�O��C�����B怇7����\�gg�u�/��%W��o{��} T^�bH�+j�Nmm�I�8[���6v��$��jƉ�oA�(�n�p�T$�=��(�#a:j��ko��Di�������E.n�:)& ��<���
U�oL���������/�{�P?X�!UT:yCi~���ҟ�o��cS\vL����Ar.�ν�ue��r�}v�8��>yD�	Zv���S�������%���cH@Wk����)����YdNOW���{���2n�C�'w���~����	�jN��-'@���9X��� fJ��z��� 
'ׯ0{��[mz+�Ϲ��]�&ܒ��q�K�BI����K̡-�K1x���*K��V	�TD�Լ�%�b`��$fL���VR���Q�/��[����1�b��X8����
�e9fV���kX����R��غÈ�Tj�>������I�Dg�t䣯��	�J�N��e(oד��4���ЛV�pD`!)ϕ��!JF
N�����r A��瞧��ɛ���!|9� �wV������>��,M�a;U�:E�5��nh��p�A��٧xә��K�K����
���4/�9��r`��LLFG����R$B|ڽ�iP��C��Y�;,���6sқ$A�Pq(�a���wJ����JՍ�>��&)y
��C�C���Y�zb�*DoC��"*>?��x�<���%�C�+�L��X:���Z��ar�i�m�\�K�Ը��C`)��9|�(�-�ʗb�J�I�髦x��L�#�s09ϻ;���N@�[X!�;��?� ����WY��uB�� �Z
��!n�B"%C����>�P���w۾<�hi���tU��j-�Z%#?��6���)`3�gb?�h>�� pU|�E.Q��˫�PЧ�����sseį������ ��BP	Pό�rc&JF޼���L6h�6c@�@0�*�o�B���2lb�#�P
%Y�\BC���nʯ,����u 1o���(/�G����C�N������WD���r���5?v���L�Zx�I��Eh�;��*�'x�!gX�{1���<zo�K�f8a�d�d9�&��ۜ�أ��FN��f�§g�]�5{/�v�FQ�:�� S$�J%����n@&�P/��I�D`�b��D�������Ow�o!w���W��m=C��6f�_DLM��f}��8�*X�m����ߢ� :�WO����$ �r�4�9Z�6zž]���ɒo�M���E�i)��P��ߤ���ZhAK�U�y��eHcqU���6PB
�Gs˭��@����	ע�$S�ހ��f�-7-�ɔ�}�1t$���%&_��`G��-�<���F�VR(��_�� �?��#Y>/����=���y.��a��� l�ʘ��%��'UK�E�"�/�$m�]���.Wai��H�ub_�un���O`�UX���9�]u���4�գrn*n��1��*q��z]��!s��YA���-�8B)����.��Kʢ�9�.
+o�r���h��5���*��q"f�:ylfJwP��h3����b��k�z���޷�H��$X�eeo�Ŕ��fw(��F��N�1R�i*H�ߪ&����T߸�\i�-(�m=K�UM���9(�ò�y䬢%��%���{
����z�H����LS7j��6���Ss�d��b�n��0I���wx��
��?�Nq�/��1&��17j�i"Y{�$4W�q�P��{νw�Uyj���Z�S`*����Dk�6����viN䒫J�#��8��A�'�mgߜA�)���Ct������W�+6����<P���6-z���S}���nڏ��T�=�0�)��S�ޑSgv��5�*�)�A���M�R�v
���K/T43Ĳ�|�<�<�����>�#֑�뿠�}��۳�Y�Ab�vd��>Y���ˮ�|pu��h�7葫0��]!(�עU<�%i��.S�+9�U�����w�m������"Z�}ٰ���Z=� �\���H�oN���"<�ˍ`ae���fi�����]^~�ݩ��y��"�T:sp�[pY��0!eӉ��6"� ���g��;���d�"qo�o�L����ߎH
�o�Rɂ$:tv��;�k�\=Z��z����!M�e-4�P�L\��6BeI-P�;нġ6B)� z�@ �?�+
�}��D���p��R��r�'�*��;��=;k��-������M!�:�E�y�݋F�� {@r��L��OJ�e(޻�mI��S��z����Ԟ(s˟cA(5Y2:),���.�vgz3-�4}^3L�Z��;]�H���k�p��9���r1����K��)����2�m'G�w��s%jm �[Y7����� 9h?�Xzl�t��ݮtaN0��f�(��:_�!�w!�����B,fw�b�;�X9$*XN+�"m�k������H�r��[>90r�3Ȭ�пx����i=����<����eҀ=U�*�s�%�<q��9XB��opF$��i�?��r�V#�=V���a.p��Z��c�>W�z����_WjZ�#r�>�]9?Y��m$X;��%i�ˤCN���s����m�;��ȡ���4I���IL�L=�*mmv�І�-�^�}�,��Z�:mZr3$�����pNH��ӈ4D\{u|�Qʌ�����A#Y9Е�D[O����/4���0�3�x>'��6�bj���`౺�!�p���<PhP�+)�����4�jI94}8GסʃI� ԭ-�*��v�b	D��^#�R�#�}b���c� ����j�<~����N*�J̶T��3���э�G�މ��6��Ec*�}#',O=���^g�G��"�0�=���۠*1��< <�1��@.-έ�S��bAR��'4�П�,�K�s����;%�U���ϋU"���J1����~uJޔ)��7q�u[����>��F&�԰V�WS6���Ƕj!����/^!r,�UQh�,|�w�e��02h3��q���"|kZ�$,ڷ�J�:��O��`��J��E��j����H(��~�Z�fg�HdB���� x�		�*�	eG���~�E���y�#��v�7���&�849,���?ak��O�����	���3�d�	\V'��⣖ƵVdL��1-�x`��۩� �ׇ��d��o�[�֥����.Ƙ3+������[���;4+���kM������󴒮@�_D\]�(͘e6�`�I5F8��FV� U_�+�l�Oܠ��N(p�h�xC�e����%)Ǹ�����D�h��>���'�e��w �bcO�v�y�G5:��)��,7�-e�D]3Ϳ8���-Djq�K�V�*}�LK����M��׫��ܣ�=�d`����P���Z��¶�5��di�n�+@�u!���
 ����%�k킴u�`��?���:~��=l�~a��4љI�ːh�[��p%7�	�OF��_l��gMG�)J�O�su&З��AfZ9^n�V�j�ٲ�����Kw�Jq�!_�	��A�B�{�6s��I�����E�x4�`	@�/[�{����,hn��|_��ݻ2�5M%f,�ED��v�>�% _�>�Cd��A7���d�a���K�p�H�^��yb������{�/�m:*��'�N�n������c7[��!�ï���'J��d�
��7@���ʙwc�<*���f3cv��#�n:�����n�8��z.�yE��g���y��~�%�j"�XG�FU{�1RX�$]��g���_�}5���7�*�.�p��ɤ�&�q��Yib݅�)}��.U�_,#�����5Q��d���Z���y9Tr懽{�T������Q���4%�훡��	�`(���Z��.�|��g��>Y֕q`��
X��#��'l�(�6�b��>4C��TqG�Z��Wk~�g]s�󽘶�����Z�do��m�Ͷd�m�&H��)y�j0�(���l �̞���w�n��]�W�=X�g�B��������������^�8��%��y�0E����`t�����鍐ҢpW�h:F�cR/�=aG�?��H�e.cu��9�p�����t�	�Z���p�&�]]+�mp;��&�)���w�y�9)m(6%��AB�W�V��7p�����#Л =p�9�;s�NE��#�?���&P�D$=�*r�զ�NH;���8m ;b���3���B���Kѻ��o]�!G��(���aQ��>����0�g�����!��&���c�J��0%�Cm.���C���;�嫪���P\ э� �A��֎���Œ�}h����\/���`A����tt��Mw5Λ�\]g����nKԩ{<�R�ٳlɆX�KR��J����iY�KC?���^�Ny����1h���bx�dL��v�pt���[8�
�;�4ҹ�B�	� �/֚�O�ȿj@�ϯ����",��=���J7��w�}�;�4�]�������>� 9�緍��&`e, 捷]<��c��\���^���qFe����xHb��,V���@!W�rz
�!o&v�A�pT����L'��ꔘɣt��ıJ'�^z'�]�-�����f�7�*����n��A}�	�˧��3�.��#n�q�U�/�Д�{\+���5�'���|Rѩ%>�n�-,[{���l9M���ܦ�<��6Iv)rAڙ�� �@*�}���$�9mC��]J*�36K�[}T�M(?0�Vq Υ�Zg��_��U���'�w�2�i4�m.�k+rx�d������mO�	�f�%��۔�dA/�2��� �09�v�ۢ�����&���w�o|��A,yr;ҿ�r�N����8tTn&.NdA���MS8<JH��΂B}]�J"�N��;���E��m1ס`����N�"�T��RO3B�wr�m����`U�ϼ%�6N[Bd��%��p-�j��~k��/��s��=�L�?�d�r�H`�/n`9�΁�QS9���%2(�Q�R�!��<�6�`��w?~|�蒆���0Y0�����k��"�"' ��}��h��:X1�D��)�VsvIt����"Χ��`��������񆇔הg���.��~r�'91���/G����>A��.Z�qө����^��{;�fb���&t����;��ҿ����1��s�Ϊ�Z�!���P�UKG�����:�F��|X��6 ��1�.���c�@{����l��W��.ŀ�=�HG��B�̩g��1#�#�k�19�P�fV!�ye�B��\S��7#���x����vG*�Y
��$�>����~���I�7���]{�!��_o9"�ÙR�޳�v�_���q�RD�K�j<3�t�u]�U��Vj�F��~��zݷ�r,�~ު��m��EB<��P��������8�L)�Ft�d�W�`�q~����@v����X�����:����U���3q��0�,�)-��9%��Ԍ��l�[6���	�^����%�ڶ�0��H
�#!�T��!w>��R
�Ć��D�R�<!�cjq�k���"���#l���#��'�g ���8F*/�u��6+D�D�Lf�Wk3C1'-;��0�k(��u%}-�'��
M�g�t -@�ń'$M�DE嫻)\9l����4~#��iY�PU�qOۺ��fK�#uS�)z[��m%2J�V��[[Ę+^7��Q����9�C�/�=������G�mDu��)Z��W:.#Ak�r�ݎPJ���� ��	����j��
�	�V��^	������Ae�-�{����``�V�v�&J[	�����<��e� ���G������r�'�������	8�6���pu�&B'��~$�C��PPƐB͒졥ï��y�<Z�#�zh)�<%1�%���<����+�'���v��O5��\>º��.C݁V#Q�S ^bg��.�#�)�C��r�v9�����D[���wK���%�Y~��
��>G@}*�9Y�'�z��z�k8���~� ��b�JJ7f�Ԛ��4�L_�e�?9m$�V���~0��2	��im
r]�?r:�7vR�7n`Q_{us�O�X��V�D`�2��}���?���^�a�p�8&m@�Z��Jt"Y�T�\�8;�Ф�Y����� Ո���]L�r�z�3��_�H����Ԉi\uuӎ�#~��%��\�O자ُh�Ӯx�v���1�?�`����6{�L0"��r�Xv%q����[���x�׵��&!+5M����
���=��kԎwX���s�3WJ(cJ]/��C�S�n���!N�͠�Ѭ_�s�I��?�4�{?u1|�	��`n�������������L�{`���h���6�X cғ�g�1s��-��D�QS��6酵(�0�B&�F&�?�aק2�p��,;����봚�Ω�%�٨�G�g��5)!�_/��Y3�	.�/�Tg&�A��,1x���{����}2Q������~�:�a:������t�QP���
!�)쯨.�?�7d� e7�f��Q��4�C�Jq� Ҿta�0�rC*/0��&R�m��1_��O��Ҩ�T�8/��߷pЫؾ�!�m|wM�}[t�:{Zz~��@^j�w�hM�,�ϯ�Z��Ð�=ߒ�}���V+^:i�g��4:)������׮�\s���0*<�4��\�����ք�
��V0����T�q����kLBR3G�!08<tM�z�8O�O�	��b	�q.���;K�gNx{2,"T�r��I���b�h��]��ly�l�$���vt]?q<{����R��-pdEg�@-,7���pX>��n�q��^U���⯧�@A��o�H�A��if�)��I�=�A9م�}��@d�kCV���e�@%dr����,s�(T7`l\)bskE��V�-�� ;���24E���K���j�x�Д�i�~U �W�؜�B�`An��g���p0[Q����=(�$l�H��ޛ���Z���?�d�x��{��{����0���
�x��Qwp蠮Y��AG�I�Mt�T��q�Vvk�+�)��`�J�O������(�8���R�@���f�i���A��IM��#��5�6���/F)��_��9yQU�7�ÿp'��X��oH�TLZ���dBz������ϝ�%��rGx�0Q�5���ze�G��m�ƚ*�Ą����Zr�[������	
�MӅG�_�C��*����v-9��]��>�h7�ǃ��|�|~ͻyߒ[ �ZףA����j���u��ís:�;��~��^wG��2�A���x��e��={m$nj�E����L�P���T�v����U��A���	��=�O����d,t@���>Q���>w#�o���0]��Ϙ�X��q�_�(��O*1ɝ�a�ɹS�kl#\��˪e�}{���<�G�+S��K�EG4<��p�|�����#�AkN	Udu�-��LN0� �h~ތET�5J ��q�@�ul�����VP)�Gpn�]:�m�n/��T�[r��zK�<Q��F��RN^�_�P�C�0dY��:�1f�����4�Ƞϙ��Ղ5���Atȅq�z8��N��0g/ۊ�R�s/��k_^�q�,�6|�J���/�~��9bf��Ѷ���X�=�#�Hv�� ���F��v<gh8^c|�K�!K��a�ܾ`�u��u�@�Ew�D��qMQ�;PA��v��l�:�w�[�
2ҷ�z�XPĒ��
.n�[>`=��Ƣ�S�g^� �+�Z�Zl�*���k�l�Ee@׮��+63?5d�t��@H��ZJ�ь�?����+�ӏ�(ꔤ�*�O a�:pH��HH�(O�k�� P��k�c��aS;����pQ����� ��W�M���:���@�}&<,;L��f���w�-�q�N
y�*�ux\vz�m�*�8)�Mɿ*٧4U��Ć������+d��Y�-C|��
,�lTd�l�u���H�����<�YE��9��Zp���g8�^l�9�X��,�ſ(f��31qJA]_&Qĭq�Z[��q<5���g�	���I��N���%� �a]v�]`�H�����c�Z[l
�/��K�I��=��zN����V�Z�!j�t�-&��u�_~�G.� ��؊�yGMX����i2w�]��B����m�*q�Sg&o~���ю���Cl�׹Esl
h�ю/��G�av�n�xL��{�Ғ4�`�:K�[��,ig�ZV �"B�)!�#�Ɲo�p��Xij�A;G�v$ҫo�m�$�$=vWJ��U��J�g�x|�EP�(6�S�N3)�+�Vm�v8�r�������brv��P��C>�ɘ0�s9�Dh�6B���y���{���Af����f��{0͢83�T�
O��!��Mܓ��+
<���޻o�D%��A�'��.�)T;Y	�>.��y�p���dP��
�������|�Q��6q�>�A�j�w��ҏ�XTX�򹕌� ����0װTk��h��F"4 ��������H����"���8�-96z���t�NCy|�"���2���m������.46mZ������m'��b�����3�(a�.8�T	gq��@=�ɻ:\��޻�)�4��^VLb���o��H�>t~�[w�04Sf�x/t��Nb�a�w���QȆ��ą�xdP��꟨���[���,���0^B1r��wrI��W#UF,���'�9��}}#�x�4���OS�5�8�X���tw�՟yh<ID����o��I�Q��=��5+S�L�p	�:����0QKOa:����ڴ�R��ָ[���չ'P���8�����I+C��(䶃6�#%"�\F��:|�:�--�uh���� h'Bv"*�,Qkq�Y���)�v4�V,������k�`'	=�]!���}E�a'Q���6��l�Dp��a���MG:b�&N&��?D4��*T����A���f�>{�-CHIE�	���ɐ_�B��j���So�όѐ�����_��;ь}5���m���W-��<��{X��b�(���Ϋ\�mA��J���b��f��u�=�'�WzU�ܠ�+���-lt��풜���F&�������ԋх_��}�\ih��WȄ��$$�i��F�z�F�.���k�o��(˝7�3��GVIW�$�%z�9�){�o_�׀Y�c�z+ys�~~����i���9y���Kr�U����O>�\U��ɖ�׾��Rn#���x��	Dk�5iKdo�JZ��٨�q��4���ei�֢޳���HQD�4��XM�2�a� ���{��\�ض�G�C��f5?�C�MMl���LU�R3��yz���ߨ8H#�D�����։���b���)$�(Z�/zI=��/����%?�%.��V�m���G��E"�W�:�(�!�go�����ϊ�[���w���ö�	�2��v۵���FR��^{�����5�XV}�C{�?�����7�t�4-���Z��J��rZjvL�IX�֬ڸѥ(E�|�cӪS�LH�*o����� �M~Z*���zǳ��.��#Fl�*ώ���9X.�e3C�Q9J���)�v_�$>.�3�����u�ݞ4��r0�89"&"9:�~�UDey?7�^=ך�-�ɔA���\�oi���N9caԕm��>Ց��w�]e�S�#� L.	}��i�Ѡ�F#�`0�G�Xq������T��m�PjB���o䄞�(���"����@B/����t���~؋�^k��=�5E��� Cr�����1#Y��ҙ�L�}g��j�����{:������K�?�O?	���b���0_߃����9Ŀ�CP��9�U/�\#R�;��$�m�O'�Rʷ�sf����}��i/�#��d����O���+��I�Ҿ	�P�{�#���0�OfT��5h������Q�.p��,0U��+��x �#�uh��.�qo��7Sa�J���L��-k��u���)2�G��l�K�\ɲ-to���Ks������~��L�lK��d��e܋}�#�n��L���*\@���j���Cs���H�)%�rCT� �+]ĕ����p�ay�*�`ap2֜`�/�f�٫�A�96UP_��d�U��M���~;Lux�c˴Aَ�H�ٶ�yy�%�I�xqϘjV�b龋�N4!趣9�	�[ܦ3���ja �"�����~"	|���5���b{�-���%q~]G�`�!b����-�Dm&eaBL�4��Yx�K���w�ߣ��2C5˙ ��a� 3��đ�n�s�<cE-|�� ���?��F���uQ�c�Q$��2'����-��
��&��pLv��_���4g��Q18�N�俀HPv�ݳ���(l,n�-0O��� H��	�#l�r <�8�������Q��ՠN�6�piG������h���4�1�#��Mdc��x�/֞���1�<k�FB�"`��!�-&П��D��vfR��G�j5^���"EM�KӞQ�����<J����s#ڵ`W=@�}Y�Vnə�@�?|�|���ה�<4մg�qSD%.֖y��;ٌBX��[K����1NC�H�O�0`A�F�I�R_����?/�.ǹ���qs�:J�-�0�Ǚ�����d)�+�_Y<�j���a`�M�Uө'_�Ҁy�]J��6kz��ޒ�J�,Ǝ��'�F`Y/G>�V��^��e\#��|#d�� F���sqWj�X	+s�^�OwM��48fێ^��#�6�<�t \��5�L����+ZǏ_>��'"���͑p�h���٤,�s���U�NzI�� ��ܶz)"�S�/�����lX\x�I�	vFíZ�Hw����\t�lIqJnG���9zG�
�$++�[B:[��?�ʵ����</=���_h#I�(C�����H�NrnID���H` ����Zj۫ܥ"�+3����qy����F��]J¢ 6�R�\�٪���a���� h�P)�O�Z><A��
x�Nt�KX1|�EY��Y a<w����vhN"�"�4���pR��Z:�x0X�$T`d�F-�%&�K����N��9���"e��2�VU�:/;	�X��W�H	��(���x8ⳤx[������EGr	1����O|����xq MXE��>#��I�x�8��'_���+�ړ��y�˷�!B�f#���_��>3/YB�feQ�g����{�*dƖ��dEe�9�0�r<��{�p#�,��F-o\y��5�*]��$n��x���L������Ҟ��, ,4��w��d}��7v��4MŶ|@@����~R��ia+���H`�$b�I?��w��n���xZ�T+�a�	h>���?.�PGaR� �����2�N�&r.ZWi�1�\�L��؛�R��AH�!u@�<
Q0�;�&^�E��z0i�h*�(��mxuO��u�_�=\�]��Ye7�#�R�s��g+��	
�T����
�<�=��'PK7QQ#=g�N!tΪQ���k�CRh��_ͺ�.�s�=NG��m�%��Lb�Q�B��O��+ʝ��N/qB��W1��l�D�к��Лn<����VO�?���H�t�[����o�k��y�;���V�,�a�����h����	^�xr���Q�)uDT9x������ё�� ɯh��0�(��<�z�}Q��q��`ӟ�M����A�r��}���>.B�k��>����F�+�5N\���}<�"܂���C	i��S`�,���,x��׮�Q�g�Y�ї�X◡(��N`g��h�]g�m+Ć龡�]|ѐg�U�#�����nb����U�l�w�H����F�_��lpKQ�oEw,~vF7C���xFƀ�e� �;e����W����0b瘌�Zu���y vm��;mb4y�`/�I�F����?�Ƌ��s-k$/���VP���G��$�������g�0�������ϋ����u�7C����M)��
��@�|��bq?5��>�l�� �Y��]_�DZ��Sx��?NV�;#�T%��<�����2"˳�bA����6'y�ok���$\�C�{y��"���y/[+a
G��yj\e�%�OkK)�E!{FG��7
�����K�Ӷ�y��B�W�<P�ֿ����*�|;X����N�4�$��T�"b�ܮ���P���ڢ���py�zGC�O�L��&M���=R�vs0�nZ�U\��8��Ň�\�b�m	@��ۥ��{d�G�8u�쀄�����	�Kog�21ʲ��a�kӤ�p����Q����)�3��	70���dX����%��_Z�W�I������2�ޢ>x<N���K������{�)'C2���wg�`d9&�j�#�>_i�	�w���B��ʯq�#��d0)cӭt�x{ԯ��^�j������ƿ0�BL4a���sU��XU�T݈#0E�l"<��?�)&#�����Q�z	�`E3��Q��7r� ��pL!�O�\)~+��v9�w�A� J�9�	�=vS`{)֮ ��n��?1K��G��iYe;Xwq2L�nv�Ӥ0�n�CONeF���ގ6z��{h����� ���S2`-xS�j[��2��N��{M����ç��P��-}gjK�6i���_>�7�j��^r�;"��ڏ���nv;��E��j��F�}�m����I�N�_��<�m��9�����e^���4,T9}rP(2��)ڰ�>TAG�W�_�X䈆]u
X�׽K�>�)=wϖ�4�r{�в*������~�פڲ�D嶀���nڷZ�D��	<��� ��{���˙V���S�c�����{�����O�m)�ANK�?VUhI2��9��b�;�ݨ��k!Y��ZMEɡ.��i�t0qmDX��:�@M/zw��޹9��kw� 	ҏ�5�(��]���)�U���r�Y\G�N<�^zû�3HUS����h�'��2/*�q���Ġs���CZ��%4dܟ��ܰs@$/ñ*�"�B�G�A���{��u��;>ρR6�<I]̤�{��P^6�5�d���ړ��QQ���c�������Z �O��A�e)���^��ir�|+��K��뢼� �m��fm��a���y��'�gh���w��P�\]M y�͋��=FA�OI��\-���_���w�:E����U�1��F enш�,��/�;���5�M������^�t�TZ'~�{����HbGF��!ɱ�����6�W��?��MT�}D���2HB��o"�_*�7�g�9j#=�`b|_��L���#3
�bɂh�����
��}^i_�ڀD���f�u�z2 �V�<Q��;�v#��pJ8C�I���!��׼��-�����z
^<>Pr�wV�}���~�.
��G�y�әC���RP3/�^1�gC& �`΋�����3��|ג���錆+Ȇ͙U?/5~DJ�t��c��"���*j�34`uΡZ��p:�g��"�ۥ@J�� �:{��?�7�*r���r�<aTЁ�^���v����k�ѷ�����kNa�5�S/L����[���A?gAz'���wց<��*� ~�тY��W�h`"�~֘��gX��GQ�Ѕ�{;���Ͼ�JU���s_��)}���i�/[��!�S+����D4�e^��<g�K��u���N�*�k^�Tx���|)��rt.�F���9x��1�;�=c\aK����%'����C�TY��mCm*aϕ�;�_�Ro�ց�vH��tM��������Z��(�4���t�Sk��{�L�t�'�o�F7q�R�v!p�O �"[�i���m筂=A���I�J�sM/�o� ;�f/Y��>7�Y��!q��I���o'��]yX#ɡ�~�S,(�[�@Yuw4-������K�	dJ���@0,T_�O���:��^�/7S-�BO�j�{�4��y�*�)6]���ټ���B���o�1q��gh*CJEU�����Yn﷑d�A2 g�J���~����V/!>p����~�?i����_�Q��F�mI~��UԖ&����et�2���`�Uک7}�8)�:$O��B���B�뜔z���G�@��8 �d���H2�f�+Q���V�bJ�?/ҧ�j��\�����W|g�a'D��gq���Z8�̹�#�I�4>���y&|+����$@����=SS,��HHl3 ���:h��zƲ�RM��.���Tm�oB���6e	*�ڬ�A���o��<�wD�X�Y�{}��TY�*L=�1���� �ɋ�M,зo��i՘���C��j[r�KQ��Sm.�?�_zo;ԟxȨ���Li�V�g�F�J�ϕ7y�5h���r��Dt�"���s\/�e_�A�ko���k\I��S�y��-��ч�B9�s�>p_e���/x����W�[��5���(F�����ou�ɚi��\������N*����T%��o�CԨ��&؃�)�2��,�7ne�d�~�fyT<3j�ve�y9ӕ7Z��HVG#���Ȥ(�}�̽�*����ۜ|�@5{�rp��{�O�6�N�h�C��FW+�ư��K�
;jWCa���/zc��ȳs�ƈ����LE��d��ѽ�A���%
wa�.hzB��2}ʟ"*���A�=�MWV�mi���@��]?� ��u�
��~�4߯X˞C�}�}^硪����e�3�٪Z�%�����_�	t�i0��`y�q�#R�J��dL�e�M��9.]swlEur�-��RLUV�&w,n����sIf<(P��m|�v*jK�*�4|�[�6�>y1,CZ�3;����\�����x���&G=(�R�̥g*�xU���giͺA�A?�ݕu�*c�VhF���>ɿ{$f�����9��!���#��m���h�~�ď�LɬG!�˽��z\f�)Z	�"tg3�C;h�Oc�	݅�}4�n?i�y����y�V� �0:XɌHB�jR��o�w����Dkr�w��W����[�zA�����NK�[�ŭ��	^t�aF�ڥ�4J2������و�N(h�:�e�������Ďq����v>~��)�F{�,g
�J���3�^U���ѠV-�E���/J縍�B�_�/�P�C H�$e��L�L��+�W`nh��K�A�!I��g�����0;�li1}Ub����у o1�m�����j�H�Trd��=�ٯ>=6���^9�p�����xcnvbFQ����oo1;ϑ�ƫL12���=�ț��u+��ì@B�le
ʡf�o<�߬��@ x8�#�0�]a 
��!s7�ϳ�9�� �sZ8{�՗��sL`�|�)�4ĥczOq�����n��	ק����0�]6��B���׻&���Y[���t����;j�d����T��W�P�t6d�|�zbU
��������4\@����O���df_U�B�9��z�V�B�s�,_�@W��y������Z��CU�z�ΰi�Nf��6M�y�w�.����s��
��u��xC�ane�K�3���|��-~P�ܥC�����̆�<D�J'��LKiC������*gۃ6��M��f��'J����.wp�a�r$�J��KI�N�Z����a�;� #��;�W
�E�D��+az�� j�����З��T�An�~F)[w�����a�v�H�+��UŽ�FD5tz���>B�	-\��ĸ�$�����{��+��}�TK��
���f��L p�Q�{���ωBC�)�a�Qӂ��taG�` -mR9ev&�{�ȱ�ëZ�񴴂���>T�i��Ѳ�a`r� �3</o(o�� NB������9��tu�� f{Zm�4?V�<6p;;�憥���w���"4����j�O�S�G��1|"����􏌅.��D������#��s���*��P��19��ȷ���K�r��<�ǄpcD������3�	��E��,q�x��"G��V$8Q�͎ �K�U�
��L���K{'H��s�U���$�2N����\E0�������mW�����D�m��� [uN�zR&�1�?�Ty�%��.�KM�m��}J��_}�4U���	VZ�e-�\֡��	}}�\�ᬲ&���G2���N�K��,:m����I�G��L���D8�j%�����`�x����n�x˟}Ʋi�ǋ�iD�������j�s���X#7l�9}�싨!n�[R'.�T����Yd��+�\^A+��O���x.¯��J�1���%y.|���fP�&�y��$�����"�X�c^$!���"�3Vļ�T��D�0J(T,t�G��H���ӡ��=,����2hRdt��݂ɽ�q�W�9`T������qE'�$Z��f�&@>n��	M8��Ɓ�>�3���tF�#�Տ�+7T��\��/��ۑ
LOJ���´�<HN���!� *�����e�������Feƾ"��|v�}[He7+?�Eعg���LW��^4+=�ạ̇}���Y'4$�l��,c����mwIِF
|S�2�I-sV�M�hN2�ϽR ����'8����7;w��޺.����LL~�d�!���\��[�̍(���\x�]c�5�)Qy����(iz|?&����'/�����i��T��$qi0O#�����_<�s�-0.0���O;�������Ea~��^^��V���? Y /��7��+l=���>��H�-#��'[T�f�_���K2�I��m���%%c<�hp�v��8���^t9��s���趺�`*.�´cr��D���.��
��$g��.�u�����z�=��&�8���+���@����v������]���.�*�e�((l�� l�������B���Q�[����V�A��~*I��`6�D�$/lծ��l���!�+�Yt�́�>��$����'�UnX10D��Ju}`�Z�)>�"NC
,�Ib��5����i������FP21�ъ��he�VA^=v{����|+�3���d�/0�Q�ә�~�M��-ܲ]jhi�A����C�����1�
%Ζ���%����:{�^ �.!�<6N4~[[�H�O��
֎�lv�ny�[�(Urp(��$`�}^=ꧢK�����2\��'�ֹ@M�gޡKqϊ|f)�'��q��T�r!9�C'���4::��dx��X�ݸ�u��x�W�ܡh,����q���Z\�т2؛�i5Z�N����ā�|N'��9����e�	�D���6H�A���\i�e(ެ�����&E�G��P����cD��d������#�#���V�9%�*0�x�oJ�H�|1�\�" $Y�YO�� 0+���K�h"��ϻ���W��T_s0���Uk��ܔl� ����z�����K5:B�L*�uˮhE�+aQ��������~�VU�Q9v��Ϧ�2%�t�+T�o��o�\ $i���j�Q��$!��x|��L�'���ם,�f����d� ΢�آŝ�oX��8n�v�ǧ���Pk	SJ�9*]���{��Ⱦ�"Ԩj��Tz�\���{FLE6!���$E9�}B�i���*ފ�����E�|�ҹo
��v�SFڳ�!�XI� Q������[����&��Q_?8�A֞�� @��C�ق�`\?�Hm`�$W�q�E���@<u��,=a��k�R��L8ed�J|L�y���v>#]���alf�iq�үd�6�8:�w\�*� ��5���ֳ�O��T ����i{�豺8�V3E*��tUĘ,%���'�3�����t��)_}���z�(^8�o�N4y4�"d�9c��.��l�5~)��w�y�Q�X�ZMnI ��x�dW��{��Ք����4�*�!��{�=��mf�z<		0Du1���S�t̕	i�r�l��U�TS9rV��c �(��� �j��I �BQ�e���Ot8�puVuLpJ���j}(q��U�y�c�(�����;��]�M
�מcv OO�a��Fh$��2�ˍף�_d�w}uC�o��K�����4)�%R��(�Bww��M�E �%]Q�����p�pm0��=���D�W��$��d��M��:�e,X`�o�-+Qrh(y8�~i,�H�� ������� 0O%=�^��s�MҞ.��47�7&@ﭘ���wJJ�wuÉ��j�~�X��se�p�p2��p���
sK�#c
;����Xꏠ��D���-F��m���MQ�j�&�l��@jI�&��&�.�aM2���Q���w��z���a���ug-�co/\9��/�꜅��h�y`,�ٍX�_A��߾���ʐ{��n�A����Y+�i�� ә�����AG:�-.��(�q���Kjs�͓�w�:��%n���Z!D��l��� ��S�"~,�����pR3�ְ������g�(1���#7��;���P~wBW^Z�-�7���x�|"�e�'M�����VGB[E��#^wi��(&:��/��8
���"�M�!vǨ��[1���,M��+}%Y�bt
_��=U��J0eM2m�5t �d�ZY����E���������slD�H�:yX�yY
�ˈo��Z�����u	��v`�?��
��V��$����j�Kt-4�a�uA��0"��&��t��|'c=siI}�z�5)�S#�p9U�a�\�X��D�\e{"R�=S��b]kFzC���?;�����C�V3��4"��`ܬ&�L�v_��r��Y�DB6$�\�[�6��r[� 9�4ч����toRJ��˻��h���WkͤB����_lva��ǐ�t�*�B <�l��:*Z��C��MZy��Dv*�o|b��t����"����e���/;:.\�ʝM%����G��&�%�b�>�1g�����l�e��A�-~��
�N����f�J�H�덣�TRD���Wɡ��� b�� Vq���6��Шzi��C�F.O-��]��d�o����ͮė������4��S豷/'�Z6`�
�F�,w�	��s0��z+rY*���ө�n�>�[�e�<)$5Q�|H����}�{*��3� �x�R��9���<B���f.�	�X�E���	~75�(���\,���,(� Ӏ�/)mhT�24���ȫH�@#���p�U�+��jx$��s*��������Q�C25w³�a��f"�LK�h2S}\`S-��*�D���2�L�ݑ���L�R��k�y�p�_[����>� =�\o�D���*�0RR%ջ�0j��n��Ph"C}�<iG$��n?o�xSJ1s�N<�C�+"�bJ��W%�T���jQB�kt��K����3|�����z����U;~�e�<���"�����ЈFB�����(�Bo'l��!K�.}`���:&�9t>
���y:���k�:���)j|}��o~Ҋ��cM�������{��t����L�i�	.`E�{��5�0_s#Qff�i�2K&VO�̞~����	������X�	�ņպQa~����> �8�HD� a���F0ةq�r����=Irͮ?d�N�趣g�f_���q'xs6��5��̬���3@~=Gjz�~UGv%�"�	�p�qw�� U�z�G)ŰC�|����]ks�RAV�	5ϤkY�K.9c�)��a�u��l�hu����f�%�����A_7ib�8��A{��t7�+�U@��T����^�7Ϧ����'kս**kH��-Pb�u�
�잤��j��(Z�u�@"0q�c�Nt���`�å�9�V������.�b�(ʕ@�x����4�*6Hr�9�������sRSPC���7���XU�2�A��;4l��IC>���tLbܩ�249��[�B�"e�ۈ�5;BeI0�۔��n��ј:RI��M���R���o%��Vdc��4+�z6�P�y-Q��n�׀p��K̑�l�.�r���N����w3�!6�ݴ/WnU��9���� )7ҝ9���V5U���l���MT?�Ξ�c!�y��f�����(a�"n.�yF�sIu����~�� /o��R�c7#/�����c����� |�o���OvL��Q�8�y_\�b9���}�-�ܚN�u��J:��5 �O�����_+�OE��M6�`���끰���~�Fd�4̴�>@��J��:��>��>�e:�嶜�=��;5�h���Y���B����W�o6}gC��%�:��U	߱�I@��q-����9
��h��;溑H�aN^w�J>�0rv��� �8&|ٳ�id-�s:&����pn�&��p�e��V��;ޑF{���D�':��<҅�&��zg�x磸케�����tvI��B��y���$��'Z�~h �V�E��\3�j��l-b{�^���%�5��������Z��ɂ��U�����1
?��\���j\8��3�ɼMw��0m)mgΆMJb�GLt �{�+�f7�=�f_�dh�J�T���QYݳ�@��Ct��;L�E���#$�Ů0��?�<V�+$/��{�/;e�k��BV~� ֶ�h���3��+���/Λd����Sޡ���u��^�� dZjq�����3�s7@uF�f(��s�1�+9����+!8���'8�kD{�%W�^;��ᇹ�6Z�ߐ�P� ��0�� �;�T�AV�ȼ5Ҫ	n�w=	�/�|$��D@�xڲ.'�6ǹ��ui���̟�
���!V*��8�M\����n6��}Ǥ�YF����e?��*�\�)o���io���������$�vq�BN��%�;Էt	�0��
�aE�����|�q(,�nvu�4�B�&y�#$6˴��%O#OF2�Cm�E���+����c��v���P%�e�w�����7����PV*�C��v�~U�O���1��A~��^Ԍl��?Y�]�/����y����ό@H��u���2W¦�A��
�I�?�b��v���`���&(���d<i�+F�	�K3plop�����S��$9/��q�P^���0�$�})��h|#�%ضleb����#�I
F��S9�ι�h�-�����kUM=�'S�d�!�l'�]e�[�K���0��p(�~��t�96/���Pf���F �
Yh�����Cں.��k�N���a��s��Bײ��^@��6f��Ge.��x�	0[�Aӽ�:>�(_�"B�*��^ذ�n��@<4B�я�����*f	/�=�8�H?qn	"�O�hB�N����$V��Q�$R��e���53͢5��t"����:EzX����=S��@�FJ�3�֢�[�/�5Y2��;$���������Q.���!#'��^��
��1jԉ�*\���:������2�V~t��ؕ�r�A�����\e�e.�]�Dmq�	_N�����w;B�.(7�X���qb�x��/~�0./M�E��@�����@�q�92vMJ��x�����C��&����!&�W��ҋ��<VNj������ ���HC�~��_����C�Wਏ닛��&�{���n�>\�?�ջ�^��D���5�'Zy��<�����g�]苓Lo;m8��	�U�-۞�˱&R��R�ǔ�X��4���L
 ��#np��&'|���^8�Χ�Cj�$�F5vN�Tс�:��:�o�-f/���W��?��yj�ԕ`�o'�8�&S�Èw��c�CZ*ǭ�cn|\�ͻB�(��+:�'�Ai�e5]�׷)GnǛҕ��@�z���)�1�M}&4��PK8��I��ؒ(�(�Ϫ�>��AC�8���W�F�SCu��2��{�-��-���z�����O<S/�KZ�g���
�tB��|�%�3�~�&�i���A�xF���f�h�õ1��%�4��	�{h���qmi6�w��y�͜��u�*Q��\��0��;P]H�m�h�u�#��M.^�y��YJ���<{e��rp%��jצ	�p ���g�}��ٵ����b!��{�oW<�[��[.��e˳�>r����y���g)4������U'R\�z�vj~]}�����L�c�č����]x�S���_"@�K=�mL��%_������o�q����b�~I�L#�Mɧ��ޙ @�Ħ��ZCC�; ���e;�x�%��&�U:[�z���e=u�}�%�a`���hd�@���H�)e�y�7��;^'h^W���8��Q��NI�G�Pf�m{���٠����=���lҷ�Z,"?�C^�ta�-u!yi��N1\�Q�-�0߱��E���~)��}퓹�8zV*^�&)����|�������K���u{�*k�!&n�"?'!��K�m����1��[##y��M�4|�`�}�7XƋ�͐6���;!��a�[����*hA��&����o3|����Gj4�?�����I�'��l �M���16��-{&j�rB�M�[\a1�F7�(��,�K���?o��H��T�=M�~Y��_��{�fa�c�����g�k������M,=3X%�:������/��l:6�^�g�<�A*�wݝxM���E�A�(�8���.����͜����'_�;թ�u�|֪<���)4����2�����q�N�.@Ƭa��1[�:J�B�!:�7�N;ń�Wi����X!j���:H D�G�ls}I�v��b�����a�N���W�7�nX,�b��)��%��n1~1�׀���EL��s�.�2�q��h@wEh���%zr;bp���[W�������:�7�e�y��h�r�>���s9C�3ؠmc����V������3��^�e|QOה�������/��#NTd�,���Է��w���`���4	$����fש�5��?0i����;�-0ჺ�zv�y�5�ea�C.�<��.h��80����%�kktV�3v�l���4�_R@����-ORN�sTg!9@��.Y���],�r������6E��V�N�a^�Z\�V�'��m�����~�fA���VQ$��>E�}7����KX2^V��;V��@-Qv&��1�	e�S |+�r����Gi���2�R8v��,�-���,�|i�y�&�7�癣�e� �#8���B]%��\z@���m���,�~�r.�����Htׂ�����E�F��;M~	����o4��m�v2����;R]��9M�?�2ФH87'nZ��Eo����0����#�ꨏ��}@+9*�����s����w�V�h­�jԩ�-�q�`����Cv8�\�K?_My◜76�ι�B0z���`��#O�%&>�j���������Y�(E)�Dഫ?G*#p�w����� �?��?�@�?�U��+�V��9	<�>4/d�	���0sm�%M������m�ӹ��r���hة�IZE��z���6�2���n��p��������<��1U��X]N��Gŧӝ8KۼN�7���gp��Q08�0x3����_M���P7�-�`(����(��� �D)v�h�  ��ށ~?��p��?kb�㻂�7;=?ّ).	�o�E�C�FɊ�6p�k��h�� �� �����ä�tJ�6�9�b�û��l��S��(ܮ	��#��q�<v�Ԯ�3"A�Z��j��7*ɂ _�5Gړ"��w2��n���*h��$�~)^����jB�������wa�^�P{�|��A�Ap��~F+�)c�m�>��V�/���Ǘ�ZS�����e����Zj���#U7v��9�[fN�LX�P��������z���x�1���+�#�eL��1E/h���rת��|�$;�A�,�:߉a�B�����p�V��|S�����`��	���ҟy��-tp'�Mã�h/�U��v����ѵ��|��ٕ�Ͻ�S�+`/�tq��~%@#���������viF�a��01V�Q�ԙ����^"6z"$�Ŧ����r��(�r�O�)R�8��f��+һK��R'�Y�פ��(�7XR��Cu0�P�4Lf�/�ޘ(.S�u��0�y�y��� ����
�t��u���OC�s�"Cx��L�o��3:�0	׊����]��J/�7HkM�<�'�F�帡�~tkȽ\����%�� �':<[v$[4�đ�G`#T���/�@�w{��*�ü�,��y_�6��䙪������Î�n���.�gc�8zv`���W״�۫����v��J̄��@�O	$]t��rC����2$m;��@��"c��x�b=4y/l�ީt��8�͐]�T b�0f��C��}�K@�5Ņ�-^�+�� �h]�GY�r��e��ѡ�F[	J]8tA�#|�P��բ����kR�`�b���=z�#t1�^k
�-EK���Z�,�� �Ϥ����m �h��Z��4��ƶ��o��8��i��A�\�����}r�8L'�8�R�e1����̝�Kxȟ�DD{�����A)�+r�
E��N�	�q8Z;i��]Yv�ED~O}�qp��9��0SI�Ȇ��;3S�����
��%��h9�5ʁ�~m/���ua��-���m��c�5C��uC���^�{Fhu���T����Ӹ#{�m)m�%6��tS��_ވ�m���H�|�K��'�+0"ς�����3H 4�LJ'5E/A���ܳi�'�;����\�����,��n55���WM�ڪ���:y� �����
˕2�5�.Ql�!K"X��{)M�ёM3���/7��c�.{��yC%L�s�D|l���-�z��PZ�S%ij��������#I�h�'���8*�ۓ4|����Z�m�I�ؤ�=�=���&wP`"�-y��٠QD r�E��'��߀�.	Z �O@
l�x�ꖱ�U�L�x�I�=��R�F�}-��6��)����f���4%�� ���d�"�eX�� �9s51�]�����֕v��Y�<�2��E�nXO��ɧLo�#�5n���[n�[�� �!|X��JE��������[�둊D�xU��햓vbO��f9���#\U� H÷P��L�cv-��A}����D���W�;��6�:v�!��"�à
`":�&�*J%Y�?�S�ֽ/8{5�r�`��"�+�tɿ��:�F�/�0����
�zs��(|{ �v�5l[�lx�e��' '.�T,�ǅ恠���(���:�=����q��.���!�Я'�'$�j��rԙE�����bGF����3[:C���J�E��T�:F5A�ju�ً-�)�-| �&��h��3;�����-ğ��D��N�E;3[m�J�O
z���E��{�5N��3d�F��muc��������Y�o�`~W_,V�1<v�i):������k�{on(~�7��z�`���e��,a0`t[�{��M�4�B��L0���Jx�.�Hpg���2��>3�R�J���f������hT���U��U u5����q2�B��HSÃ��3����ēO����ZA<j��މ����-�n�]Y�4#ΛIe)*7Q�I� �A���c�v#�,��̋���@"�b����M����R�揻��rv�(t��;�
��FV�����b�GJU�6e���n���%��֖!��������u�t����lQ��/G0f��{��SR�"[Q��I��M1���u�'�.��@w;r�����&X FK2Ǖ�n�����d�x��hY���m�Aw��٢�����|��4�KP��˶�#\"���+AI5��LG!����_�,��G.��[��0Ũ�/zsL;��&6Ȣ��9&���bm]
Vy�k�S�Z�6/����h㆑��%M��f�X³�i�'���.f	��L"�|f_5Y�I/m9٠kr.��ѳB���|��P`�?�`?2�EV/c�S�]�z��$#gY�:����{��J�g�<��MAs�%+��XJd�N+���3=NU�E�!�Im�d~�Y��x��f���>k���ݑ*�g4`n_B�ͣ���^���w�Z��7W1�ts|��PE��v�8����%��i(�Zs��w����ǹ$e�.虂$��U�*��_6��۱ �w�P�~�Y�o����~E��̙f�f|0��~	&�F���W��|H�l��+�lz��+��\fTDia��vCQ��SB�&SQ��p\��0֦����zC�gN�9�, ��Z��N���#�������#n�?c�M�73�_�����J�ۨk	����������1�}q/��1�g�N���\�h�L�j@<��Y݋��(�D_T=	[�����_�˝x�cȤ@���d�� >��)��W'h1����xj���2!��H�q�W�6�')�p�Fޅ��b��9bW��;P��KcǨL�����"R�(��\*ii���J�CS��R���P���%�Sδh�6���(G�����C&�3ܛ�h!���B:T��lGݕ���_�az��%cot9� �7�xR�M�̕���h�Q��x��'���w��vt@׍��������l����F����A���d���+�ʤl�si��R�xx����MS��{�W�ם5P���Me7�|t|t��j�����v����8=Ӱx���N�۹tى���_�	^щ�/���[��v�eIüoˑg��g]#�WP
+�ރy��[T*]��ۄ��oY�{u��Ew�F^�
L��2�Ղ�5�5�Ld���ߖc%]��g#�!�A�իI�yǀ�wP�S�gd��/����V���f�ߤ�<��Ϧi���LZT�K��J/u�#���q����n<0�%d�4DE������P�f5��\��h�#:�՗Qq �ce�(����;[��g:�Xcq�L?�p q�U��f��^bWB^ �:�"��4h��>?���*����}�7Z��%��g��� �Ԉ4 Vai�z����,,��}E���')(���6��cCD(���` z�� ��q��fgl_O�bh�x�ꐻػ�>-�д�&B�!$�W���S)J*f� ��Z3l3�����+2(��D�遌���"� *J���-����0���7��Ş�SN]�|�
������(P�z/���dRGhuL��� 	�ډ�B kD���lQvX������<t6ǰ��
�a�����p��p�k	;�#S�2:hk�ֺ&��-!s��8< ��<��H+A�+�UW�Ay�7߇�8��3K	jd�I���ԥ��hӞ �pO�S�z���y�M�ތ��e���~m�}R�����*$�����v�h%�C�6�����7v���_	�(���l�И%�6��Xdg�M򷘸�K�Yjx�s�d���rw�?GI������cmx�����D�Y�*�:F�<y�	���9�&So2d.�"���8�h�l�G?(����N� p`�C��=	Ȓ��y8��T�V��C"�#i,]|���l��gh��"!�&�(�v��X�pE���~��T�������i�?"j9?�g���EN�"���+ɥ�0��D�y0�M�/@�	�4���)u�4S؜*�x2G�z��k�bec5�QvO5������F��
TѤ�����.8ճYa��
� x��7ތB*� ���k�~i!�>�aeM�*~1Pѱ��t|k.O�ñ�L���f�� ��_s^�k��� \$�`�-���r�A��N����m����6D��?綡*hA�^*s����^}_�̂�	7�͋*��]�jN���bjo!��7���6���2�!p�o/���=!���x����)8���ov�+�gy��>�o��l��u5��I�b�s�K.[iܳ��O�b��^��K^@PƁ��!~��$@���A��J0&�烡�T'g�:��7��w���L�b�k)dȓX<��R���������)����R�S�|�ME�����k�j��+[����QJ�;�]�4��J~�$X�C.6�W���s<��N5'yJ���d��P��ݯ��Y¡Zv�V�N�0�'\�S�߆vh
���ltG��Xs_@sM����e+�p�?��F�G�=eM�^G�/�n�!�`@�qZ�?t+HՖk�t��Ex5��o<�06�m+����,wO)%���5F�^$T�i �X�d[d�#�Ѻ�ވz�k��E�M�,����|~�F��_׏8�<�<��0�W\�0:r���t1�+����d�@[h���JC	�U%�@�j"�;�9T1�~(��f������>�[��դ1�j�Bu>�������A����/���ĳo�5�RWnVپ�UO�C��!0_]�6��2 ݈ҩ�솵�01>��C���~o��ί7��ؚ��9�v��{�r�p��N|���3����@9V�pc��Sbuj{����pâ�Ƈb�a����N� ��|H"'�5*��{2�!��p;���4	�V?PO2v�(��7h���c����MIH7�ή-9� �қ���n���k���'��\G�$h�֗,���c;v(J
%�S+q��<�j	&L��l���3���v-o�[ɢc9��U���k�lCC#U�Ƽ?�AK���y�|�V}�μR���B���m�CSS��Nԗw0�4������( C���`�;�Te�M�Q��d�Ae�IC��Ь��rzܗ!���c-�	����8l�9�
�H�[`�����l�[*�4��;\�C����ܬP����
[� �N�D)�	C���@����,o46�B]��w`V�õ�yY�x"��6����g%����_w�lӝ OP!�[=��F/�^�Zs�O�����,��W!��법��[�n�zڹ�ʴ��)���듹8\�k���)?���K��W����&��\���:�`A���9	���UC������Ln|�]N@��֬�Z�Kh!���
/`�&ld�S�OH	�+�U���@L�_c�E�\��Mx,j8�A�Q0��ڢ�ᅉ^W��8�ȅ9PNi;G
V�T�k"�Ʀ5 򒯾9l3�q�	k�$�n.�0i�`~���(��/�I�ZКG�2�,W\=	��K �J`y�}��"��(��GkROF|�Y�h�t_�Sm^O�+�M:b�#c6��E�����~�
?T�4����5����x�M��ItW�|S�P��ݹ��M�<�󻹂 /MU'�U�e�*;H`��bqu8�5^��<f��gYR˅�md�\��>�4��T�<����%'�T '�ݜ؄F�}@��If�l��(�S���#Pe�j_�G!��#S��|�9�2ΔQ�O��(�Ʉ�	:�Ib��k߁��	��T֞h�`J����ⶸ�R	f�|S���
���a��8�/��ּ�.��>߮Vg���v�1_���1��U{�uq%Q�W'��"!5�hw�D��4���ߌ�+�rƙ�+��3�����V!�1[,�_�=!ɏ�k�ܣ�0�6�v����]{�;�|���������J#4�T5�O �W+e�_���W��Qw�p�M[�3[�,��ʰ����N�!{�A���zB/"֏��5`��Уb�`n%������|??�����Gn�a1����/�G�n9��pp����z���A��ߺ�]�GK��w����M�c� ^\��B`At�D�>�{�<}�(�}>�n{�W��s~��Y�]]��D�፞L
2Xx4�Qv}�}��A�$��k)3b���%�����5`��=�ˋ�әz�^�i�
Xm(U#��>��0��j�u�
�N�L��ҝQs ���&-_���k�xU2՚r"P��Z�i� ��~�ry3�A�!��"�.*?��1��r�3��d�< tU���kH�&��WuI�/�D��_���	Zz!ŉq����FP�x��"������b�d��Ar5Z�5^��f�̤�H7����^��w��G�����&���T�;at��%Bx@��	�v7'+��cT�W�������1df@�}�"��Fbx������e՗��ÕAנ�R���2^rh0
`x�~���yw�^�.�Y���D�>
P�)�{!Bi���J+��7�g�y��J�ł=H�g���jf��ʺ�-��3ˬ����X�|I:?I!\lQ���=�^ƫN�]���ܼ |0��)B��{����]�Nf���
~�5�E��iXD�^Zd�7�M)���B,�c�ɚ�Gk�'��>]��ϲ�Ԉ6�2��Y�e����UY���B�X��8�3˄�1��G�ͥ�����5j��g�Fnxr�1�{�N&e֔&ku�N�c;�7e���JIM�<����)��[K�����u�����#�e �#U����P�Ʉg{�7�
K�?�pO�!`��=0|a�qZ]��&��WD�E�	�uD��cY����aT=U����pt�O��R�$�F��U�ޮ�L<��ዩda�t����؈��S9�Å��̊����)3Eěq�?�
�`�j�-��}�<ŀ����:�����Y|	�r9��п*��.��M>y����87M]�=@E�<� ��p��O��tt�q�b�JAɛ�#����еٳ9��.�o�h�Um��$JX���F.�[R�0д%��1�C�OlD����/W���j�J>���$;���a��6���$ 3z+�*6��!B�c�1Z7�D��t���<$;֐$��e��uJ�xsZ�~�q�֕+B�.@G^��	0.�*^Z�t@Vi�U`TyHz�E�2�
��s��)� 4�KM�NkZ�#bT'J;D�⸥��Ҟ�
���]��O�}��bbdE�1Ɍ��w#���on �b+>^*ʱ�?���Z�љp���5��w��MZ��W��<���_)��p;����pe�J<�m�,IU3TX>��J���S��J m��S]g}9�Mk��G&2�&�Wӵ��Tm߱\��w��.0-�N�� *�[���P�O
���{�W�ؤ]�4$���!m}���(�^ �-<�]t���d����>��i���~�ۙ׊����!VC�q�h���B��edu����	T��r�i�]�������u��yA��X��:#%�����W�&�	��� ����>u7(?�"�
�ٍɣ)�����L��ᾱI4h+�w��*�mS�EUt~Y�S��xZ�r  �St��oRv��vL�������?�An��jn�>�x8	\dk�=�����e`A�7�ru�wģ;�&��Na F�*Hl�QN٭b,���2�
[[`����c�����sT�ĵ�Mf�y�������;��Ku+��3������x������R��Wͣ|�S��t�Z��[�_�$�	|�w��Y�����!����)k���40���E��K�15V�c���R��E��7��62�᠝��b�ybY�b�YȔ+���L�P���}O^��Ȥ�m�"ר[����M��	�,���˄2���� O��׌m� �@]{KN:\0��^䫜�S6��_������*j}�^��J�$�x�`��	�2U�� ������N,���_���C�Q��(�,OV��,�&*�?d;/���}a�6DC�!�*ߎ55�?請�Q��u5��;�(�z��`q��}o�J�3�0.1s����{��(�q�3��&zG��N[���Nݞ�$"ȖTWb�'�wD�������QS����ȄօK��=;?��7���;[��O94�;݂r�dV�D�8���_� �%\V���I��:��n�-���LN��%�F���c�O��������1�u	�T{��:>��j��|�֞a΋W��-�1�򂔙�����&����3�z�FY����'���蛭@�-�:0C� �+�h��$;��E9"i�$g�JY�ܬF�\Rx9���諈��e��2�O�RS�~r'��Qz#���W���م������� Ό\k��o�2�fa�ij%2���&Q�i�4��I� �� =�Ƙ
n�0-O$��Ҁ$���:ˡ��$�O�G�Yo�UxVpf�Vtn���H�}�y ��A�T��E�#���y�)�{���HwC����Ң��`-h�?E	���CU�-Cn��1A��J�"r(���
�a0��ɜ��I����!�ū����p�>�Pb�����H�q��Z�<S|��_�D�?���9ԅ�ɀ�bc[�6�t��9ZI蛁�m�H{�.�X4}b�-ȱ��۸�9�����^=�Yx:�E���,±�g��H��7��~�&`2��V�����Pf���E{���;�Z%�������W�]������I8��I�2$�흑rp�Gf1�(7C�	�4��"x��Y�(��9��[��lBO_�݉!�i��'�[�������r�l%},[I	�OV0hf�E��n9�@E6A��>�©�<%wZĬﵦ9੔S��u�K�@�^h�k���P>R����_��%:i.��Y�M	�a�A
�w��J�����a�bjbo���<���H����5Wk�/�}Ԑ�O�O�|�c�a�BQZ���{��Vٛ�g�5�2^1�Q�q��'Rg��@��R�r�O(�����MON���X�WX���~�iV�/�d����]���+Wp����B�ׯf�R�����n��d}s��k�CL���x���{L��b�/I$;��?,�����L�0�O2q����l����vC��_�(!���5�{h����տp�M?k���5Q�hӈ�Q�ҺF#��{����
�'���B���6Y����eo�l��$ci�;
�.!�ĀK_,��og�3�4�M�ǋ��K���}U/�d΃y!0f��ѓJ�J+Q�]�"��=��枳�iFT��l������r �P-�pY���i������]>�AFnqL�c�fť����4���^"]����ԏ;ا^��
C�9�-���6s�B��gPe������˷D_�8����b*��@R��)U
���^���iИ>W�:׆e�D���>�P����?���j�u�)}MQ��Fs�jZ�(ע������vt��-`����I�/�z;�bٗ}3�s��o��ઠ,e���\��"�太�%*�O��ʤ3<���+�Ȉ��az��"�����;��~��#fT�J�~$�@������=���������c����A5in�<#�eO�
Q��ؐ
/%@�bsV>��$~��@x��O#�:_����H_I���!P�Iљ�q1�D=�'ti��f�:����w����z����2������xk��8�3���������&�2��#�QL#_p��۬m��	�VQ�x�ڤ��ë9��<�tY�Y���>Z%�oa4]5�4Ij�h�G�T铍��B��ǌ	���΍S�{NB>��:��k� ���[܆g�Z�W��]N��Y������wF����`�n��s�'P`�<N�R�P}1t=nj���"/T;�������X/ �lݷ5n?�������=Jv !Xp1�t[c�f87��(�/���(u1�h�]@�k�.xhT��w��^��]�nlȸZ9>�QB����vn���V�*h^���EʁK�$#}4�/k�}�X��cڃ��$��m�7��^�����>L@d��ϟKX��q���4��²�P��Ѩ��%�"�7�������~J��{H-�|�~.�9��A*��[E�̜C]����3�ER0�h���o��?V�.y�u�k����+���=���:�'��[�a�s��P�[dp�m<*�����L.<[�
��X�!M_ �&A��a�¦��^}�)ؠu��3���:I�����Ӫ~愅 �VZ��8�|:"����,����}���u�c/牏��|��y�.��.����-S�b��s��04��J5��������l�5�I\�EGGg��t4���"8-k�bw��X���"3'�D5���H�=`�CkR ;�}��΢�?4��m/�K)�~�^޴_��Y���[P�X(���P��6]� �/�w�=G�?��[�L�9�A�P [��˛�$��+\TP���O��z	R�R�I���+z�τ�l3�/s����~>]l#C�(Q��:1����WE�H.�7`1����*J�/hĂs�xP�����o�ps��$?�Ĝ�=�`K6^y~DE�>u�Lp1r
���{�A��7J�h�x�?��3�ϴL[�&�vK�#���$��sM'�T����nZ3ܣf,�Ƶ�h��A։F1� �c�ٲ�О��{i�(���5d�>�y�TF5��T�;*��XD	��6xl�;D�`����N��'t"�R�8���oCHI��Z����EU�im:Q%��Q�X�T�����e7��}Wø��u�.��#<�gt���D��а�N'[Ϩ�1-m�~���Ƽ�Jo����1|~T�?�'^�ћ���4�H��4�6匛/ő��xX��,����j���;ܗ�l}��i�Am��ܱ��V��q�w�{���!��z1k^H;�C��O���t.��<�rwH�`6m;Z)E6�7_�U�۴�k����2zK|A���-�����9��;�.�� ���Q���v:�B���n�:Q��d��O�;z���85�.���'��1COs��C!Y����3�7f���R�� 5��?�L)K{^�;�����Q^��Brَq)�D���}t�ɩ���z��X�D����mg�4�}8����Bvr�]��z�����P��#_Ȇ�)�[O�*�c\��#Y8e���������������)c�}g#B��`�����k{�vN$SM��l��V��T�u��U�����$�����5���1bQ���JpF����0Q#���!�]�xV�E��<s�
,��/��XI�n����t}��zv(::K�WjT9��{������&G�u���alh��^J�\q���m�xއ�g7RbS�N\7�SX���	�1��-ۆ�\g�OE�$�)��Hee�D]f��֥22�F�dSO���ɰ@�e��>E(�7y{��lϣ��1��2HB@|SQ�u{��X��6��{��x��=���gxc;�Ơ�>�j��x��%"˻+
P���^02�q �����b' Zj�?��9����_�����^H�%K�ބq�Ծ��xI}p���������۾���^F7����`�3i����H0�7ch�p&8�J�)X�p�V�h��Ϥ�4�:�yPB8TK���M��X�w`Q�j�o���͖��$�J"�rA���ȗ����JE�:FF�$8 ���v�`>��;Z%�C=*IX���h뉬o��9��ϕ1��_�O]&�L��y5+��U�O�����捏�_K�Eɻ\A�*��Z�[�Ŭ`�)�Q%+N˪��12�����N$�`t�rI��[�����r/��˟LvN�Wec��%'�6nÐiY�!��צ�s-�-kf��]�}�	�U^��	��q�%�cFL�H	����j���TS
��T�M���<-�+����cf���NV�����T\��S��i�樔�Ԇ@��E�ί�L�xE,3�O7G�����^�n���6��C�.}��6��1X{}�x�j�"Lb�������S�"v�q�&p�I3����.W�ZD�[/W��*��c�d���m{	�x�-�`L.��dܜ%�{\
��f׽�Aب2~�D�K��7�ƅ�z�u`n��W�AJK�t����P�X���n�[TM�~�5���bg�������e�pn%#:�3M��Je�n�,��x�p�ݔ��C�x��MJ�,\X0�L�>��
����=���i�-�a�]Ӕ˔�s���`9���Q�^�[�
-
R���D����w�ی8R|�=��k��(�&]�@M�0:w(m=�ǥ�s�����Xˊ�wq\�ٖ`0]aZ�0�70�y7y�3������yM�q57���L~{��J�f;{��4�a��C�C�M� [u؎4��r,20�]]�� ���wd�
>�+/��Ö��-�b�ă,`�Md`d뺍fr��C�a���wq��3sw�/R�sLo�`��F{�f%6f���s�-;�b��9@��w7û�ڇz3e��nϾ���Zn�<��W�)���C�m�������.IY%-�5� .�G���ܲm�W⦟���a����w4i�v 1��x����>�&��H#��W�n����;[	��-�n���yY׃�$�7���}ÒfK�C�d?�?KB��T���-#���[�]�F���Ǽ��My��+եӄ�M�<�gy�ru�A������P�F/F`<!��\�'@ӧ�i�A+J�i�}>wj��\p�?�,'��F
afKr�B󱷟T�<���Z�|�qUbF��5yt���Wєw�\��������=��
C�j]�`���Ů�[�~�e��c��(~W�a��x��e�΀�lD1'ߺH�1~Z�]0#������d�
�p
$<v�ޢ9�����OUo
��gf�*�w������N�����2�L�O������Թ5���	��buB����^�Et;�}���c��m�y4-Ϯ:v�fင�YM�]v��&����hN q���T��P��3N�O�µ	�1�qķ^����`�q����R���X�oN��W�Q�ݾ����"E5ҷ~Ҕ���Ky��i���|93��4@������ڼ�0����]a�L�����>�R1��u�j�Ѵ(N*_�郵���}��
RI⮪Iy�~r�w�>��v��uO��%
�͍C3�)i��d�6=(׉g�<�Gﯓ��4ع�ʃ�4�Q�ѪX��i���g"]��-v��mK�CQ�ޱ.�S�Q�y�������/%S�����7	c{�(m����)C����s[����}-���p�λ���M&ỡ� Qթ��K,�w}��ʜ
r����H�����E�������O���݁�k�R!��y���t���I�T	�br�)]��$���@=�v�L�!#F�y;����N��WA�ۣ�z*�M�ߚ�jQ�L�`�8gf]�u�H��#�N˭��nɎ؍�����#��قX{�8^J�CH٠���ɋ7ӣ�䢒	*<����ĳ��e�r�}O3�1�������fڟ����nvo��O�}ي��#8���ﺺ��B/����z���|A��P���b���+�4#?V9�;���I�i2E������6��~�o��*r���_�����67��ۨ	8��A�9О��Q�?y8�������/��s��0F'�y*��N��_c�c��w����J�{���#ǭl7ՇA}��K[�n�&� `T�C�K���E��ֺ	��皬�_l�w��#�j��}k=�Ƴ����O��#}�\�?$��"��m�;ͮP$��c O�,�2�M?la=�a��x�p7��Yk�~Z1h�&w>5���r{��%đQ�@Ml���g�hChU�����(t��r]2䘝E*��zX{�4�B��?J��r(L_��Ɠz7�sNɵYT	����˛7�V�����Y������ D�Pu4���"�x�B���o{Gy�a�u`JמEQ�������j2��4�d(��3JK�z�m��S6�W#�h<-,���Os�owd��=wz�
�@&�l�<�&�G'���h���W���ѻN�UM�y�o?�w�g`�t�:�M���߾x��M�.��v2Nğ�l7����L�Q@�n���n{@O�����E����D��g���Eg��H_�C��V/�ď`A��wJ1/| ��(c閬L}R�iDe��\�nv9�X7 x�"��!�^{A��
3G��-�P�n��A�K"��y�R�S::��X���<����;s�R�R^&�l_˰c��$��>VR[��u�,#���b� ������C��=��(�p�	�~���'�Kg�hvtwO@��T��'?����1�{pӑʸ��I�|e���*4�E4�RR
 �u��I𵇯D��ݻm�dN��L|���q�A�(���βhs)A`0��޽:D���w����S�he"��֢1��Í����V��!Khq�!P�Avd�6i�'��;�-�㉺)�B=i���Nr̿¡����zֹ P�+i�v|�U(X<��J�:@]�o��Y�c=�ON��ehs1/�j��eB�C8���� �wo�b=�2.�P�"qM2��l5`�l��n[w�.�n���\H��v	aC�9M���/���K#���$.�J�s)�qǼ�f$�*�%*\���J'D��s��[,+5����=�=+�n�:,�}\��7�@�$�h��~T�Wf�9K��bEi_K^��E�u�$�X���AR^��-`�k�)Ԛ�e	�TVc�� �)�� �X��'��X�^
��j�`��R#��ֻ��7;�C�DC�K��jċ�vb_d�ok�	�z��s��ȓ���poE �z8�G��#<�4����*VWJ����r��ۃQ8��Ҽ�;
ȳd�Լ�x�;�n���v6��ym�)�ɉ����u.]}ͩuU1�_f
���/�x
�* ����"q�_��yv~�ӪS�d�����~�@����Y�ڋz�Ʃn�ق��Z���>z�y8��"e��3��Yi�O�3\�F�41C -�wi5�<���9I{#��9��T���]�XbQ(�t[�Ac�#Մ5��޷����b�uT�a(��p�1���C��S�LO��)� ��V�<65���ުd�XY�k��8�2�AA����<>d<K�]9&�Z-\@�%�ؠ���U��j�jX��3V�O��@HZ ����2g�/ �2�eOxۥ��ʒ�KiC"�z�ri�C9����J	��Bע�����+'b�>����'����-�`��F�َ|���#b�☱,\�y쏄���y}ή�H�'�X���	��	Ƥ�B�MN��z6�����ߞ2#���1LfH\1����Mh�a3��K���:�g��x�୪Rt�R"J�Q�`|�g���=�~�=���_�RGYbuy��_z❄�������e���JU�Gm�!X.�a�\���k�ґ~�y4N�9�������{�q:t�^lL���� �d�a���C�W�cY��{���a���?Jq5�k(Ka�81���)d}Q�ɿ�T�5��Í��ب�,m��k�)��Qo�;-�<L��Ou�c��2�� �爆d<m��p��1�-D�P�0k=^C��{�N�ϋ����uR=W=*3�('���|+
�� x��gR���(BŒ�%���ED1�ߐbH��NYsޘ�E���24i�3�����Lz��djB����e�"������z���e�\yʖL�qپvK=F5&���v��Ba��sc�hXŲ�����0�aǎ��w��e��f@U0,Ă�E���ҫ�d^��?��XܕK�<b�A<�|�)S�$��-%y8�>Cx�g!�S��O���j��9�m��mh������q�V��k�����4�?�)��f����o��"��ǩ_�/IY�*c%3b�PJ8��:�b�wC=9��BM�\��tP�n*
��I6uz�$���n��U�o��E��)'O�-���*�ϴI��Zh)�xI��h�����i4N����J!�A�m,�4;HEdy`���Mĉ�;IsG0� � o�|X�=)j)O��!��)�l�sa�ͮ���ݦ�v�dM>5a+e���B)�Ȥ�^`�wW3]^Q�G��[["�E#�4��ƖTq��VG�s.��gi���4�K��Q�ͩ	�H ��1���������_��l��Tib�}Qk�c�z�xy6o=�*��eLm�&?"�\�k� ��W0��F˸�A�lܱ���%%\T�}_�|v�=T_��C�2��Yii�8���)_1Lt�N!1Z��C������1eW<��U-eef#jo]�x��5��p��*~�׀�c�9�'���O����#��(>ڵA�Łz���:�0�L���>E���3��@�]��+��E�q�k��k���'G��u�NSz<<��vpL%_���K�UBa�wo���Gb��h�:�B"��� )���_܉�<�K���Z
/H|���_�r�~B^W@�]/�S�)������ �m�e K�O	$u�\_̕}���U����\g��
b�+�r�
�p"�$�+~�P� �k��5�d`�m����� 1��{��ӏ�~3��1Ѩ�|R� k9�(���0�9+ͤ?��S�
6�:.� �
W�`����݊˽Y���5��>��U����U�t�`+ �\�M"������
z����x��%V�2=����JMٗ�(H(x��^o�M��|�Y^�Cf{��5�N�u�yS����۴r�wK_���ڠ\~���DU�L��]�k�볠�~9��tR!�F9k{�]?�BQ�6�>Q2*7�,~����Ӝ������ݪ�9�=�q���<��ݶ�ɚV @:q�xLG1S��E�R�4�R;D�"f�#�@�	-� |i"(ۆϕ�J�<�kb�J�ݫ��y�c�L�%u����5��}_���\�=�Prۿ� �'9�;�����kE��|=�#y�M���Ŵ|���Xʑ�1�O�8����G��J���üt�������hХvP��i�.��n��J�&�T���)!5�1�@�{Dw����}E�U��L'g/���C��XR�2����- )�܃E���_k-�}_�t�r*��μ���(������"O(%oE��M 歴VnTj�_������*C�4@�2����P�'2]�*~�ͩ��m�(XH@�F���`X�:҆�������v�]��9�ik�A�����HsV�v�iy
}͝T�t�Ca���N}�{�:���Y����c�|����8qVa�5]ᥔ{��!���hJ�g��Ʉҗ^��X�gh�+,���`���g�vv��(���yY�՘���Vm&�=��?��h)��Q�,�Mx@d�m���*�Л���n&�H��V��(�"�>�#5ƾ��R��o\J��C�{�{pR�jte�)ߖ��Ă��3*�.]*]�/rY��ڄ��m��Ns^D��s�b*�oާѺ�%��[�	X�=��08*"V�e:��a�\�{�?��-r�ak8�$�7+"���w����������ȭ�V�
�C��-��T�h������Cm���-҃�,�b��Q�f��l�F� \sٲaՄ>e��r��'+�1'np�|���8I��kD�tE���Ts��s����0zv���bRz��0n�z�q3��Y�qc�����D��!t�7�b�-���렵��GEK���	��Ձ1��i/��_�
f����H�vm|���i%��G�dѮ)�v$�MsYf+P=5p���,�u�4u��t�٧�C��
�Q�u�gs�J�Hϥ(�ATz8$�)��wlm]P��� ����
�,�欆��'�?s�hv"��x{2uciЌ/[R[5�<J��Q�L��@�$AIB���̔q]��Ɓ��G�_B��^�W4��y�S�['�{���٨_t��%N�F�s���S*���`h�q>��Q�n�@���rN٭	f�t�߁�-�u5q���/�J���, �8�k�������G����)	��#��f-��c�!'��.�a�)3-�@��Z���=�b]��Ƶ(�;K�"9M����"k9Z�ՁLuxP�C0�VN������@��=�Ն��E��)'b�b�Kp�"z`M(�@D36l��o�^!`ۋHq.m�_�[{Ϸ���?�9E�0����穨D�`q��4Z��Y�O�z���;�=v7So��^��y.b�HS��r|��h�4R�=	Yq��Q��9��2�/����k�t��{w�'���F�-��B>JH U��`�t�����1���΄�|[�w�~�����n���n�Mm�wx�>mkd�x4�q[n����X�u��+�Dׇ��擙���
�97oH7F�K�yC��������o�ъț��T+������L+��X�L|���]:�;������%�.�������b��m�Iz��1%��6���+����%̂�4������dʐ$:0�7q�
-W]�V�ߧUǕ�Y���9Z���~9��2�v�<��'5u�,�I@��3Zz{�&�t4�@D��	іR���s+��?B^xW�L���Lԡ�h�ӟ���,��B�݆���0cO��MJ8�p�Su�[�ӯ/׹^ޥ��g������#��x��#��.��NSa¶�~�o��c��Ŧ�o!��im˼0ؙ���­!����I��̽������*�{,��p�jO�E2w��n}�gQ%�����E�Q�
�S={;i��/���Q���X�I�@`oS�Ɨ���{��Cg�-��lh�F�5�6'�2o�M\,��̱�����z�XkU.%F��ީ-5#���RVÙ�&a��QN<0nG��4V;Ld����iV4�.kM�;�v8j�S��5 7u�$nƿ��>6�N�mD�-Ġ�y}�z�!�k��s�u�`�f��/K^�D�4j�ۨ�Q�4n�@v��z�$�hCw�JP�$;�.ka�(4oy�Q����M�
W���5z���}{ecvXl�O��$���k��Ն���>4����q�����`]8]&8�\}}�����<WΎ�v 6M9�Y�ŉ`;y�uT�"�6&����ѥ�%K��Dω������w�״ =�`^�ʓB�4�5՘{�,:*9UŒ2=�U�r��e*A��ZrNjѐ�Y��&7��c��s��SW��n���B�-N(��yAy)X?��+�G|C]�C��Y��V��SW�N�tK:.�4�hDY�!io���qK#��n1˫Է��f�������L2F�|G[�.3L!"�+߉l�M��m���M��c6b֖�qx���$#H�ǖ���ו�uR8#���'S�]K�Y���W�Z�߼p�%��Z.S�-,*��C�R�W�9NMFjԤ�#�h�/���;%k��IOdN��Fy$̸�L����D��J��X���]�"w���f鈵�ވ�E�*�O��?�Mr���`�׶��
c>�k5�v2ګ������E0|ZTH�e͂*��l��ɋm��������iE[���UaG���:<^g�Vj�;�h7��Ҷ�c��Z
C�BE*�E_(�k�
�=�	�J���H�t�j%��oӳ�� ��m��<l88�����j�&����c?��ҲSE	4͏x��ߗ���:8vЊo)���et<�U��gr��0��+g�� �[v���	�04�nG~����8풢6����s�GOm<���㋢���Ra�M��R2̣g3Æ��<�`�od�Vź�7��yvx�H	���a���x өį�K�8E� ���-�W�T�� 2
Of��î,�X�p�i���xtQ78��'OpJ3��1�����&j';<����J�u�xｗT��	DKv�y%-�tS,"������R����V�Cl�|S��G�B3@i�<BbM��F)i�Y&H��^��1�4*�������>��(�����L����3�s�z0��}��t��-�_�r�&
���Ə���-|BW8j�
��?S�Z��A�Y���r��������4�Yţ�>�X�sʗӖ]�����+#*��#�ۭ�%�:��'M�{'ȯ�8g��S)�b��tC�ڔ��H�:�}��� �>Z=Ѹ0��g({�~t͡\!Y��\ͦQ+�>&B�<��*n�54���w��ڴ�C�Wc�����lG�h^c�ӓ�4 27���h�ꉧ��SMa��vy����>���k:��FLn��[�������fWQ��m�% ��P�Y��j�R?݃00"�6X�f�1���r��eŝ����0�]R8����c~NMQi!ϫz��&�:�89�}�	A3�8��>A��V˫�@Wx�=����JU�س��2��δA�{�;�!&/�؍�r�[*�+d���Ip��t�
J�@���N��[�co�<O�(��1=�YE���G$����}�����7 ;t��b�J��iq����\����~�9XG��~o����,����{��4 y�Zoӈ��l��=A.��s�D%|]Z��+��5��E�wKg%��6:�٘+�4X䙂ߒ<��G %����Ml��'9���Z�[�.:3��r5O>e3�x��=��w�T!���_͸7�}�6�WB
~�l�56�}���NVEǼ����'V9D�s7RI4t>%��)4���%�6�,��)���,�g�1�i9=�h���lY�忊˶��f4�9�l;8�daJ�y�P"���Ҡ���շj����:""��aD�]�Q�fUО����ʅS �P[����1_
�O�;%)�<�����M\�80����5�s�1F&��̜�%e|�rd�ܷdA¯���GE͟�]��F��~W+��?)���?�W��WnP��vΞE���ʹZ_]����	��U>��d ����[���1��	V>�����|O�mL�f:i�5�i߯�݃H�� /dY����3��9�G��`�r.6���&�R�D!@��R�{{�TZ]���+��A���ps�{(�ഠ�BvZ�c�Qܖ���	�������S����y		'O�Z��^.�x�-�i�	�V�DA)U���a:O���,�������"�*��Ҙ��@��O�%J��{���-�F\%���TҠ����'�������؈8ޑ�%h��*fgv�A(ںc�����r��G�禮핌��a�Jb��.IK�N��l�B��U��������㶈��tW��Kv��U�x?ov�5�\7}gד�=9�2T�㮄��|�?<���"������s+Tv���onn�H	��$aÓ�ri�������~���6w}���j� �s	~9wZ'��T��"A�?�"��8�D��]��t��1B���LqfɋU��S5��V�o8^uhy0���5�z7��Ļ��� ������ȼB#n%Pv=��p�˨�)bXi�\��*�Ĵ�䙴�)�{$K�t.����מ��zN��fel;�"�1,����F#R0�-��CBܙh�f��O7���k�N�]���Z�d[��E��0jd�i��YXWv4|��m��.�X\��ۯk��`ɒE)\3�L�ys�5�;�)og)*u���
�c��k�9��	8�]�r�l�*� ���Y\�	���.�nר@�<��t�]�_ ��i���%f��M�l����H�4V^���^w̎͡8�]:��gޛ�Mhϼ2��M�*������Ϝ�'�<Z�N��kkC?�U���%nh����C{M�L[[��ֳ�T���6�Xާ�ᓖg����9�K����`tG
���F��=�c��ܜ3�X/�X�{���@Gcs���y?��ﯖ��Oʊ�
�u�U����+�.��J/kc�m��/&R&�	�x���|�p��z��$�2���/ >hx�M�k��`Ѯ�X���E ����=Z`�t:��"�t<�!��A0�YG��3��rGT5lŊ)(�p]Y�hf�#p>9���$��m�Z��'���|Bܝ��ؽ�/q��$KI:���U'Og`l���$�%�'�/_d�cp�qMƝ�I���;��VLD��Ɣ�V�K�J���T���J����>q�o? 8#;v@���̠�#�F��r�f�Z�l/[u�"�I�vg����[П
I����YT��!]7���,��A}s�Ǥ�-92e��H��H�f��I�Y�Q$�� W^�u���7�ei��B��Ti���գ�]l*��%~��c~���K=����\���$���ֳ�Ud���d�7���[����`��3Ot{��D3}����œ_5�3���L.��Ϯ���	�V�����Xq�A�HWz�>3X*W"7��H�'���9z,"���U��v�I4ڔ�EB��X��
'r���L���d���տJ@��q��5�ȕ�TJ����2I�S�-T/y�g�& �_�~f����U�[F�P#_	Lq�8�nR|��9��Jʥu��t�1�q1k.$,.�>��o̺\J�W�OS��Ů>��G3O�)�����#F	1搤A�굊Up.RJb����Cv�O�U�dl��{$oA�$��7J&�����-�1�����Z������?Fc��6'-��[�����G�?��Ԅ���Ʊ:����N� �1�DI�dz��<��a��з�a��(Dѿ{o-��S��M(52&n����.Qb'�F���-�t�,X(vD:�f�����Ӷ-�_�����.�ܜ��IU+K{��u���ݣd%[ɚ��Fֱ�!���Ih�1;�$'D�DA�*�(�yv�,~�����3�C� ~���)f!")b�/M�[O?��/�n�7�C��?�`9{��u%vfT7
U6�����5���j�hh@������E�I��-�3�ʒ�O���gO[��R��ix%ߑ�3�I�`�����{ىX8yJN��_v�	�����['����;��Y�,��Bc~��1+�Of$.7�$��7���#�x#����m��t����|�`�]�j�'�&����J�eS'���0C�c-�S��0�h�k;�T=3����^@I�C���s+G/�������
��?Yl�]�wV���z�7������3vG��z�Wf�>�Q�ؕ�"�6����w۾�Q_�����?����38����n!V�L�����&�<<��pWRYֿQ��	?���Sa6��_z_4ˋK��V��S�a������4�t����s�55�e������j��O�(:Pی8<�.�.�ac��& c�j@�~ߦR,<�E�{1��4l�
�Z�O����O$�#?^e�Vs�sj��W]��c��c9�R4�je��V��⅃ܨ���j�T�(l��Z��
\ͶS�#^ueB����M��g�D�E�w�7�����X���p*�
V"|��_��~�C-�<b�/7Y�k���%����r�i���*��Ӽ��.,�����wk�N��}�I{7�g�wR�6��~�I�>-�j���+���,ǃ�<;P��sl�nЕ�V@��:&j��&��y|��zo9�"֌���qq��L����8�y��h�7��2��%��7u��|苮����ѵ�m�&v8�'x��$�p"�+��$r�gXf��0?��G�3�����s(a~vE�e
U��B}�JE��{$c�?��㍔�m����p����{�������d4[Jp���#{�-y�Q4�oS���q�za�Ar�+��Bͯ��շ�zY� �ԓ���x����T���!o�HG!7n����4�DW�ܐ�E�E ��7?0_�:����R���� r=�@I�!y���2`'O����DQ�����^���EdTSh�Gl5��s��չ,�
O�R���[��f.=>��S��N<�u(��2�n枢� Wޟ(��&�@&�����P��$����;�����v��q��%5����*?I!+X���;���o�k�"�#�BM�W}��4�|m���-9j4|���K�ǃF��[U�R��+L٩�&Ei��x��x1K}Q��:�ɘl%A<���]+�,8:T���?�iq~�o
�P�5�z�Uo]B��oZ���A����
�3�,�W��X�Z�" Ƴ��A%��F���Bc|p]����mb��Kq���̂]���a�3��`�x]��~�K G�U�9 &�A�Q3:�)9�� �N&�`~�R}c��J��h��x!W4�Oh�o$0�s�嚋'�M�R&*� u¥S*��w���'��F�RI��<�t�����L�X~q��|�溵�zĽ/��|�x�j�mhd5׺����=��z�*/�������b_躒�*'�8��{x�芗���mc$ǉ�\�=*��G '������j��{h��%��l�˹�L��J�Gom�U�E:��֒=�V�=yJ^��*�2S��s�aO�ꡳ�@�y��g[��=���\*�!����	J~)��g��9`��uj��{����y�����e�tM�)��ĵ���Q�s_ �"~n�T���d	�'h��>O�#��V xR�4/�Pzm��1l�A����y&F���\���j#�V��s�����E�!�Ԙo��'�@��ԂCC6���;����Eo���ׯB�:]��[��(&�Kn�{�o���b3y��{1�{
Y�o���|�b7���O�T]�uE��k󄃱h����_�ũ�Pv�id+�f2�S��GH��T����FaQ����.��4w&H_��{����A]�T
Oz��OG_h���MվY����z�D/���������&W�r��W����n������q�_co~���)�Q�'E<�F�V὜��.��{g���W�cg�ၳ�%s)B�هS�V>�Q����s��XQ������P��G���@ۣ���U�r�J�sT�9��|E������^X"{��G����	~���")>�Uĝ�J�y��k��-�$�Ba%0fe�8r�/�ީ�UbĂz�����w�v�2ɵ���kE��=�)��t�����s-�zխ�c�� �v$��!x�0?�x�7� w��e�#�AJڛ���A�T���-Oc�N��G�GR���)�����=�fe�����5��|��mPd�V��M�L>*��Mz����Q�ԛr(��vh�?Yuq]8<౑�?k�ȨaBO�>N�(�D˹��K>t�^����5����S�0��T���00��B�$~C�����r$�R{[_�_ƚK�"��p4tv�F�&:�@`�i��D)>�q5p���Y��P��=��DJ��kP����
��}mV�� J���u3��i|�u,�<^��'COi4���$~��.M[�C���G���x����38<~�YR��������"�.��ف=t�i�?B c,HҶ�oJ���$�5���+|��6}�}�"�����h�H!7�G��;3���m$T�{�3݇�P9JCN���h��\T���Qj����h��@pw!4Ԇ�m<�v�n�v�3X�{s*�f�1	$1�b���Z��9`f����j,O*��N�[a���e1�����)K�U��դ80G�+�I�|���^ब��l����j*�no g�K��` �h��Q?��֜��Qpk���9����x�2����
�q_�8`���mOJ�3��=7��!	��e��L��$ʇ>�[� ��`�l�k#�I�5��|����Wx��L5��aB��e-D>)��bum��&^nR��������$7�s�!��$ǫE�៶�����{�9�(�����8{�@�`��^��Y�o�����ܿ��@Rb!0��cm464o4#�v��nAFl<��ۚ���V�8 z*���O(
m��F�ę��(�2���hաJ5�,��4��:��]���C��LŊ��7�LzE 
/�����K��GX�g_z#G��Я��`ܰ�Wy���<Wa�q�,��S�1�\�� ��� ������<�iJ�&/ӕ6 =�3�.��1���f�Y�|M�
�0
����1��j����!2�F��S	��/YD�M�,�R鑕�[GU�	 2 ����A�w:%7a_f_�5�뽎[c���ˇ�"=;�&W|hKH�+�Kɲ㤙��_��0�
ށT�	[��^�QE� ��GL?��R����)�T�Y���To�=0�ϞvV��{� 膄9ɡ�⩩�BI|]o-�R�V���D]�6��4�<'��ں�q�F*8m�]������_�xz�`m�{栒b�I�j�M;�15�޳�d\�?,?��h��{O�>�\�)�ά��0co=������:�c�`��0}�"�Q4t���"�_� �RF�Ϫ#���3�����e!dE ��.�ڽ%��h9�`T�dp�W����S�B�|K�^%K����?PN.G�����J|Q?����OZ��8d �P�� �1�k^S"�5�;�6J���3�(8��~ɝ�������yhQ�x���Re��7�ZGBy9���D׫�Qþ�-��ʓ@�3��%�ܿ�Cs/�G�p�|�%e����/w7<#��$:�%.�7=9gO]���m!ʙ��f�9s0������6���ެ�M�<�hÊ�}6m�V�&Q����lUT/*����������)���S���� �����Thf�N��0�c�3���M��:��4��,������YUyH��c�[G�O��:,EZ�6M)���2�]�S흏'B�l]l� 	n�.���y��޹j�@N��G�T:�ũ�邚�v�1j ty?�L�"�fqK,�:���\�A�7_��9{7�����5n�Q���7�̳�T� NE��pq�E��p�?�)�[+BC>�К�n�)�� &�]޲C9��y�k�Ȉz~�@)>�U=��VY��t"��0�`��*�����0;&�J�P(��T��U+�y���% 93�q��K�>������%��)�I�`��.�)�\
���	@�;4ܪ(��Pɋ�a�ʔ�3&J�����3�NGE�j�z��N�q����gxk�R�F-u�U��	d�KA���m�oY��b��^+�2>
��r+��������n�s���DI�%����F�C��r�#ڏ�!��9�A�Q�A{���ꌽ*V���q�&Qz��	���	��(�7��)ɉ�ʪ���Y��7��{�.$e"T�ߪ��zU��G��.��0��tuK��F=���p!$)��D���E�^p!�ު :�G�J�3��D�q�(��g�W|���=f�>���΢E�`�Es����D��F��~�r����׆�� �?��u��8'Oa���
:��MT���[]�b��-��U��[��֡`;�FoK.sYV].u�je��W!���:_�pg �)�sw:�ٗ���9j��=�����Бn�C�T�k	�v�{G�:-�/[w�"��vw9t*��	8��颰a���8�*dT�b���h�w>��x�3�LR>�$��P���xj��hƐ&zD��E����ئ[/������LB�N܆>W��Q�#�p{U׮�������� n��۸R�р(��m̻�W�k�N�l��n��o�-n�M2h�󌽱�ЯK��"��y�FKy.�`�o���%���+J��vRl��>���L��)Γ�"M
�F�P�!���3~t�����׉����F�7y�}���5x1{��C����c+I4�\j���u��s޲�~�3�nS��������bŲ��(f��~��y ۴�O��EH�BF"���Y���Ԉ�'Ld?�K��DccՆ�u6�IP�=����BK������ܙ0�u��a��.I^6"�槖� \u�s�f���v ^��6Y�����x�CZu�B�lBQB�a�, F'�%�ɟ�?sb���Ń�yZ�H�J�*&���}$ ��ƒ�V��ܒ�Ϳ剎1o�>�����f�<��z�:��$\�o�>3���PP�j^@�M0-g��r#E���_#?��B޷-v��n�EAh-H8!��^,U�J�<W���k+ΐq��E���W��U��i�1y��i�X��Ds,{��C���[��a��a���X^�~bXe���B ��}D�h�fa{��#��m-��2�7�'��1��R�3�#��ʼ4��Q	Ou��'�6p!-o_ucI$L����[���Y_�{E������Kc^uG5��($���@��n���lG홂�ak���Z�f�b�;@��"~��ɣ���ҭ����Ab��Œw��{��@���;u}�<��B�Dz��PL��� G���q��W��Hq$Ioφʺ�p	΋]�ݨx-�;�v&yI��j�|�-�.2
�E�"ۄ;��`&�N���2 ��D�_j�a��X��0(�Eu&吅w�$h�iO��ʟ\�_���\M�I�-i>�R��I�Ŋ�ַ� �tp���t[�����
3�`�
�+��k�����L��s,�<ĩ8[a��'"'\�h:a/�:_�����U�pFH�>o#jDc����$i�]��+�Q�K�W�%�>So��"�PX7���ɰ�mP�o�A���x1�"��c�E�cp�̑��j�ѥ�:|�s�l$�FF#����~ bķz(�\^������a�.�a� ��q�_�e���D&�� ��r����u��(�-����@�G`B���\C�8�6��.�7��S�����9�т{�	�J�qbl��F{|vx2�*z��4 K�b�kg�I	����l��r�RP���=�W�	�,��ט/d�U�o|�U���1x�9�Z�Ν6�f�64������z��Y���ʔ� ����S~��z�d��i�0r�'��3���	��Z+�:����"�%�=��`�V��v�4���Ԩ)���j�ݸ�~f��ہ�q럘-e�%a�Y�v!���!�<ȰǪ>ȦP:��
~~�5ў{M� �6j�Q�z��pT)-���|�e�����e�>�� ��a^ƌL@�ĭ����;���n�
H2&�=��N�v��]M�=�+'�q��{��W��I�틍	C��,.��]�JD��C�%%��Dj��7���˓	{'��?Ge�,�v��d�R�ۣ���s"ET�X�^3�O�-���>oqg*V��V�)�I2��[�ߒt��ˉ��|��p,=p�ϜꦘJyq��ߛ����շ׽9�Vv�i�F���@<�`H�	���7�p�1�uF��y�lZ���	�����>�T<�5i(7V-�e�����t�%s̭�^[����/�uaOP��B�h�1���Oᨿ�A���
e�(��ѡD���̓Fi�`�v���I�"t��<4�{�p�UufR�#���h8�\��k_��h���U!��tKd2����Ȱ��n������j$�E��CL���2z��87����^�\�1Ԁg���
�ę>*����K���/+�6r��ϙ0W`�0��s��к��@!��kK��D9�_�3r� �6"����Ŵ�K�Յ�x�N_5���a}^�X����#?G���Y�O�[Uh��Ҽ���:�BW�Y��cވrY*�\��&�
�NxBg�?�H���"��a�7 �c�f���r��Y�e�>����މZ�D��o1C;E��؟�t�"aYc@�Hϊ�M�L��^�
���e�F����.Ka�����]��	����ƌ;i��G��A��}��0���m}]�J|3��r��B��c+,���9�\�;0u���~��;3ʋ��������'F�Wg���m�`ʍ��RZ5���3�W��Ғw7�sl{�y�1K��F�Y�8�{Й�f��^�0�L�4��w�'h��_��41O �>Fi:�ͣ�ZXC�wij�#�1_�"�ř4~�B(�-�n��i��v����t�h�(~����~}E=���K��$�H�I���쵪v	�ז��������m�<�OC�����ʃ}9|��D	 c�*sAWx���9t��n�~i�j}����l�[���lQ��q}�F�����oZ�9Θ@di� �L�!je�`�G;�rVj?z���B�%Gwxu�քX��������r��W�]�h�$�	��a��7���VkS;�R�.��ġ��>J���1��6'�*#g�S��^{��"xu�r�
Kd���2�m�Ф����ҙ�N@H�,�h�s2��O���.:> p���@��dC���(=�Ҿ�#� �Mg����f�i6s| S�ئ��[�r. �[��S�3�v�y�wk�����
��Pe�Nf�Ӊ�a��qv�_�[�o�����c�����s��l�ZV����vX�0H1'|��a�۩������a�$�N?��Fq1��%�"j/NtSt �Aתּq&�m�Q���-%�U�o=��A�B���ۅx��*�x�Me��h,�]e�*��x3Z�Z��u�����Q�S��}h�rn�@p�ء��S�+��>�6C�#�.�W�'�tJ�	��-��#,�x����T���#��Q-��F%g�Ġ�_�x�������?
x�o-"�U��Ƚ�*'�]��4���|UYg�H��ӯ���!��ܼ����6���GW=��{��.�O�.�R��&�f��)KTs���E)�鹭��"Uu|7��2U�2R���Ÿ�L�����
���أ 9�Y�y��
pw�P�vE����@�I�1�����3���1��|zS��_Q�������+�0UG����:���۫2q�˽���-��H�#"��p�+�L�A|�&���{OCC��>*A'��ԔM`w��7R4^0|�+	Їպ�j'�晵�V�[z������F*z'_e��4ca����a�� IY�[i|C2��߅���!�_��X4<�2��X�З���I�-�#$Z�����@j�W(��� y�,�DG��A��0#1��Nr�-&��h�͕늩VvkeI��n��״���&�[O,c+�1���¤��?��ݶ���F���V�F,v_!�x��kXp�U��V���aV5�À^x<@�L��ݱ��%]����i%%=���Ov�xB���$�����F��\0����}���r����	�3n���y��6(j���~�T7�kNΧ�$�O9��3�T���6���!"�f�^�dr'ʰ�� +��(8��J��m��� ��괅��\T�V8}:�U�}t�$mb�n·�FI�;���Ku���L�k���ɼ*1� �l"67-|��m� 7��*��X��h�A]5�"��D�{��{��zꇗ2e��J3Ϟ#����Z�Th?N^�����j�`��nõ�J}���Z@ex
�w�*H���(����1���a��s ���i�9-m��Hk ��������W,�Z��C��}�������%�~��n�8���-a f�*`nk�_�
����8/MyF�B
����a���%�v�ܗ����S�Au'�^v�*���ht�V�2��u�w��x^�<�x"�b�/W���u�K��#�o4��,�q��P��t����	8�5�uf�鋡s���ar��_�!7�^���a�tZ���0ژhQ@u$�`��V�:����[���5�b�uiko��拈#�a��^�ջ���!������IG7���U�����O��Z��F��Me��k��	ʍHw�1�WY0��hnA�}7K�W*�;C���K��H���r��yG���[9b�D����}M ri��F8�
������a���3	m9�T������z0:5�ꍽ��FNht�E�ށ�^�Ne]�|r�j��<Ʌt����=�+�C�*���$���3*崤뭈�R�@��&��섅���#�p�����}��U�a��˪p�,~<`^�˹��^���y�Ē`G���W�+~#*��O��_�dMQc��?�Xyq��ٚ pJ�$�z�ܣ��t_\~��d��^�0� m
<��U���ǔ�c}�|���&��&CJ%,�h2�$��|�3�ǭ�l*�p�.9Mܷ߇z��N��HN/T���U�Υ0��P
\G�ËE�eӎ���Ɂ)���u�L�b�½�o[�Ϥ�MN��ބ�{��z.�>7�P�����1���&���t=P9�n�ޥr�n��Z#��z)�$I���A�7?��(��a���ڢ>�Q�>Ɩ�h��O�D���ȴL�N���>J�X�9��?r�Ii���kk+XO}���$��$���pq8k�� �����V��unj��s��Tj�7�pѸ����JY�R]�T:3/��ΌYJ��Uț�-�#�v�ixDg��oZae9��d3B#éVĘI���{�g`4�)�r�H��P�	"��4 �����|�⎠�\�>~��8��r��l�2������k[����Z�v���+�G��R6N�ʚ�*���v��ң_sՙڎ��ai�Q$�P�[4��!���.�%�h�z�-W�5�`z�������ЛZ���.�ֳ�X�ҝws��Ĉ�(� �м�+��+��d���E	t�/u��`���=Q4��k�:�����f���D4��6�sc��Z��)7�_z6Qe	��j�B8}�dud�������鶴G�a�k���!y�`lV����2%��آ�z�9�Bn�8X H�Q��g�㢨��?�� 9��%�
��Ag��ز�U5X�v�X�%���H�7��C[��:K��?"�ۛ��"��`�{�H�7�Wr1���h#B�M��5%ͼY���\$�k;[��JZ}X � �L-U}:�hO�˵St��8�{����y�$Q�)h��w�f�$�KE��xߊ���&��.��N��,�E���Ҋ^�a�'��Vl����#'�Y��3	�o	�\�n���Df��y
����� �6"�z`�6=��~��
?��O5qU��������4�KE�ͧM�d0d�g#X����l��k;��O�t >s�z8�Q���Zu�����y��S��ȸ�����=�P)����{u-���=�����CR|��f�<�0.�M#|"/^ ��@k�q�W|n�-y2��A��Y[���:C�kM7S�>���T�c,�J-�::�fe[�HS����~NB�+�9�x}�>�g��k΍�������ƾn,�lw�0+��kL��'�.��q����ב�F���N����^�\x1iF�)ҋd�4���ô��UT����E��>0|�308��향�+�;GL�&&uf�2����-e
��6s!��fԩ�&��ʘ��z/7LNֺa�W/��\��*�pQ�+�35�1�������5H[��Ai~�kBX�^�Ře������h�7��ℍFY>��`����Q$j��7Ƴ[��+n�zg�BO�����nR��j�6 #r~1?>C`�J� ?Lڇ����6�@e�/X'�)o��IC00��湪�G�wd�͊����#���ǉ�K{�3������@ޓk�0�n������tmk�S,��e�O��~AxN�W����1��8Dr���1��Y����__Kӝ��D	3�͌F�Z��[r���st�B�A���F�l����گd%�J��r ��=��!��v�����Hn�Y�}YD-#[���t����-ԁ��>��р�]S4����r�>x��n,Ο�����z�Q���A�	��#�BX��1��Z�/4f�L,)�|������3O�Ȟ�Q�o��g�Li[%$�c`EM\��M��1��Mqָ��i���t:i���N�y�i�[5
m��+���s������03�͵�?�J��΃�7����ei�Ub�j-��Ic� (�m
}Z�$�Х�Ri_�=�~3"��%�-יbזA���f�7'�)7�-b{2,!����V�8�B���o}�@rcy���i8���5��j���sb�Aq˚���+�MPn��7'��u��L��%�m~���1#Ru�f���t�������^u��C�v�-?t�.�!�wzB��-
��#�ʜ4�83�J�PZB�����ߝwޘJ����I�CX�N�'CWq/��#BӒR�E�$�7{9�M��=�:�g�L�
H+��E�4$@ ������W��t3��6�z\m
��4�L�4fz���E����}�RE�aI�R���ݰL�Pd<�F�'b�/r^���a���JT�������
�t��y�U�~���ظ!��K��ojL;��~��ފ��rMp�˹J���i���7k��v�-�HU��n�`�[���und/���䔴g��ad_e�Zg���p�N|����v?���q�������zp��?e`�]u�9�Sjf�>�K�p�����R�P�2|ogPʿ���O���`��,�t�pV<U�����%��<8���)�=��,��P��;�T�y�����ͣ9�+(����i�3��5K�*�Ԩ��?��Wj�>2��V��������Kb)d�az��t�{����5�'�g�UP��Y|]�1�x���@�MҪ4�Y�V�T3Ⱥ��l�dMd��[�s16p�u~�\~��
~�b}P�G(7�L��r.b�*�;�7e����&�V����y�FB��
���ы�N�#G�%y[*hz�ǯ�nR|P��g�r�x��ߛW޼�[�J�sm�א������HW�����s�A��]��jur�g)�˷�O(A/.
�̝��������l�w�@�_��w�D����:^7B;&+VB�j__�%*���4�Tp��l��5��?�v���+p�.�+R33V$��^�}��1 m\��`��ˎlJW�֡�r:ۃ���]5=���,Vo�QWo�g�����DQ?r2�x[�J6z�2`cL(��,����g�|2xA����h�-�!�y��	�-��{���%��Y���E��Oi⫠p.��_X�	b�*�֬f�H�Wp�Axp�1@��ؿ-�4�Z8�z��|��ޝ�S�g/:N�<?�LRǃP�Q>�y�]�ڞ(�`��&5��U	j�q7F@�xݿ-	,Ɋ��S�Rf��������S�Pzf�
���N7�2�� �躚��=�A�=�0l�ߊ�a�G��h�!�xm(ͥ�ښ�V���`^J�1�#���zd�^���X�A e���GZ��R@�&׍��k��Lbx��\G�_�G�6D6$�PRa�	�>�1^!t�<摠X<��<E=s��{�E���Ó}����M�,���`�Q�Me%����Z�ex���|�7�6�̛��%�-a ����p��x�Jh0Z3N��>�e9P���po�X���a`祡f����j
)����q"�pԻ�*�N]5z8e2�)t�����;9���fMl��io��L1u�UFF��*B��;�en�mW��d�Xԝ���� �6��Mg2�����%����X��D���\a	�Ā*���S�À��5�26�r��?=|WBi�,�/��L��Ē� *XJ'1��$F�R$ȳd(�����*}�y4?� Ni�3��uVpl���'d��D����BU�4��@���j�Nd(T:hvhJ��.�z�#����[�zF�-\��u͋2uD�ݔ`x>��<}��&͇�HM�A+��lEq������K�W�&�����`}���19�ϻ�@�	�b0R٬�b��n�8A<�^�2f����J:��{��WӬ܀�Yu���>�&���Y��> s�B�i9��Q�բ�_ �� hzm�g�#��e��%���pi^�e�bP�5���MN>
<_��>.�����/�f{���Ca�� ��.�ʱ��5��B�..	��.�G�Y��x[���C�s}B��C������&����E����'�q ���=(�k�A?Ƞ�Ƃ�uʅBR���9��[�V��؏j��=3�/(�E4/.oR���(��)(��u0K@M�U��#}���5��!�L��x��M��
LV_9iz���;�%�|�֐Yo��w�HU�r\��@CU�48|13�4#�C�a<��%L��Dh�d�`�ч�3�}q�r�=�kR����IɉL�8M�L׮~�76��::����tc�.�	��	��9t�Oo�;�c"�ת�[�=�M����K;U'��XP�A|�j_*V�%L�A)=X j},<�1+3����(�8�9���Ў9�1�Tc�� ��) DN��V�/r��}腈������ޣC�+�����r���1��w�H�)V����#R�v�Lˏ��y6+K�����LJ�t�o�q��l��7m+���\7��*m��Cc��w�t�� ��+��Sw���8v��.�%/�{��i�;�K�¾��_�����wi�b�@`�)(���[ķ��t�xr�ł}y��B'|&F�ӕ�W��v��H�~�W���͂8����N��2��c��Fz���F�>1OPui����ϖ�	 H��gb�)s0/)l�~�ҼA��b�;������ (/�Gp%S�MF ��%��9;�0}�'"��Tm��H�����8-�����LtQ��ɿ�R=���ujك�`=sCB5����v_-����Im��M}���^M������'�5C�ݍ�g�nb9q�O�,��{-o׎g�P|m�,T ~��H쟭��+�.�X��`�B�7�a��
A�Q����U�4u���͠cG�d����G���@�2W8Gc��cS$ֆ!q��HJئ�&oR<㣗��e�x[O��R���$��
�"(��w� ��N
ܥ�VMN7�z�y��2˞3,�A����*)e�-�՚s���$�[v�S�grjz��Fa5�6/Ϻ����*����j�ON�����̉�^�+Ƈ����h�|���%z}"�U�9�N$�`�'�l.�9�I���>�\= ������L��/�RV�@�ʾ����V��6�[���1�ЉYhJ�#�(W��p�
U�k��3)��K#N:�K�̺PH�����VE�GSH~*�X��#����W��s�Gn�hM�]jS8�?�B�Ki%_��J9�5DJѾ������޼Dg�n#�{m�յ�!y��������~X���3�o5w
X�6�0����l���"*�k��ͺ�{�W4�h��p�ք{"T=�\.2���É�d8����׵Ľ�4�*bS�V��3)*�r�(��l�tzly;}^�FFý�<������RU�I��?P�r����M\�dd[�����g[�nk嚼$(��e��W�w�zI]m��uzd�C^i�:��F���(��X2\��
�p��8:��B��
���kA���g����&~S�5�o��9���4W�*�YKC�h[��-�b-0`1��ٙ�ڵ��/�VS-���Ƀ����J�x�1|b���WF��g!�^)���n�D8������Z�k�D��C�C�)��$���)4a�K���>tB���l^X�6K�,����ѹ#��v���6���?�۳�`x�Cu�ĳ�na�Z�d��pZ�v�N+ Q�3�&Ra=�R�D�vQ^7Uv��~���P�c��e��:��-�@��/�غe�Kƚr�).=��T<�+���]�t<��"�7nr�`(=
���3�4�)	�MJ>ɲ��
�llw�rS�M���I���AWZa�tK�X�6�Y�	�P*#������D�w*���PЃ`�Yzhx�/�
$�ߏ����0�cU��sBlǊ��ñ�-��U�e����M�c l_}�<C�no���w�? @�SRm�K\>j����"j�T����3^R���W��*�����"�O���V�˘�������}Ԕ8�J���ڡ����(+���/�b'g�AU3 g�`��E�`�?p>�S����7[�Ƨ���ixص�`d�aǥ�zC����+��q,?,��&��ڋ�v(�����c���t%�ĩ`e:J=�F���ol'�!�ߎ�"9h������6��Y~X�U�)��`e�_�:_���k�?q��u�|����c_�dZ���\�*>|�O�j�;�x�Y�.�J��V|��i�]�������p��i�����5�����)߂��;��r
W���3�+	�������>�Ct���W9��q�_�dA|� �!J��� 1]�q񥖟��<H[��7�͝c�J���8|�/���c���T)R92��'|��4�P���z6_ق���ePM���v�<-���k�Ql����w�Ն��i���c��x�TG�F�D�-�1YҼH; �A�a�sM���*���N���v�v�\"��3`�����[t��Z��%vgv���!;KW���w��Z�̓�����fٱV-V7v���j�7>*����ɩ�a�2�F[��=��r�>l�N�]�|&w�O�[�L��؏���a�mƾQ3�UUr�̭5�]7
�
������)�������dk	f����7U�T;��Q-쭍��-e�ݹ����i��Q��
a��$�'��
F#��6Yo�pY�6�χs����#\oǙ������q���C�ᴟ�5m��/��<�d�s�هG:��j�2��;#�v���Kn�9�G'��Uկ��^]J�'�������o/�>�$�[��m��kZ�kq�{��<+rJ2m���A�n�=ӓ\]�U�C΀ ��]���6�u���3D�����;��h\_��B��*�$�@����n����+K.B�M���һ��#}������}��K�+#���v��84��u[i-/T[�XB�k\�&j�>!�!kRI��W��m��ge�Q�Y~��t�����_�~u�ۗB?.���K	-��i����M���q��f��u`?�_Ī1JaS��`�D��Ű۟1���܌��a��y�*���3+��{�OP��cuLO>�z�����U����du��6����w��\���\^iN^�vr�ߊ��F�L�w�۪b���[Rr�_,4�J���4����UW6���=��|+�	� YPG�#�%0nR�ȭ�ӝa�L��H(��~ݗ֪GY���CqA�N�q�3�*��*������-����8z�����ͅ	Z�P��>�pv�M�a�MX*���ie��Y	X#��&*+��� �H-\~�%'���1���0 ��l�4 ��԰��T������y��"D �y�5�	�d<�ynJ~`[n����TzΈ��&����0�����g;��18r<]�t � Q�Fs�S�S�ʋ����#���h�hL�	�;�bw=��Є����C�� v\�K���J�+��_��'�*�^�(��j�A�c!�R���:��3�V?۳z`Ƙ� '�-���T>���6��_�GF�	�I?c6|�F��9M�(D<�'����j��G)_<���1�\N��8��9�������w�8��,�>��6u�\�S;���ܹ�x��k��3�<���U�y0 w��%�5C�T^������`Ć��c�����]�����nm{��L74��q=j��1էId�܅(�}X���`FzuW�����'V#� �n5>���:o��͢�+�w�P�o3�5�$�y�:��j����;)L"F:M¸��J�V�� �\Nk�{I��f��١���{H��k5������6�����$�- d��0̻ݤ@��xOɹ�H�)+g^����p�@�F�[�jT!��r�������2ǰ���h��>���ր�d/���x��ŰM��^��~DM�j�h���L�s�n�,��Y�� �6|���]l�{q�Ò+m��Օ1rV;���c�Sp��3��l�g)��������4� ��R�5���7�k'-�����#	Kv�22��eN�j;)51���H�FL��.N���V38�u)���&kIM���IsAh�o��@^�m�~Ѯ����_�ޭt[2���0+�eS�&�N���F�#�n��`��~iy�9�/8>�G	���|��3L�/%r~�B
qߧy���>�Tހf�̜%��]v[��؅�?�2���^���X������u����np!1���y]�{.�`��o�V(>�N$s�Z�p4k������� �!i	�A��Z��Z����$�t��w�)"x��H�����+��Q�F��\)�����"�0k���Λ��F�� ۆ�e�`���~�e��S^:ٸ�ɃC�h>6x���_ڒp�+�V͂y�G���^��^J�=u�f{}H��x�5t}I���Ά=5��*�{��������O�$�2���\��_љr�>�"m�
�$�����<`^ ��?���:�;�6���'�j]�Q>:z�~�%��\ Z ڼ,0���я�g��L.L�n#��`�m�s��2��K��8�j��~sb���^���V��"Hx��� ��ϴ�':Q��ID�S6�;��آޛ�?�]K����"����8r���� �c�J♐����^����4����G���(p�ֽ������>��	xq�5��yz����@�ȝh=����	lPs��.C�%�;6����:�{�%�`�����������T?���<%�%ч|U3�j��:�J�6�k@��fw��^(�D��b[UF�ꢼ�Ԇ(��F���Mރ
��3?-���
�?F�Z�|�{b�>�0!i�?�Yg����dn#���aR5��q�'O��I�����Q'� Ie兙v}b3b����u�ѩ�ЧZ�PQ�3"�*;!m�$�G��R��)�GF`����
�q%����f���h����{K����.��)�ZYDM�M���@!}C��>=�T�I���t�"�3��f�k�O5�r*�M���as�o@��E_qg�!X�(ц<�J�>J,���"h�%�>�c*���^���6��C��Û	N��n�u�X���Ř�霴5�%9��YL�^�ETÃ�HpY���2�&�.�k���Hz��r�Sh�{V�n�ǡCxf]V�|����B�H��fu�b^ApEk.�qxg<R��c��N銽n��vM�����v������!.�"n��􆞀�Ϝ8ΐPK�Sgfߴy�~��ޣ�Ppu�9���ۊq7~�t�둍�~���vD�M��O�]��U����Xp�֪�n�4fUum��aذ�p�v�!�^���;#0(G��if�7�@�� ` w��R ^��2T1��q+���v;|9_����[f�qy�r��3��ūa�W�Q��fel�b�inZ2����x�e9������FlO5Q�f��xd�^?H8IB�ӹ�$)�o8\��Ǳ�t�״d�p���i�wX�w����4�Ե+�����}��oPp���� �R�}�`�h�Ž�O�̥��4?�Ak0=����s>0Y�ɭAhq<M/}y�Z�)�G./����Y��Va|��ô}g�A�sw������Nmq�3�Yj��|�m��+�Kd���J,���b�C;��K�ɢ+/L��	���<k�ΗI��"/�$J	}�����m���e���������TAW����[�bО��d-��s��oʌ��40���~� � ��͎cFm>�ǁ�2���&Ź|�+��|fZU�Ĵ�@&�sø�QOÕg�m1�nr��o�La,ld�hZ����i�S�0�u�&j�h��!N#����FU$z!�\�̃�L�����7}�X�
�Z<�0`C���.����x��_C�Y�3�w�����F��I8k�[o�~��|_q.j�_h��Eؔ���d���}c��%��$�oTw A+�j�W�Y8������"���[|Md79pH��f��I�(���BP�Xw�����ia0�������܅Y	����\z>�._̚Vgl9I�.���k�-O��jc���UQ���YTå�yo��Sk%�!�b!��1���\)J��{�H���c�� ��&Q҉��5;R���`A$Z4�3w�J���[�*E���'��mu��Y�	��Nɸ�V�=���y�ߕ�D/��1"Q��@2k����tV�e�u}�N�nnz/TK DG,rNL�t��Q��o�{q�Y��~�a%�v4�b �:��Dx%��{> 4Ġ�&�[���8qo"��j�(�0m�(-��nY?�[�v���y$�z�M�����2���N/Be�k�svr��	����}|ao
�C��]��f�D�'p�~c�g@��=KW��[z�e&��AH���bh|qel;�=�Z�R�`DŚ��_n��=Ƅ�j�Na�hle`����)��{�;Ò����C���j��|�rW�'$�s"rȉ����kgu`A��x?6d����9@�}z��P�F�3�|as��5ƹ a�6�+k[�v��@��u~[��eT�]o�qP��a�#���gӍ����z����x��3X;0C��ED���v�k�"����g1=`[Y(�-2��jr�sϨ�MȄ*߃�36Z�G�ym�Z,e�,��6R��ܧ7ZKzȲ��N;�$Lw8�c�4~��a��:nٞ��d	���Ѡ�0��~�6�2����)�{&�i�\��F���;��O92!mjkE�fn+��i���쓡 �<uKjG8��tMT��R-  ��k��ӵ$mFUc�_�3(������˥�Vqʵ��=gQ��v����4�^��/mP�@1J���d*���R�ʩ�d�lv[�M>�{���{f�7�����9�׭p����%8���ڔ,>Ĕ��k���N�z]�ʩ(�	�y8�9�Չ��T	R�������鮥��/���Wu�6.��e�r'�0�-� � q'Z(�G�	�{�	2���y�.�$�o���I7H��m�%<��,�I8�K�u��6�~��l	��@�]�͘}(�J_�����D�jT�TZ�p� �?{�M%^t>?�FJ����U�;MG���kϔ��<#T!i��c^Au<>2�,���/:̵H�����iW"'7yF����7�s����5��\��D���vA��e�P��|�Zj�h�t�������,�5���mmԓ����c��1�܀۞�2�0�@��AQ������T�����>!�t/O��r�;�P���w��n0ӷ��z�l�?��i��9d�5d� ��*�&���­���5H��[�2-*�b�mÖ�X��Cũ�_�4��@�%����.�> L�S �k0˒��\�D�-���J�\$��W�����+C�+��l�D-��4TW��$�NY��_%�JUmt��	us���7	Դ��_�E������	�ܖa��Jf%��?o�6/���H�>�7�;�Bu��!:�9� ��_:8���>ja��P<���S�������t�W/�O}�	��t�G��~e0��u���`�d�P�X��:(��t����Y]L3���2�Qr�s��_��+��ܛ	�O V���kI�bq&���FQ��i❉����&�y�i���;��zPh2�Ts�	��'~ڋ&:y����o���*z�d���c���%���ã͠-f:?��u[Y�k�S��<��>C���dr��?�� >�X�d���Hf��G�̮Ĥ�j�'|�|�Ԧ{/��0�Kє���]���:���Z��B����#M�[��9A�����mN��=`��2�~F�0o���>�O�Lq/Dc+5��c ���5�Cྏ	y!k�(--� ��X���]R�{~w��D/� ]"�A�j�➒�P=�tk7�������G�ė'qn\����6�.�=>�J-�Nzk6�A�x�ߢ�	��U�ld�yi�q5�����[�A	C�Rƞ��sn�\w�7�}  ��,c��`����G�L�p������,��mDZ%�,!��9�t���x�"��x�%���J��Fħ�>�Vv�N�����=���P7�F_�o1�]�H�����F�yҜ�� �Y��G��w����F�Ib!�w]HȑS�+�?����0y�k��-WG�֮1x�C��²��P�����>\�6
8�����ʩ�	��6I�311	���������CE�B���9f�,A�ԅ �gatO���2��Ve�$Y���<)M�>���e�%��d��O+����u�4���/� �t�ۻ�)����� ôQ���Dt]��H��� �<n�u	&>>���1�N7���N������C��Sf�Ñ���� y��O���6���KOJʑ��d�0ߧbD�xL/���u�-@?*�����C�@��+�!1�|�uT�{>srD���β�h.���IY�,l<oJ������O�5�s�~��^"��έA����`�f]���5GЖ�ȧ��ID�D\E9��WI{<d|n��1����}󏃓|K+���~�&�p�|���O2�&��Ћ�s�*����l}3|�����S�ViK�w�0�G���&},�|E:�gM'���.m~>�_`j�T���q���wݔڍ�+z�G�
&6�}z���)�ȿ�8x:X|!����s!��N�y�4d3�u�j� ��ְJ9����
?[��� �z{s�] =�2���[&'H��kA�q�Kݹ;�k�t��x5��'в���!�F��~ɴ���ʣ���)R���E�/��^�
.�౸}�v�Lg���bid*�JS^�}Aos\kn��/{ΏM��!��i���%����uCm룆vL=��Ӆy(�
��T�����9%�L�y���h��)�:�G�u�9+|<�� &�\Ҡ��?�gB2��(�6��b���M-�U_I�[W�Ph�`X_��b���WXg�����i_�-�xSXk�oF���<�����0�{P��c���vI���%����-1#���ÑfX�9Z���Љ��8����%�:�6��sRNz�u7�%�(�Pd�O3�M{��ئ��"3��Z7���h��*�;���s� �N��㴇�{[9u�%�k�E���"J���[`8����I)�X�l��
:m�l��z�AHo7HG����/�VX�5�b��!��C��J�L E꥓-�q�w�q���#@&�ް�v�kQ���W2�9���F�c|���/�{�L�M�iy&1�[		I�{�|#�_[�i�4g�
��Y)������ �U,����P�U����[�7U|�����X7���� Ǒ�SZ5��\�HD��������[^ z���<��՜�$�d�_��(�
y�h�o"�D�3z2ɑ�n�}�g��i�H�+ �`�����_�?&-ś/w�'��,�cl���H����궩�JE��-NV,T��/���S|њGǢ̵��"s�1�&�w��V�=��݃#�SBm�
�!BxJ���C:5qf�~�y���g�BZ�Cti�� �#^_�P�!�Ti�t��N�����3�GJ0f��:��UQ��9����L��'P� ^4�A���RJL����a�]D�dM'fu��E8��ۀ�����O��e��O��
yz�7�3��`1.�S�$�pҴ>ƈ֋�����`.{e���V	�׫�sw��>�O����$a_c�}��Ţ&c����E�6,O`�>G�į'�3Aa��]�i�Ƒe���	y�G�pB�+�+�!�-�o�*�sF;���v�'@kf����z�_��G�6����i���ф��~O��l�eI��ZϠ �"�C\j�%#�d�]d�W 5�;�P�9ʶI�(jS��[��L�����b��§�9�J�έ!�"���t�x�G<����1���s��|ZL]>hn3.1c)�<��1�BLPe��� �_e������G ���4Ԁ@�j҄��ж�yCG�}�/$����0�����eR��X��jztߔ����D�JO=y�	�	�?΋A�����+�H���9R_�����}Q�@���T�C~��0^wfjrGHF6�6F�
p���� �'�fvG��ㆥ=S2%��L?4�K�<��\�;y}5���ʭ�e�_��R��i{0�g�O��p��}�s�s�vxb��Q3�ȲA.25°)��ō��CÑ�cy&.��D�_�n�?,I�H��C���w܊a)8��N�6��7�`	��D��ق00�I�@�|��1[�#���d�M����\D��g	[ Q1ȃ<�l�+N�,��U�ht�B���6+�#���+��/��_���R����Br���Aݗ�[�.���⅁�ō�w�*�����u�YIe�Kh��m�)kn��ޯ(K<.Z8#$�E�m��L��܆e��M�˒�闞{�G��OG����S�
�m�w�Ke���n<�>�z|�ȅ��!�_���oЙe�l0��=�x��u��ϴ.O��n���+�<��b�	��w�(xq�=Kr���^�c��~*����e�q�n#Xo��3�⾟K���2qqr-���C�AV��.��p�˒S�(.����Pp�l)��#�e��}�N@��	��d6�noNO�����~֨�1A�|Y)�r�Jۂ�_k/�r0+��"}��0,5�0ڱw'<�zW��4�8�y�dcza��4fK%����HQ���ra����9�/6%�&�B^>(�	D�a�_A������ɻdu�]ё��=� �5����R2�H��ۿ�x����:$@�OS0�&��I?�T3gX�
��,�����%E��Hx����G7�P��oY�+�NjSϒ���+���Й��jle;����Aѥ��W�K`�呱u���W)���v��{J}���$��_���`3�=���`�W�ͥ���-��S�"�0`L�8�o?�&��{�Î�>6D�:^-�5o���ck�.ef���4%��n!��%g���(��B�������OA�j�t�:��<n�Yfz?��
Vp�9��Q��~��'�\>v����^�ڂ	��ҿֵ�t���8�`��kwRYKڐ�-�l���6DG�Y�_YJ�5��[c�f
�~�L�����1�8�7%��@h�����q���Ψ/�q�2F4�]��E���	� �[µ�ǳ[dJ*)��,ٍ���m�Q��D��6�kϲ|~j���T	m�r��3�p0��΢S�4�$�G8���b����N�	ȶ�^5�&b�{��Qj����}�q���}�»� 4k�U�sv#>���(��*��M��ε�Q�{�Ft�g��`l,*���%�a� i�z����Wp���M�#�*�o<��^�/ߕh�CT��-QW�&�N��.���a��8�6�|�����M~��t���7{�Q�Ձ���xE͐i�~�@a��'�U�{�,�L�����/iQk��C��a���,/�]%�ߎ��)�-�ｨKnR t.o�k�}�Ȍƪ�i�?17\S�f�W����|B�lSr�^�1S\b-��b�-��D��揋���银�����;Qlj���/t���_�)���i���7��%�)����߱W2�	�g`ru���ByT����p%:z�pxZ�kba���C���U�n��A��t��Z`�$��@17irmf��a�ד/���x��;Cl��э��w:b�e��Ʒx���Þ�Zx6ΐ̔�*D�=i�N㸪^;A����� �^a��2����jJ�Do'���+{��Qc�Sw�qQ��E5��> �b-H�Cj�Ӑw��M�d�4(��q]4���gʷ���=��oP{�@P�97ɱ�E�j�W��v>Ɵ8[q�K������aoc���[ل�`�ɦ��贘�V=�-v  �}ik)��T�>P�E^͆�h^������FZ�Uz�+�G�s�VHP�`8�WT�{6�O`��<0(VNUz�����5GɃQ��l���
.�����:�<����2��T�]!���2�c/Ob��.����_I������������q�'����ش߲�B�3�䓀�ez��^�R1�3�=dXo����dk�)��zJ�u"�=�]1��7��. ���'�yU�{�n·�S��^N��hH@��R�g �.'Am�Z�BWz�?�ו!�?�pSR5��-e-}��Xѣ�|�";����:"�Jka��0����gDz�V�d;`pǭ��-����a)�r�%�
[�T*��,(.�Ӻ�G�:�	��-ǩ0_�v�E'�������0D�)Zz�E��@�Y�N��_x�
�w�h�;%�m��?��}��P�*3k�rs吴e+U�
l�p��l�T���qI���/B���w`]y�����6��Y��2R��cV� �rˊ+���k�_���Ƕ���d�w�i��GHo��_��+bv�0FV~��(���O�G�^JhW�E@u�"���h̲ȓh�^�΄'��wV�<B�I��Q�@��C4�͕�qB졬p�و�@]�W���iZ�L��8��z��#�h���\�Q��S�s�8�)�Ht�\�3N_@T��UgA��pbb!��1�da�C����ҩvS�7	�!䵒� !�R �?�n��;r(�����`;p��P�=L��������n��?�J5��(���r3@���7!��t�f�f���2�F#��RR_��1���L4./(L��
�C���z)��Ϥ������D#(�<��@���ȼC%K~��� �k�o��H�j���yUbr���!z���8~/{�Ց������V�C<80t�.�5+�h������H݌�K���B��㹖�Y��PQ?
� ȷ���~�T1��R�	�n�WlB6n_}v�R� չ�,g�T*߫5��d�P#p]���wg;bQM6�������=u@�h���u;�?M1m��p�o��0�	y��O��%m��c��zUk�:���:�k�L=���o"Wӹ]/�xO�濭��u���q��6����F���G6�'����
��L��N�Ewv;k�5p5�:Ԭ�A��;-�à�C�0C`���W�(�\<���CR��出��ێ:-a&�V���䦙�`�s��,���KoZ��!3f�-{
f���c�6��pk������79�i�wM�j浺������J�a�lF�^�Uɷ�%\�\C��C$z�&�4��N���i2ч�J�XK\��st��2�p!����j�x�٫;���V�l)�h�H�}�T��)`1�M��f�I������� �j~64RG���R��")k^�R	z�suF\ر�.ڒ��f����'��=�P�%�6'�Y`��q,K�G=��ۄJ�]�Mk-ߏ�N�ޛ+6!3������D��ŕ,"��b���e�ٔ��|z��t�F��E�9�)�v9&>^�D�N�[�%���@=ۓ6#�e3͘)9�M�W��@G��=T��^�hR���	��S������y��)J|및b���&|I�a��ͦ��O��dO�
���U �1��v�t��b.�s�5	�߶�9�V�K��/݊��1�� ?�9�O�/�KJ�T���'�Z�پ9�$9��ĪMS�&5���0"N�[UOf����U$�s��ϙ2u��i�k���7k�T���������~#1
E�_K��g��� (�ʴ��D���΁��T��;�?����xu��4�¯��ǝe��$����{ք���4 t1�H�r奋��4�dP��}�E���~#��&�-1N�����9[�%�I���d8��L`�xI`����Cy2����&r#&��$�D{��\���������Y�T޺F�؈U9Eø��M���u ?S�g���>�����I���Ƌ��ڭ�����u����'Z.���j�kq��$I)юq����f��֌�q��M��-b��U�2Yi߸��C��T��y����uY�O����_=ɗ������+%�6����#bI�M���x{̎��H\)�*�d����c���/�����R���m�_H��f+ig#���e�Au_����Kih��Wf��#�����V"vW��g��t���$l��kn�(�5MB��y�T�s�ӗE����uH&91+�z�i��L���Sg�}�:|F�+�?� p�,����͠�Z�ﲄ��Xv(���:s=�i�����g��g
�~�����f�Z���L �<���n0r�<��Vԋ�D�T(X�q���=(�R[x�Wf��xsA0_���J݊�zL|U������:X+�"�����X���s���*�<��	�V��f���Vi���v�-{��mW#)�<6��%��4�$b���k�+z��i�g���\eX�Dj �T�z_=���=��	8�*���X;�0��;�:e ���}=�M��]�J)�gG�3�-������z�E*Ywn0cϱ�݋FG*���-�Ҿg&�Pc����Y"�ڵ!h���A���h�M�H�?��W��+tv���7L��`!�cQG����\��[�d�e���{%|�����B��_����ǣ��|NR�eYV#z]����Y ��Vl2��E~��8�dd͗|�	&��6@�$�૞�H�p�A���*��H����k+�X�B���7�f�w�ၚj��>YN�qz��UE�r��9_��j\c��Uz�ۂ�>C`�_��B�_���}ø'�k�/��(ݏ��4Ϣ°_n2H�� K<�����~����a��)F��^~�C@9tC����%���!�h������3�����Ԇ���҇��Ź2�kf�ܻ�:�D4�TQ"��c�g�j#�G�l��N{A�tn��Q��	�$��]�ظ�
����0�7���5[�y�Z�&�-�F&?�
��G�-�u�O_I��K\�W�`F��]���p$��� 9���q�C���VG<�Ba���T[�{fF�m��i��J*ͯ�u�=k�=p�����(|�PEL��<�x�jKK�X;ͅIǊ����t}ދ��ŧ�Ǿ5]���2dQ�i�t��i�xI�M.��0��0)N��Xe�@:�߆�Z��6E�Bs��ݐ�k�T�����,�i��5Mh�T�Y���w�d�+�+��+�g���\�vf+�"I�}�oS���U�.W��N�
͊]Q/��=�n���|ړ�N��V����ZV�P��Ǝ�:��OY��BWh�ڙIī�(1be�Yd;�#>�e2�b�a2����sKATc��鵟=����(@��Q���pW#S��{),����ك�Ax%��~ K�o��y<���y.(<d����0�^,�����\Dm���%�����c>�.Iy��{R�P�����jA������Ӯ�����3 -m�MM�Υ�RF��q�Ș7Hpvp>��}��u6���u�Х㏔�F}�_L]FhA \���]	���⢂iB�U������Q�r}�%�I]��39q�g��8�Gv�g�_�
?*�[�� )¢{uM5�	e���6�=]���Z6���n5���>�%"���C�����Jìv�I2�(���[Z	J�~ �*bِ���S7y��_M�in��K��C��X����2�R͢�	As�#�xk��M4W��Q���uFED���Ab��4�"ڿ�ٮK�X~.͇�5$����d����,�������>#*�fǺ�V1ln�\���(U��<�)�������"$&�vY� ������nn��F�e�A�x�3F>9�a�MdRk	��gX�L!��I]V�}����U	ǐ�0�b�~jS!S�.��I���z��W�X��ō�^d(��wm��S�����ʶQ��I���/��k����E%#�Un�6� �à��U-��V7L5���(/~K�>)��z:`���U{��m@���S'���8�rZ0)�n ����c`e�{�s9et_�&��j�O�P8@�\���,��5��x�-�ah�Ih�b\]Ef�O�ș�vЄ�rZ�pWU�O5�����5��,}.a}�ن�<�إ�R�P��~���W
��E�׶K���&�����b��?UĸE�h��%�AP	$Y���<�t��O��:�Ҥ� �#��V8��Ӄ���W��(�W�J�sE'g��Q����B��6vvRMbZkR���p�Nw�#&J�P��'A5�"m&��� ]ɓ�jH�RW�h����l?Kwpq3���Ȃ�����[QYb-לּ��]XT}����ȳ��_�b6'����<�z�Ҽs���7P̈́ѓ� �Eq�t;m8+9JV�T���;�vj�ė����-�F���pҗ�ShL��?<��e�����U�W��K���!� ޶�ZA���g����C"�d��Nj.�Ƴ�Q��t�0R�&<d��`z�uf����o%�{Q"J�]:!�"|8(�U��o(�����/�j6GU�*!��'VM7�搵��C���А#,��?� Z�d�B��z������z)�P�c�vG>A��`���X��3W���w�KW�&-\�sY*�Eժ@:��5������b��7F�$B����R;3��x��P��t��lK��l�Q��u,��t�>:;0��A������E��F���=x�Ԗ��/�:�(�@�'Gp�Bb"�?�Y����M�$4�Lt�a��s���n��1E����/CHe���f����$�H����;oh���w�)�u�%��atN�T�(Y��m�4��@��N�kU��K��5�� 4a�9����M%l#����:�b��V'��n�>L@V�(�XO�+&�yٕ����wBTJ�ʿ_��>�!�Vt%K+����t���7pP!����<C�vc��S�}����B#��p���/��~R��z?h���2w���N�'ޣ���/�)����
��ݝ�k� }���xּEwlĖtLЏh�Kֻn��Dե7�Vo�7��Gcѡ�g�1!�U1_��%�k
J��q���&�����B���Y��y2O1�����:ְ�����d\M�B�y��χ���K6�_�[[N��9ݥ��!�S��1����?�8����|:8c�~���(���w��ܻ�P����z��KV�J2z�fOx��8_�.:�@6��|�ؕ�$o�`4�}'�m�څ\�_�xK�Zx�+�:!uʆ�b0��{���h�´�"o'�B�i8���b����{�z�혣�2�n*��a|���Xan*�܁�=�m��bg��`{��Q~�8g:��5�z �U�E�_�{�>������ x�pź�?1��}��JУf&r���C,�y89�5���3�(4N'Qv�=�5-��*�����mI���,,��UHg�z䍐�����W�F?�9� !y �����#��s|K�0�`)t ��>HTJ4�}��āj���s'�މ���x$)�x�t�V���6��3m�F�\,c�Z;�4���1�<�� ΀D��F�{	k[v�p�U�
b����k��5�ʖ#�Л�|`~�v�g!�@��H7�,{Y.����q�Q�k��'���>�ʋ``w�/v��?(�U[��U��7�G9�ߜ;L��5�<�����6W:+�ѣ�,�N1�^��ߚ�T�Ŋk�]Ⴭ��:�Wͯ�fP��R��o�����0`,�ԥl~8�
O>8�}jlߙķ!�4#�j�.��;HH��m��+8u�2X�C�� 8��Q��-R_S���t˹j���;���a}h�R+t[��i���|�E?��r��H��"�����Zږ� +�G$�\޾��`:�k=��נt#;��*r\_[��Dh2���������c���|
����W86�&np��)���� )^O8/ C��y _G��k�^�2S��㾘z�7��� Y��6^=�%o��RqW:�q����s��b�˟�CóH���Ŝ���6d�e��:�����Ƙ��oU�KL˂Q&2���U�K���%�Lxu�:��e  �C ��]	7$ >�x�K��D!��!���/�N�"�����(�I��`�����ؐ�n\�).�O��M�xꌅ���8y�e�~<�>��v	df82�.�r�yd�gL�?��H�428AW��R��,�mOx/bIg��_#@)��DQ�C���S��oS�) ��/7�Qt���z���@,�]�YHM��Y�lowd�&XƲ�L��;����~I�a��eŪu�~v"�~��1ƽ`?�3���o'�����$��D����E�����҄�>2��F93y9�y�;�3���s�Q]��_��(mF���:��r��BGiO�����At���8F��3�<�h!���-]���@���u$Z��M�xu�{�Y��`hT��S��[��� ���W��0��f�y��r��9$�<�k��-Y(��&<���)A�1 ɗ|T����4�	�E��o�8s�}x	پ�<?��z����ŕQ�2�8Q�[�r��2C5v�o9l�o\�ݓFI�T�˔p.��
���"��*����д��.P��B
���n�Z_�(���KX��3�p�nC;��c���ȠJ�	S	���+�P+�iaz��W����㺂@�
"N��ʈ����͓�=��f��
p�]2����C�S�P\©��x���y��#Kz�{���`D\,�߫T�R 3��Ye��@XK�iq���d��&��8�*!�l3�G��~j�*���,��A<����@��� 3`�X���N`�."a{+���YY��E�X%޾$I��7������N�y�4�ru�}Q�	��0/���U0/��b�8&%�0ßlV�= ���Pud�A����r���d������O6�����*�t�M#V7��A�^��TJu�k@ǅ�{�jNf	��N7!�:�Y�h�y�*�M�e�V��m���S���q�Аj���~N�l����>��]��.u+.�x`�V�=��r#ʐj:�R�Bvu�M�|�����T�ſ��C�2���wl����/�S��i"#�-7��t���ۺˣ�4��nQ8M�ի���v�nu�r�Pt:�:�-r?�\?:R�ZhHh�W�,�;!U����P�2n�8zR��?��t�א�wr��f0��6�9��=~��bv���E�e��&&;���b'��#m
�4���H����8��U�q������M8�{��O,a�c�	�Zn{�Ƙ�9xA���5�:���t�'���O:����l�.�F��S��kT�c�C�yZ�s�s^dh�R{.�����4i�q��H�T_��n��5��C@Z�1F�o��|q^ _	e�]<�=�R�*OM�M��$��۶���zгl'xu��;_����_7�bX�9���MB���87��m�>��������ݾ�u�/[�+�^��ź�]�Z0$��|%$F�]n���r��,HB�7���Ւ^.������)�\�}	m�{�h�F�R'%(�_�Gޗy<%���&�G������W]_�@�DaN�FQ�g�"6�rY9���7�|���6@�#l-{�JlgC?����?�2@���!&�W<��J�|�!���:4�xs*�Bl��?m'�pH])��l&^#���G�-�春�	�y�ו���
o�*d��<��m�T����Fj�A�� xA`I��uY�B�O͈�0��p�e]C�3���~�����Y��f��V^��z��1���UA�y��ăE��[k�U۵h���O�4	��tه���E"]S�x�U���T��!*�,�=eA`͖x��ǥ�b2��F�"���|*�<YTܷ)��c�($=�}p'S���tfxLb��&�=K��� e�Y/0�({�2�g43m"'ϗ�(�҆N����K7P�S�0r����Y7�5r�pR��z4i�Ab�U��kW��b�bj���/-���k�y͆�]!n�ۂ�ľ�{?܇
�d���%��G��'��)��4��e��5�_F���>�	���J����ʷ2q �л�����N����QHqA%���f�6
��l�즚'�H�\#�q����F�hc��G#)li�?6/}�m��Y�Y7=�=Xvp�֔UO"��AS�p����#�7�}�|�ߵ�7�C�q�=��{|�(m=��u(���E�BM�>-�g}�x�iN)���_���y��9)�q�]`��HOe��c��z��J�j����
b��6�Z�%����D�����*�x�Y�V��?4I�FJ�Zk�"������6e8˄��<���8u