��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��ᕫ��H��gq�f}���+����c��0�7�*�y�HXH�+��Y�Ar�#�<�k���bu�-��.���O�;����b���7pE+�������v@��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T幭xX��8�hG��kr��'�n�IK�v3�[B���fP�e�q���7V�&����J��v�(� ��n^�ӄ�`� S��JK��W�|�	�bL�Ԡu�%��x��@:���Vì���Cb�ƈ�x��tHjl�!!E�쮸-R�uD���`ꗢ$X��%ʀ' �D����NQ�G�v�	x����C�c�Q^�T��ȶN�I��:Z�ޮb���u��$����u8�������<��=,�=�ߘR�7P\ȇ^Sl5��?��#�3��I&ug��F�@	p� �.�Ŀb�Hωg�t'v������fu��}�̈���1��N�������]�f���`�jX���J��g _���(��>t>=<���:c��!tlv��$��Y���S��ܾ���ݿ�b+� I#c��U/
#;rRB���Wx!RC*�ʋ$���א�e*ξ���c$oh��A�qï�[��a�&yc�rd��w��g��!f����}!�L�Hn)�0�D[(��-�T�B��fhd����3 �[b���ѱ�Y_��o'X�+f�>�>Ǡۮ�hP�)	��)#
_�żt^���Ө�a�����tc�p��sd��(�ztf�l��
�':�A�S�-���5dY�F<[��=�ܟJ�F��ĖY�S!��<(%�0k���p_���P�'��V�]��f�Wt�����t��.94Gȁ��z%[��r�~��6����m(h���O���-�pWq��$�p6|�ӿ%H�䐠c�l��e�Q�҅?�g�2�	���8�j`:�7�;��}!�v}5bx�6�����%+�*$��Rc�����A)ռYvb��;(^�9��vL����by$���v�!.�nq�@�3^ �픿T"�� �c��f��b�JπC4ӐXW��(w������L��q.&;��W�Ͱ"˲�����c=|"
���"��-];���t���D��(�͕S>}�m�-cc�a qW�To����͗��Ж?��LN��QY&�M�⺰�p����m��y%�&��ny�0f	~�|���a��Y{��i_}��5�D��n)k��R*i�p9ma�cz�8o4#�'���p�q��6z�cW� VҨ��99�d��ɏ�6��E@�v�x��h���
�x��IW ���N�9�Q>���^_@*1���F�lx�k���$���)^�2���T{���e�3�
P��4vi��_��|n���c>�W_K�>��	�YE9���=�_�� �O��/�G�%v=����:؏T]C`���b��UԱ�����g~g�r�=&+Yv_�+�j�8��QP~����������Ғ~�.p3c�%����^E�L�K9Y��R�H��eg@�?��o�A%F����ki�ɶV�Oqh�c�I�B�1���1_A�� C��9t�(��	�xl�Q=��BmeJVwL�
�q�ݞ6X��o��Fk6՞
�������༗��:�[�<�5�3�5+����?����y���RX$i��g�d��ь-��#Z��[�ץyv�� �I���|�w�P�H*$B���4�Ec�}n�zX���~������8O�u���ǈ�w�F�i��s@^���סSN<w��8�&�uR�h+�wi����0~�o��_�"�[�G(@�z^;��������!����O�.;$G����>4�8�X.���Wk�,ٮ�f�O���K�Pj�"^i��(v��)�k�4S��[����;�5��[&y�;�N�kY lx�a�9Q]>���."��o�]��cMGl�Sxf��~��f
�Q�9�J�1S�o{}��o_+vKQn�ϊ��k�bu�	Y�)�^j����r*�;�.eC�0��ޛ�e�}	�`$�#�UwT�A&9��aM�%}ń�����ёp	����N��#}�Q��[&.i�N���u�B Wӈ8F�L���k�ӵ8U8�*�;M�1�.�lZBk����X�w`$�*1�(bT�s˜m��J���*�kz����,�k�c7��.��c�;>AZ���9�R�	=Cz��t0�x�ɺn�y�d�K�^����Y"��'�\(ifC8�z�>C.�B�Z���	-�Hg�m|�k����ߚgd�1�:t@�A��_��=[�A�h��h�R:�r�nK}c�A��%���ጱ�qFH�Ls����|�sxK��1�Ι1�g�Y�ʚ
)]����1}���f7=�-�=�5$)�#�r�սqBr� J��6v6\�]��f=��%BVSs���3C���{���c��J)�> ?�-��"�G�]X���Ll����f��@�*j�C&�d9���?n�0.�k+����ګ1wNflt�&��6����ȀG�ݹ�#i|�Nx�ޑ��R����D�eo)m�l��J蓝~O��	_�d�_2*����
��:P$fz���ݲ��+�����-i���_�pI? ���	��K_�M.2����.w޻���h�T�&:�oFú`� dW'���w?�/#��·[�Y	&R�v��f3׈*�X��Wܲ��Zåh�<�*�YP�<�G9���Cl��<��x]qo��)R�7���X��[���by��֖èȷ=��р���k�]�I�!��*i6#���㜈@� ��EN�0`��kYa��F8��+�W�u�I�������Q�g���}7�y�H̿�9o[	�;
0�غ�3��OŝlNx]��+}��"E���A���"�@WK�fFK#+�	� �ilG�Da�J�Mp�w�@'���I�s0�L9B�����wxhg��42�e�l�Y���Q����� ⭔�Ym���E���E�/5I~i��8A��d��M��۪; ��������Oю�*��D^���A<�ms ��
e�������x{q���Vn>�^+���;y�] c+n��4����^=/��n��,��� =�=�)�`��ϣHay��޾r9vww}���}e������:'�S\�Cf#��{,���m�\�(���1�;V����HH���k�8.���+�!��]���DqChU���)3O�ob�H���P�8�v9-�Q��K6��D�t�Z��ԝ+� �u�Y���P(�YNGNjB#�/o�����G�a2}"Q��맆5q<�,�%���_*"�DG���^�r�zNZnb�T�ߣ���Z|�˔C
�ƴ*�\�;J#
�X��k��==�	� �?�F�Y�ј��&� �H�O�ˡ�j���%��G�m�Ҵ��f��uy�L.TIi9����9�u��5ۓ�V�`�m�̸"�X��q�3�tR�������EՓl{�@F�/5w�D~O��FT���Dc#)���ˌn�' �a�À]3h۽���-�D��5��{_���L5���ы/�W��<�ӖJ5�6�)J;OZN��|Z��w�����E�(��ϴ<�v߁Xf��.;&g E��fB���8��Y���n$�M���XrK��u��o!>M{�ue�����X�'p�s,�c���53�U�뿮�|W ۷v�ԏy���C��%���|�������Ը-��p����	��7�w/�Bb���!o�_������SP���5��b�-�L�݉��%0��	n����`ݚ��t���g�S�n�N�w �Z��5�`(V���}�<7�ÀքJ������ǋYȨgf�p�Q���~�oqĈsJ��h.u�iܘRׯ=h_kjk�S��b;��`����j�ъ͓�TYŕ����n�p9@��ժ8����۷���}�02#h�̢>3�L�?�LmqZ�}[�����{P�k�k��=}]æT<�������K1�8�X�*!/ѓȸ�0F�h	��	��$����Yƃl<��g��,����ǻ��o���cK��)��$�9j0��ݺ�1��y=Yw���"����'7�K<�=T���x���-]��}h�,�{��QL/e@��ϙ���1p��K�DKs�
��\$!P�$�;S;)s�a��fM�2l�����^!��XX����N��zbb�ٜ��e��B�4�5��/�6}v��o#��t
B�X�0��9�,P|+�df�]�/�B6N�w��=V{���ԅ��cZ�r�_'�>�����l5���($F��Ћ��0C�R�4��M6�]��$������/�/��q�}jX'go[�������oE_@�ʑBG>��]y~��3Xe3��e���3C�.HC���V!1��T]p=�G���b��@��0�?��Ö�T�[-��d�Xt���@�8�G�/N�eR�^R��)��/�#��U�V"a��?�z֏n�ݠgkǓ�JלYb�����)��۵��Թ8���(��P���	�w�mq�W��W/�ڭ��Z+�y�DÉ!�2�jlZ��R��j���ݜ����Yψ�e�k�!�6�#�fL�̜I�Q%[�k㰚�w�ԉ?�6��t¢¦$��/����h����E���8c�ȓX���|�MiQD�F.^�$����Nu��y�RS�@�l0��]����W+��fB��ژ��E��{�ZO�ł�� Q��b�!�������X�?�t��.c!_��	�,�a�I�V�� �:��;�8/�9��b�d%��s{��J��Wf�ֺ�B5!f�0Q���1C�ȗ'1��/}����� �A��&D�b�(��^&F�Ѿ~@#4δ����o���s��)�-G�\��;2s<Q��5ʝ�p"}5*W��I�T9Z�*��r��%�c��.����5A5�W�`FR쐇-��F�f�-)�q|�P $�?��կzs��Ⱦ�W��In��
��##���	��ڬ+Q���3I�
K��&u�����oت ,�*۬Mvn�Ap�֢:j��8���e;�]1WX,��&�z�0d�7b���m&��P����� �B ��2qٳt�['�
tV��09�P�6��(ϐ���"҅�@��%(��`]4��NZq�*�u���/f<[���N����R�')'�����I��rO<��S����%��cX�-M�g��wsO<924��'�j��(G�����L��7�N�	��9���h�ԧ<~Cv|��'���,�-��)�V��¶9԰�hd� �Xy�lJ3z������~�w�R�Y2vf��$0���e,�� ���������>W?8�t	J����g߃b>	
x:�l�L�n����.3�us:�����G�y����4��oL'�~]s=�cԎ-&���X���������=M-0sPݺI[��'�b��<]�:a��@�<����Vp�LC�!�RqA��[���Oն/qp�.�8�D�	j�^���z��e6!��CS/"���J!�`4�'�G�A�
Ɣ�e���ٽr�Sn,��z���%+뙔�v���J��5���b;
:	����"3<:��&AD�^~ �,�t�cN=��p������^���}�p�|$X� ���6���S߯{,K����.w���@.չC����7I��c��>�P���lL:��n�eh^��2��� ���e���bU"Ca^����H�Q<o�r��S�A'���3HH.��9�_{�BR7^����y���K�(���mǚE@(��6Ġ#����1��0Q!McW'�� ���Z)����̨��2Mv'-�+��.�w�ـ�H��{���Oj|=7xT*�?&���;������O�.�Dv3(�`B3Ғ������� ����ȟj ѩH��	�� �Ȃ�h%����-`���&�A��[�/Ty�Z>�`ؕn�aH�Q/0���[��o;�����_ˢ�!M{!`��ɯ
���N22r�?@F��0�� oR��Q����ũc!�D%�C�}���A�L����)Cm����@��8��́`�Y��I���M�t���[�t^�_��۝;~ӡ�/���^�;u˻�$�Q�{N���^�$
#�s1xE�����4���� a�O-ՉÅ�Ē0�*B"�M �Zb���_v��{$������V�����I���i>_�p�:O�rm�F��,�{6��RN=��S$����9�U�B	�J-/��/��ru$���]���̍�𭆘��KD���1�� \p��d��v�t+0����}#�å�5�Bm�(��SJ?;+'�Ҵ4�c��n�� �:�U�����T���fr�:���#)�"�P� ��gY�e�gF���w��SzB�0�����ʏ~�;��TN=x�.��Q$gl��<ra���3�}� =mi���/W�(���.��. >�����Iw'��c`�P'(�\<�71�O��3!��H����.ϰ�$�{��=�c������W�M�	'�w)�9ۚ-��$LD��'�.�rKm	�C�<�[��[]�ϔkT���\;_��R[t�鏚�[�v��Bwǵ�w�/��lC��H��(~��D��pXH4z>|��\�g:ݝS��)U/=�S����9 ����(ά��C �[�O��S�'.[��.�È�#��\2{f�ct��S����wr36�U�� 4`���6g �a���MaO��I ��E��0 O�=:�;*�0���T��CwkC3��l�wۥ_w�P���ol*�	�e�{�E���ɶ�w�b�d1́D[ڤ��;���@��Q��"��T/�����Q�p�)�G�#��PI�gy��ը �m��Q^��C��]�q�o�Ģ����+���jP�+�"^Sj^��f#��k�/Ix���'J��$�	�ؽ��\wg�\��37cL�m��'�>�,2���^H�8V�C^m��v7��h���c���E����aa� Eޙ�Q�0 _q>����lawq�k1OA�*��ٹ"`p7�i��2,������p��l�+F��$�{m�3���#�ܿ�6$��>e�9V�|4`�&y"���F����Yp�����]�uOe����W�Y�X�l����~�P��O(��c{l��z���'�9D�bn��N`S����d�"�����[>��,6(�s��Bz�Z)Wo�E60�,.�}8	�=��$V����QV`�	8�!q�`�f��P+���%-��Cy��'rR�{&�^X����ƀ��"�0�0���d5A�
q���0r�݀��h�J��d!&���aycyc�A9AH�ӏ��,5a��#�4!Q=��ݫ3;2�?��_�򢁊sѻ�$�����P���bߡQ�� Go����g���5�<����	1��-�z`��7��_�@{p���N��r� !�r����C��;+f��:��Ģ͹}�>E������~75���<�z��Ul�kȢ6	-�=�|1уx�~Ӣ~ /.2���;��D�c��c�>�w��t����l�������q^�Q�0���ּ$~��!�g\����f�a�ϴ�6�QG��Ɗ36�\�ڙ��^&���*ĩk���)nޭ��D8�� 4'���6�O4��ع�+H����Y�� Wa��@*&���
��p��`��y} ��&��N�����`�2�}��װ7\	{���i+��2�K�$@z��CY$i����8Rb�2��D U� \[���g���������bǴ ���:��'�]�Y6�q�*�{"�� y��e��Y�'Sh��}�6�mW?<�o#�u����{��i������99�*b�S�W1$��Ѭ~�ɌfI�o ���a &��Zf��{70����tl�n-��E�ck����*����Vc�.?H�Ux�C�:f��o�r���������آ����[L^����S�1'f�'y��k�N�7D� �w�'f��� +�s6I�@����>�`_�d	�0��_ ��A�Aw��TC�\6d�tr��A�#�m�éV�|u;@j���X�irG��o��SƤR����2�+�:�W���Da��иWW+$�":4a���	E|��wԋ�I���
�NT����*�.B���I|��ҕ}�ԫ���P��� ����Da���+�j�b����P�X�=>(l_���*xCۨ�5� `��k����O�o�= �i's�&\	�d^�8��PU�q�|�{�鷯�f��[����|�P��@�
�{��VP�� �A�Zr}j,��E�� K���o��u�΋4�?2�WbW���L�6=���!�Z�g,FK)jΏ�ckq*�ʕ{ae��#��	$'��A��%�>��Y1�dչ���i���\��n�a��N��U�Zx���r�>�\��8U�_o����Ŷ#��T�% 7 ��S
��+E��hC4k�o�&�
�m0:����w%��CBa��		
�e̝A�<�`Z�M=I��W�~���=�Dr9�"O��ˊ��a�	E�&�]���{���u��P�Ms=�+G��*�O�w��	X ��6(�4-�7�Y���[�	�(KE��C�h�YQG9��>��XKb�?<����'��>��F�¥;���J�D�^�4=�8P��NS��V.?� �LͿ��^P�\����4Õh�n��;y?z�4�ɕ����A�%�#��B�1Mq�9c{�w�J;�ҩW�Ny٥|)��� �e6��>�/�;�<A��h��������a����˽�61�]�,���e��N�Aey�ԘK9� �>e�����b���I�	�����6�
۠A'|\�&�l��\� ��]�*.����C6A� �6v߃�9��O��
���I@VK5l�b���<W��R��;i�yřϛ��/���)�1��Y�Ef )��y��$g��|���xQ��*�4���/_����3h��~h������IN;=`~�8(T���/�)YZ���=wdZ��m�OS~��V��%f�M	?�_]��=F��Q�*gqb9�5
;���i�BN�,`��Z�l>�T�H�
��|Y`0[׷`E��2�A�%���&Q� ��I��7�������.����I�^�"׉�����! �M>�<����E_0)_��jI\H
^�m	�ËAyf+9������т����)J/���q�ܞϥ �%a�U����)������#!>|���jW@���u޹�a���L=5�Bz�i��l1=�7ʴ�k�׏��G�m��U"7�{���9�V�|��*c��~�o����l�M"�<�����W3]���S����T%m�M�pj�^�z�@1���<�)>�V(���M�d|-V������Lkє��7��_
tP˅�)�@v q%/cA�S��3B�)����S���z�.�y֌p~��h>趷,��k�1��0�m�Nd������~i3��ؤ޷�|k8~��9?5�kҺ띱�X����b���D��nc<y��_,L��3,~��:��6Т4c˃ǿ��1���Qi�D�P���n���a�m}��у(Iābc�cjy�Zl(�i��hPź49�|h���3�q�Zd-��ZƊRY��q�YBy�+|ly�9ť�GB���#��l�t�������o�%�r��y�ڽ6<����{���l���}��6�����uqwU�?�l}�ږ���z�Bq�E��|���������~�F�tg�\��-�n�|G�_����J�!�1�� s���/��s��[�^�ѵ���}^��	<YchL^��:��ޱ+��7�Z�C��O{Wz�:��bΫ+m�[s	:7:��Й[��6q;��uȫs2�1�� ض�����G�^<V>�@���������HsM
"��ΎV���+����))	���L��^Y+���a�\f���_Qn+�7�:��ʜ��Ëk���KS���[iղQ��N�O�8��#�X�qM�I��+X�;tR�!���ʉD���j�q?b�<Q=��Z�J͗H�-���C������*�))�I*��H�d$tG*�w��dF�*ž��;DK�4���T��a�m�0��Z��l�$ݦ����ͳ>4>��`*���}Yn\fY�/��r:����=�R|��u����Hz���^����>���Ad�gk/ԯ���ÑC��h�N/�pz�M0f_��,��7T>�:�>;�G�6@�S	��O�� Ό5	@����M��N)�/��`���y�Gل�ި��`U����w��h!ws��)�b�����4��_���>��)�)���r��h�)CƢ[I
�.NI�����|1�G&���p�0(Z��P�Z���na;���q/�X�'I��n�';�]��S Y��tX�΢\_\f���j^Y	_ G����xk!��!�S��V�*�:Oӡ� �ܤ`�5��v�Vz���/|��`�8�Ѩ��WG_�Td��;��2%������Ne�F��"�l�0���)K�dt5��~����5��9F�Ѷw���{j)l�o�/V�Y ��)�.,�	��䷘)f���aQ�W�Y�y��c7���$��W�&��/j��}��U����s���*k^mP���{�\��ƀx�p����ከ�;z�
�h�'1��ђ )ٛtP[S�T�!�Ս˗�o���mf@�U #c���&�F6>Z{�z2�w�J�]N�j���O��^��9�H;��yl�.�Ix�=�Ǧ���.��[|���VD�~a4�����B�Z�ՠܵ�(�����I�&�|t�ϖ�m]�YA|ćl����Eڽ�C��~]������I���~ d�D���ɞh���0GlZ��@���>51�h����5��ǷC��Ƅ��wl�%<I��� y���G�]U���&.m<uL*N�8�/6E��3�/^�%��>O���KnEW#]��E�?��b鱏�iM�L�B���:q�������QW7�V�W|�����Y	-E'�ZVlE`j����d[�0�X>���aY5�u�4��#xH�MlV�[�7��z����v�?�>m����w��H�޶�Z�OC�>�*ϻ�����mN�oi����"G�bǪ�L��S�n{SPLq�?(���T�0��x��l�N�9錔M C�8�\ʩĢͯ '����܊t�8s�0�IŹT�z����eD�k��n:w.������G����8�������1$����085U$\�0����o���T�UbR{�O y<���(�V�f[$�J�k�C��<I��Թ4	0����.��6��/�-�KT�5J���Z[E-6=Y���M�Ivi}�I��?���E��w�+�>���y��P5'}��j�p�>?�_anc�@#$dEh�-IJݠ�)�UpА�u��[��/��m^���nP=�$�/_�O���g��L�#�P�f�wor�Xv��.+w��M���,j%
��|Dq��ln�g\�"��<�+nm�#������,��Y���R����|:�2�T����{�{0���B}r�T��gY6�8��u��� �=�����Dt�7��B_w��	;�3��[��D�������ko���T�
�`|�`�/���,Eʔ�g����� ���^�����ʱ$x4����nN��=9o���\bm��Fν<���3�7ѐ���ٝ�8Ƨ��.��XR�����������J��̶��AݬȁM3̺ӬZ{-#ZuTY��UFq�MA B��e(���<;˽O\w�+���)b�G�*~��N�i�5�=Ӂ��1񢞵���)�q�/��Pw�a������R� �v0�^K��2�wL۳zհ��}�p_�'nP�iZ�M�CN����o�qBi���!�J�x���Q�БR�e���Ԫ�j�o�v�X�h`�r���:�qIA�.=���۪��4-)�h� Z]��xW�R?/��/y�f�47�jJ~U'�
�V9�PQ.(�=�}�U	 ��ra#��f���j*]���T��ٮ��I���W�NdX����\��V��m��|�}��^�<�5T���%�Z^�NF����YF�tC3�E���'~X��K�fz7�$l�{$ѵa9B�J��ÌmU��
���5�60��kD�����"������/XH2���pt����}�r���㞲��GL$���}�b�k������KX��*��[l^�>�}��`	r�̮��9cc|�HJ�d�o!!�Q���.��sQ���z��ð�"���(	����5���j��c���=�������][f�����w��^4V 6�������7~���a����I���`>�ț��v��^9iδ��BNZ:l\hb��S���~��V�OP�o}CoB�d�ρ�)Գ%	�[�JSؤ�d��bh�|�X�������,�Sf�O��{��nIt�)��T�8U���7�xU��w�-�"�)j�c��T�5r��u�0�%������8'**t�F{yG��L���jo�x�s4�Y,O]���Ǻ=f:��	�����>줵U�곛?*��F�vS�� *��5�"�z�h�'̬��~��&���5 {�����x�$��(�,x����ك�^�!Q�ŝZ���V(�x\���`��p�O'�X���<J�h�g�kvcU�߭��]{��%9���k�`�|��u�r����ڊ�;\%�=L��O�wV��޹v3���\):��ͮ$���f����HT�JX3V9q�� .�
��Zj�v�&v�����Ŕz�Ŋܓx�̕��G��9X��Pv��o.�!}�oQ��ю���O2.,����92��y�P��5�Պ��	�ThI. Q�vQS4̭Z�Lˆ�oP���}�A�w���/�ƕ|�&����e$|�7���T� ށ'����?��7��<$Їx�z�e 	�Of@,��1t�[�U������",�Q)�!��u�z��_�&��i����>`��$n�Ο����*pD?��⁲��@�|[>�X����B#�Wj�]~T"�<)|�?��/J0K��\Rn�������)�Uh�Mi�߽��H�Y�¨�<ߎP|��g{�_���k_?�+}�$�i}�w_j�|��7Q���^}��.S��  h�?�"Ӱц����.ybӱ�g�&w���lf���A�]���/�uq�+K��;KX�͞9�vi�@Q�a�nxk���|�v��\������[NPR�o\��$�J�T�kN\�O�|��!���a��#�(b��w�\��4���R�`Vy�e1��	��+���-��w���խ�e=������	#���?7[>�3�]�'�$�� _���u�J���W�	|&O�B�ru�	�X�����9����#8��ٽ�q� WR��t��Y���'*ڂb����/�P��QT�$�f���yt&	�K��Ɔe�NE�Ph�_�2�&@�>���@�U���`�MD\/UІ!$<�6�݌k:�����Yy��H#9K��_'��G���Ax��h��f(��N 1r��tn��|�]S���&�	�͕�N�����|���9B�͡��KU�䕱/9�����'9����~i��y������W0�������!���'\V����o�Oj�e,za��J2+e V��>�r�Tf�00CLt8	o� �0�2���k����A�J*d�IIٸ����X� � Z�#x�J�Я���
�{�6�p/K&��K����A4��