��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�s^W���0A��t!W�I�a�D)A���F�`��x����cfa?tFi�zA��EYǧ
:�J�\��=��-P��8h]3��ν�=�!�@�� �Э��H)����������7'b��D��ix���X��e�Ł��MG�!v�I*^	�����usog��VF~C��Ȇ��v�L��Γ�
�ӊ3��} 7Ǫ�A��/�vd .^Ɨ��@I��i�@I0߂N�59�֕���qц��0�Z�P������ۡ,^���,f@oD�%�����1K-�uF�
$-��خpȃ-��ÓԈՋ@8<�|��u�/_2tQX@@}�2�Uf�׆	�����>n@����.�75�%��)?��`ԺU��$Z���zr����@=��v~w�%��c3TV��|-�b���d��/������jn#��B�đ'�� ���T�~R�k���iy���_�}�c��8f�]�����uf�����hP��DV����ykZ�6Z���IDD�>��浙k�g�<4��	��VѲz׾=:M�Z��ƅͅU���F�^�5����-��]e��5a��g�!j���YZ�ʭ�I�t��9Nn�����woV\����"�<^h�:���0։�Ȫ6�v��'�be2��|e����'�R���G�7?��!���K��,X�F��|d\'�	����s�jG*��ז��}������⓻I�����FR����3�����?
ʯ��<8�|�ܷ���Q.��N��t�J������L9:�33ݦ��Uc�� ����giQ�����r�5uR��
�!���V��O�� I�z:�8<c��F�̠x�JX~˸j~'�Yv����c# �(�� 8s�T�WXrB�]4Y�hL����'�p�1�� �5��$�X��V�$�OC��'͕��K��$Y=��$���k�P� ����i���п�>Y�G�m�t]��
 ��@-V�g�d�ycD�X]�Mm�/Z��
�s���x}�1ꮿ�iǽ)Oډx )�2��ྒྷa�\G ��a}θ���V�%���+�T�� �(���c�-��ԩI�`Vg�hv�b1�X�`\C�ٝe�H������騧{��R�ƽ	�Ro�BxSh��`�y:��1:�B{}`������d�b?������c�L�!d�����n����V�7��Hi�G�����1V��%OzI[<��l�6�.i�����3*��a�l��	�;c-�J��"�+�� L�=��D�
�~D���2�:H���@�%��� 2�B%_��K�Tu���[3��$Fߌ��ך �����@����K2���=�tָ�<��E��y�J�2�����z�����E��\*��W��kˈ�ML�<|�����z�}��D�n�N�$IaB%J�p��[R�b��E�.���., ����	%�!���d�O�4~��y�3*p!<*��t�+0u�Nm*�,�5��;�<�w~��"�;Ze��-�̠��?�	3,[�Q��~��?8H�	򿊺H�w��4��* 7�J�������/�����k��4(Dٿ2���rl�<L��Wh��ܖ}%�B�K��FD��Y޽�M���z��FƐ
�� ��E���s�D �c ��o�<������@���R����0�=��N7 �l��?м��� �l���)-�9�#D�i�_I�l�L�����z�y�����Jq�}��r�o���zY�F�+V"j9��ʚm����qGxL�;H8Ƴ�����is���'�kS��@|��_nO�c;rB'�<� ��{y��(��%RL�龜��~tRb^eɅ��!����v�x�K^��� �TaU����w݁j���h�����
юt:���<	�>='�*Uٰ�i�Joֱ	�U�6ґ��qi��&1�Uyx�ՙ��J�<�¢�����h �tԿ_��@��S��#>4)B����r�*3l�&���n4�@9�tޢ^2�8T�r<+��+�rL�A��5�](��/��Q��,�n�7G�2@��HfD;�l�*�EK_�l���x���깚�m�J�2XG��)i �[��j@�
�;�^�u��T�_�/f�%N5�#�2g8�!�1��/Ԏ�7�'7\_+	|�r�ޞ+�5�8�d�w��s��d�*�d�`�WgS����8>���
�%�bথu9R��C�erʋtn�Lo����J�<���S�L�͜���Q�]����#E�XEC�T?��\�m�È�</�Y�֔�|�׎� p�v�
JmQ��,�"�fr�ql�J��3q���#~�c�N�Yr�/��Uo�R� �9f�Y�q=�iD(�y �r�W�%ǽT�9L���] +�
$�������n|���Y��s!�({��s8��o�ز��v�wsAn}� ���������^����8�Z�!�$�w��V�6�X+�E{=J'#ھ�5vr�K2�]�"6L�kH�Z���w�گw����2ȰxӼ��׏�+�H��
���S[m��rX�S`�8�H2:�3�>%�W!�6�^�?�)G�?{Y�Ul_��K1s^�ţf���19�U`�+�x�6��y����=�W�!��va`�^�BB�����薢��^� U���Oa]�7���8 �j �M��~H��
v���SL�`4Ý��,�l�ıaZ��9u��x����?;��g���r!:�T��	�c!H.	�{�写Gd�2���nk���A[\�۱��<�����s��I�\
�[�۴z��t�X
�3
d��C���uH�Hn@�E�N~
_���V�D��`�-�r�mt�]�!>�Z���	nQGl�R�D���&�Ga��v���VJ���IhZɽC7g���ᒳ� N�k>-|�.�
�R�Q".�nL0�`I7:M ���J�y��`�T"�pl��O"�^h�T 2�&��_�H��`�}��o���X�AӴ��!>	��/;d`��T4I��j�;�j�F��;���7 ��(bv#�h�S����vTa���Π�dCH��/���Z�Pػ�'.�u�L��C��<c�JG�G�v���J}��	b"��]}B`��t�e�����a�+��v��d��`%���P����)�蟶�.'�p���S�a�����!O��*zW�Ҽ��ƣ�����,��O芪'�E+�9Q��,"�դ�S�~�#��u�g��'~�I����H���x��hb�ѢEK!H9S���@=���.H�5�������Y�
$o~a�>z=��O"��2'&����>��d��3��T�g�YbFZ��za-E�����m�t�䕺�g��{��y��k���0c t�e���b�
�9ZȊ���e����ʚ��!Qȓ19ҋI�f)X������3`C8m5]
�|{��u��#�dJ��x$�{˩�@ �������T	q�jpa4�PU>�3��X}v��kH$00�=�}|^=̜��T�U�]~����X`J�/��A�Ӝ6$�/���J##���?�*D��jaA�u�j΋!'{}Ѝfr�N��Wl��F�5�#��9��������l��(���{��#QA����-e���a�@h����j#�M���~炐.0&or�ERQ
:E�,�0Zg[������>����!&��3�g�@v��lK��X�����v��)��Z�M0k��ه6����Օt]�3$�(�@9Z�9�ћ-I�P�V �?�D�ˈ���>'>����&�{O��!?�6�K�������暿���4�j2�9��@&�ۣT]Bv�&c��S��?U�T]�a��o�Oh���� ��O�~"�#���]��p�p��%f�v��Wʊ�'����#�?��Ø݄c��9�杍�@Д��r�t�Zy��+���$��K��ȷ���2�PL���\�ߧ�o��s\���k��)�A�&-6�X��Q�k72��ISgU��:�aqJӒQ ��/p�h'fc�����J4����s6\?�u�/DlJW9��� W�<����->��62�����ŉ��*�X_C_���~([|<r-O��[�4Fc�[��H�y��I�K�-�}w�r�M�o���'��\����Cb&�s�7m� ����я:!&����>��1|x�?�{�)�N�+�{�Νt-�-K�<�^O��o@-�������#�f��׏?k�J�4�[��ǼB3B#ɆǣGi/������!$�yJ�Gk#u̶%��:U`M<�?g�ƼP�@Cz[���� ���$j]��D�KcP�9cv�^�f����,Tu��HX2G������к����h� ����Ã�2�i�pn��eg
)r=5�c;I���82�����q����f`4t���s�,���ͭq�s36��6�8G���)ʨE4�'vf��&C[)��}�Q���$���r��b
�Q(���ɟ�'iG��z���$�l�%�PW���W@X�d���xP�:��r\�#����1U���ڐ�M�R�� ���n�hI(y1!|�5�h���.p��wv��H��~}�1Y]	@[t#��"���E���7Ęc6�5��Y�l�8O䶏�i��l5�E���h�I��i�dGa��fM�*^�t�iV��[s����: P��;%=��!��Jm&z{1U� ���2y��R�:E�z��\٦��3-@��w����Xn�e�t� Wr�y��������]��ʒ܌|��S��yIX�Z����Q v�8d��c�hc{�3ܮ_�?�Os�YN�<�K��h�N����p۞->(���_�!�J�P�����RMDx� �yda���S�m�Y�dc�l�@��3�:�ք��	n�_\�k�7z[�ؘj���/��+rX�1!7�Z�C#I*���)�ܧ��!�Z���o��ă�D䁣�@��/���m�Vl�y���j�h���g����e��F�3�b*/9��c6����Xn�����bC��f�Ub�3[R"`bb:|"�|d�4{D
I�=B�UO�:�<7&�}���y�/���g�Z��s��Sᵀ>��a����O-*Pr����D1,{>w@�n�Q�FT���8؍5c7��ө��S�)m�m8��sC�*9�H�ę�#��b5�w@
��g�������˜�E�y-�a�����v2��,)��|�Z�A@��i�fLV�r�uK)�hPq�f��0��/�%Ru(�6�4�%����5j���ƨw�����?��\�ͺ���{�`��&��)�uO:aA
����-���1�~|.��BU
�+��U�D�C�Y����rin��NE�m0����=|��-��]�l�0lk�+Ug
�@��f�%\>:�m���[NV�f���$7Jƌ���g�Bl·���)�@t{���4տ��b�rˣ��;�����f��Х�Ȧ*|��3H@���-���D{��7�Q��f�ҋ��Dk�{R'�y/�Et������tHӤ���%kس薘;'zž����iu�)�n0�e�O�`J��Y���r=!����^Y�Y��;�R�P^��T^P�U�f��Xϓ��lR�-k��A6l�^���y_�k��x��8Y~VtA�Ç{I��Ê��1-U�]���ר%lP:�O�%xnt�]�/�<1q,��v�z�d�C^q:9��.�Q=�H�j~cߘ�����ۡ0z��"z�ށUg4��GE��$�m\�^/藅	���^?�%�k�]IEm��9�Zؼ�����������SI�Dl�{�(�K8��&�
��;g��ު�GE�����Au��8��Yf��^�ϐ,�G���yvP=S�,Y��?�1)���
hy�������|�E�e���E=r���cց�e��P9n�y�ޱ��G��UZK�/�/B� '�
����):�}<�	/�V�
L�ò>��������&�m�H��a����0,3��C}t�z�Ʌ�(���&�i�}^@�fM}G����������|^y��^��p\n��3)Y0�>������[�YN����$+6�&\�6�/V�`<��Z�j����[����`�Lb7�uȴ�'^\�,-�G�.�� ������&��8��9�%����p�˷����|r���߷��=�NC��/��!��҈xN�����L��
�\������d�=�D+(Ap:�j�o٦yA��RP�w��%��D�\�pS#������՜n��^ G�å<7$�ϥk�nDu��ךB�׈~难~�K-HI$A���=��#S�@�p,���4-�7����
T��h���+��ct��6��Dn=�K16�W��݊��a)C��H?�my�(īy��t`+�<W��%�����HI���àev@ꨩ�hr��]$��G>~,QY�4+dX�%1<�g$8�3�k���>o:�����#�wA�lԩ0��<_���,�3�6�D�n�l�ƛ#,�S��P��S�Մ<T����(V��*��Q���Ӑ-�땩O�IA �b�Xp������yˢO��;�*�x�6w,��9%�_�r����-����rl�`�u��}�`��s4t®h_r|���taf	pP'��R�_˭B�?��p��4�5?����������6���
�}%��Bf��d��~�H�N�/�g۽��@�N�{�U�=���~#}# �Rk�M��vu>�#�d�?�Ϯح���������w2n��w�rJk�����Z���z� n\>�bc-q"9(��rUJ�*,N��W�A� z�:2��_�A��B��lK�0ԗf�����D٠xTQ���'�� �Ԗ��w<X�9-d�A�\6�ns�t� \���K%�E��ӎ�8�qI���{ �j����)�� ��pO
��?�7�捑<aǺ��K��T�����y-v���ٯ
��BgaA�N$���Q���r6�\�� 4��9��;L�2�����X2:*�5sbV����3A�%�l�4f�I7��ʐl}��_��:�}š1-�,rװ�;�����> �rԽ�3����d�V�?��ΨlFM� ���_��Q�	W�q�Ր߽���=�_6��	&�9�bR��4����݈����V*y59W����}�_��h�6I/p(��W,ĳKE��#wqs��n������2�uϾ�ʑ�W&��}� �o����-�	���2������Q���Cت0����f�)�W��,4��戳��� �ߞ7%^�yf��xy��vKR@/9 �5r&Ϭ�[H�!��3���-�v���?  �����nm[����ֲ��E�Ѣ���m��=���xSVӕ1t���I���,�y��D�ځu;7�&ڢ��,���-�ES��Ip��(���ֆ���k�)��~�B����CϪ�p�[Oev�}C�U�F)߽����-�V}F�>�P�㐱��o��0�lm<y��q�l��]c���z)�^�Rc���L̶._�G;����a�����,����F�-=���xHu�d?��n<��|�cwҚC6� �/r���_�W3�+�Ѭ
�r���R�n�^ne<�hI�]J}�ǧv���C��Ξ��;U���P�}n�# ����}��P�wR�hM�7��6t�q��% (0xq����� ��_����@�sп����va��?-�Ƅ��\LW� $dk��*��L�L
`�ůG*��H&�q���`�x�_F����fuup���"7�*�\-
���Z�Q��O�*H���=�v)m�ett�pK�߇�E3�����d��=��D�73a���~ml�U�.嚙�p�w����|s��њܬ��γKCFXX�����;ؤ4�����K������J������/^�=âka����s�tb��g��i~���^<o	�IY����S�cZr����љ�'֍{�z��VXeob�$ۂ;D��)h��_%B~�sl�2�xΓ ���nuϐK�sX����n��$tP�\�#{-%UG��w#��%?[4�M��n �V)�X~E��П��9p?���'!����Z���fDq��'p�S�gj�a6�վ��X<i��Q�}��e����{��E��BY��1��2x�sVdt��'�$PYr�qh�(�ru�����@���+q>��- �}^�ϧ�!?�Q���n��9L��a��%Ah�b(|: =��RG��sL�d�ճ�&�I����te����.�5%���*hp���O�r���d}��0������'�I�Rm�EUd� �F@۪�O��c�{��\|����7|�Ai.zi�8�L"Z��z���[�aS8N��c�u^��Nb"P��z,n�֦������
P�Xù2Ξ����B�(��^'�,�uM��Κ�Rƥ$�=u>)M�$�"p���@�=�4���l�i���(��p�dͻ�S#eV6�M븋F�Q&+c�T�x��	�m� VkPK�S�/��~BG�3��J_���f��K�ӧ!�U�r��U:���@�?��0
��Q����;I��uw���y��Y�l�AP��@t��;����y��-ǳ
c���,���@}L������%�"��^�{4C1��� ��j�4D�(���?4o��~a�P������KM�Ľ���g9Z^���������6A�C5f0%��-u����v*!��z�P�����W���2A���X����9���i�FU�I����]$�'JX���+O��@F=�˸/dyyj&�s�cOީzS��\\���_��,f;�kS!a<y�Ò*Η�՝PY�S?��1k���#MLF�7��nЄn�NV�T߁�|+A��D�6l�bGi^��_����?��w�2ca��d�At�����le_�c��l��6H&�^9� �[�s֠,��9�(�<��&�� \�F�2�2~�%TN��(y��$����`����{�ڏN�:^��"7�(kƃ\�B+b�9�L%��lˇ�D1�r������_M)��<��3mt�'�S���^{zJt��K:΂�&�����-��{}iO���4�����dvߍ��q�������o~�����oQv�_��_��jפ�9%��d���J'HI���G=�������-D�h��e����0���@}+6L����^�}�K���˵i�3��-�i��\U�n�n���Bë��8p�p��HL,�}���n���'�Q��%˰8�dm]`8�[��ܾSw��ps���q��j?�5�`��n}�G�7R$� �_A2t�aO�")A��<�3#�{���u�<Yt���Ҥ����$&�}���v�U����-��7��x�X��:��� U9xNW\�%*|*���56�����ֿd>��>A�p\����)Z;C&���3�7'�����BE�Ξq6�����I�0
��E�
}�)|B������W��A�mR�V��FN�m���MH���wJ�9Ef�����j;X�n�AIJ��)�*�o�nD��q�(5ë�Vؙ{pz/X�cT5�j��sp��ho5��d���Bsn�Z����a���R�x��
��Bb����j����E�`@��jc��ul%���EB�jw��a3��m(��st-f���OD	@�9��k��� �j�;�ΊkjUG@l�~[3��ҭ��W�SHmL�yPef \hN@�m�W�Ò� َ-*J1�1���y_����V�S<�������D�4�LW��P�0 {5tl�3BZߡ�3ҏ����mM*P����]~��cQ�"5I�D�8Pg���G��.��P_��㜾h ��ܦ��2�����H#a
Q+CUda1�L���!�ռ��%��ܤHP�Q�略Q�ZB����*n��=�U`�~ x	�!�d�	�3%Td��(���^_���u��#ڝ}����5�V������(�S��!��Ҏ��ʟ��J�rzn��j���{��h�g�9��Nیe-D�<�
L�`�z���0��?�����[�61��}���DWYj�c0<��"����\���ѿO<U<j� x�4�x��-M��*��\�j�;�!N8A�>3��;��pLz�א��!67wo����+�D���(p�F]߰N���N`Vd��̿ �Pa�g�jO�6U����Z��4�v�+d�]�~+�0�1rY���؝C��E��TT��7�9Ґ��Ծl���f��ߠ?%f��8�i���V+�<��_�D�c_w���GT��xw{~��G�����.5��� 0��rݸ�G"�'�S-J1�"Ԡ���=;3�1}�qQh�S�n�T����VO���n���-�܅�� 8l�� %���JL&cU;:�Rn�*����c�Cۑ�Ad,	�<�K=����>�TPf_=~I�Y�P$��*�yc²�s1W��Nl��漒¶ʇ+��H����9���!6��v-�}���`T�B�%�dM�q�,�0��>?����Vѝ<mbQ����������<�
j	Z%�A��� v�d����9���(<K�p;���}�<�A���$�9ln�FZn�R��i7�Xu�
�VsW��_R�������q\��G��,�ʻx���f��Z&Y(�@�I���`���p��l��2)'~t���XdcMi�X�>�(�1bF,��'���4��+%" D���ĩ���'�"�F`V0Tv"��K�x8��gp��*�x)ާ@��0�XU���3i@0���g�iN����h���)�^��²�^�Am�����S?+rNN`�g��ܨ�iB�fd�ԡK0S��β�3�d�Ԅ�@ݓ��l���sɳ��G�#6��]�6�ڇ]�掯VHH��D1�f�J|Ó.�V��	�g�ڋC�o�/0�.@��˼'�����nj�-^j}�� }.R2��j�si[�"B�d��^f�b�����f����kr�cv�2��&m����5f+g���7�&�`�����;�}�hp�]kC˵o,�f��A����~J�^P7�>`�J��hk�]Vd�,_s��? V�QC�g32n�ɴ���0��č�@�0;7i�>x~+M�\��;��@򲥿H���X�K>�������H����*\\T�?f���i�6�.�T��O��y�9j����9R�OQ!��G���*�j���怫~)JDulw������ny�P=�d�M�f`0:�P<u�Y���=1a���3l?NZ���Լu����0/�P��.y�l�Y�8}�/�eM����w��E�����N�`c�y�n�.�&$@��哮�A|)bP�`$������j��m�`��Q�/ t��y�9oV����j�h|j�N��+D<�6�%/��2�M&�aYNx�jJ2�r_�4���mp�:A����*ʜ(��J�'�콄���.�%f�EE�r����.[�y�P��b_H'�^x�(�p�d�3�`�͉έw�|�9+�˛�c�&���������xl��:����?>�ݧ|k�@��֥��=��0	-	K�ߜ����$^V:L��O��qlM�x�w���t��
�^#�8���յ������'�B��	�.�O$*�=�3�S"{j�wI=?�]tp�W��$/�<;Ԃ~��I;;�Fz����?*�i�Q�lb(�����F�f�z�TV~`r�͡"��xX,'�iq���ڈbS�g�� m�X|�kX��6�I|�0r�+�[�<j�p1{|/�����R������l_��7>�����|��ٌ����/I�c|�f��p'�����q!�X�*��.��"����Y����9�J�Py�)�ȼ,t�cL�!�>�߮���t��ח��`2
x	�����uYƷ$.4�����Tkz�������:[pyh}��jTk�(94ĥ�w��O�P��ܗ\����B��Z����Ӿ?SIP0\���3��gmY[�T}\�]�_JW�D�!nl�<C�)��w���+�N+M��̧�O@���ۍ$�;�F~o	s�����;�EWs�C���k�QJ��Q��%�vE�i\�W����U�<.�z�%�Pg:or����������Vⁱ�[
s�ת�����xw��^g���.�X�]��QŦt=!�Zh��}��0��Ez�y<�v,XK K�k5ֵ!�J�:Z�D�� Z΄fP"��he��@5vK2�{�So=.5�{��-`*��?o1K4��x-��sȆw����u!3q��&�@�����`��`v	��tW;������F@��6b8�ޭ�l�PBB�A��t��W��[Mx�z!?1����O���w�Ҫ@�K ��A�c����l��y�&�[�n3;UG��xk�MA�k�<�ДSZ�Ws0�E��b�R�?���G�T<&x� �ɒ���q)m�H
��حc͟�21?�E�M8��$8S���]����)]���N�c%-5����I��3�/�
\�)Lf7��z��&8K=[���FwI����^g��J	��+-V�=f�E���rA����t�m��W��CxU�E���K�tl��#�ʐKI��̌�}O���w�b��=���[V3>C]�ǘ$�5w�[u0�"6������o�X��S��9��Y��I��ʙ�s���}��^������;a}P*jZ������=�%v`������
rr5�?o9uKe˗0j�ln��4F��Gtf�0֥�O��W�E���eUN6+�/�����22�v¡��SRy�s���	y���0���{Y4yr�����8�,�x���W~u#�c�����ư9�>�d�#�P.3���
ѩ��8�cV�;3<���n�������m)%�s�(3a�xO�فa�J_oO�+���9 ���ߧ���������T�}��(���9��4�MMM��x:GR���K� 9.J��M;�U�Ǎ)d�KN�?E�	��6_kV�����/(U�;_�9�?�;�O�?�E>�nQ��¸C�_�-�BBV��:�S�"hRE��4�I�X�� !���hN	�g��a��Sz��5����u������`E"�sWp��\��m��������iq��	�дԏE�4B�K�
�����7�U4H�o8ҍ��"kD�G�`X$[����ͫ���b7�$o/*.Tʣf^?@W����6@��N`~ңe���ü��*���k�X6X�F���̛ i�1̍��'������U�$�^\�nİ��v&�r����s�M*sSo/�K�${�9�������/oS��#�O>�
�"��B%W�=;�ߋpl���D��.l���^gn��Y��F��Î7j�8��A�v�%�AM|��y�y30�`�v�9������ �ؘ��# �KN�G�\Vv	R$ׁ������^OѻT�q���^ϊv�1�	��,Z�Al.L���0���ۉ��ݒX�L�f~��T�$����f�v���)��%T���x���P[Wa�NOC�SlLP/l ��x,"�#k�GZ) 7�u��g�EJB����p �ƆcO�ͅo:�@$��"�0�六�����?e,�О�4�YuR�yx@��2��[!�n��3لRX"����"A=4�	�ρ+�#���XڬG(�z[���X[m�D�^��,�0$���p�#�.��vFh���t{4��,�
I��AX���_�� {������`�R����E-��$U$J�ϤⰅHfc��U@D!K�c"�9��ؼ���<��'����.���r_z��]Ze�,a�?�u`��Q�.i_J-L���A�gN����(ʻ$X�j�w�,U�?r��h��z�ರ'f6I0��w\SҶ�������6���%�q��N:J�1p<�x�L�$�����p�_')���-�ŷj��@X��ݴ��tg��+�S\	n^�jbF��A�$X�����ˍ�%⃆���\�?�d�!<5QDU亠��9�֑�E��f�5Nm���K��O��vQ��d\�+]�nx�sp��uY�X��}� �z�{�zn�0��i�m�py����̷̎���`�|�K������)�Dm޴_Ml���<�#�D%�{����%̗s {%�%��\.�N_���{B_D��M�m�� �����GZ8�E�p��EU~*V]"E������D�s]��dԄ�W�
}Dx,_4��=Ŷ���z7�P+~ vܿ@n�L�o�~,�X�-\Лm�����Xud���bX�&5�$S��_�Lw��B:Y�7�����G�Xl�����0e��U�8y����N]��Dy<�V
g����	��^ca���$i��O��
Nb�D�E $��Dm7������DP.����2�� ����GZC%��_I+�1U���Ng(�}�E9 0�6��ѓ(S��c����2�j��J��J cj�Ӊ�j�_�A�����v�Y�N�����EWM� �s0\�W����F��n+��@,�-D������Ă2��'�S���@VD����@��̆sʭˤY +(φ�9RYp�KQ~�s��h;E�N�R6�h-ώ����M�*��"�Ÿ`=ͅ��̩h�Ѫ��\��:\0�]6^hm!�h}'�#t�?c7w�c��o}�M�#���g���'�a��ב���b�3�׫uz,s��7^]|��@X�n�q��Ț5%���Q��kP�c��V
/
џ���������깪I��쎬u+�6�jR�� ���h�,Z�},�-��hu�εIV 2��^$x��l'7��^�i'|�ƚ��zDH�%�,��8dT{)7��F@><G������Y���z�X��l]f�v)׊CV�^���@��z;�\��(�1��Z37r��AtzM7�e��ɰ֞g�?k�Qu-'z�A�֤�$V*p�q!^��JG�3rݔ�EVޖY�mT��D����W,d�{���N~��T��G�7��8xh�T^bu:���8T&�2�U��5��զDZ��= nݏ���`��*(%OH��L)ŉ�,Í)N�l���&ݨҬ/�^�9B�Y��k�ت���3�c�Y�	eE�-=�S��/�VZH�V&&���i��<�Dx�4ߋ3�0ϱ�����7Ax%UC�s�C�k�jh��*!:�j&;��m[V��?/I�]z�K��w���,]2&ηIs;z]z���1�9~c=*Gu����\����8� F�j�6 @vh��_&n��� O��K�c�j�����l>+7��r�ե�D|�y&6�?�����H��1�gVQ�jI)M=r6Km�EF�I�޷q+��Os����`Y�,SQ��
t�=s��i�z��5@� ���K�H.�z�D^΃~F��t�5���ce���R�ؗ�j\*[�&p����4Λ�y��h_����ȅ`~��Y(��
}�Y���]�2-Po�L4�{�1�����Ÿ3S�Uu�ȩ�%��'��Y����C�t�j���PC�u���U��iYZ'�f�IAx����p Z+�K�������:6S�)(@���́bA�4�⮦�h�sz{w&���O�����O>�9��w"X�J���oF0?_(8hix>���󟒂&\�w��L��p5�;.����k%�gJn��֔���9H�A���(_�Bj�@UR�}9�ɫ.�ȧ;<\嫄�<?ӵ��/U�mW�p��C���6�#�mك����8�b�/�Y3�ں��6����fN]��s��)��P��d��� �k�Uu:���m�`�)4�gSD�;��J�p6{ٔsO9b=Vum��7���`�U�����~���.��'P����\�<��A-�nqҳ�v��[��װ7���Џ
z���6D~*�~cᦔ�׸�ZoӸI۰P�-ƛ0�=�C������=��llW�ﯛ�=<�g0��@Zb�Ǭ\"- a��&
a�S����l[�_�qBMx�.^7zh�	@M5�b8��_w�2T]�%7��.U�}��Dtaъ�c�9���]��bi�uL���+��ǹL���y�Evdʔm"TJ3�"��q9f~n��M�'�bH�z�ޔ���c�7�D܀F&��!s��bY�lD^1˝T~���tj>S#F+Suם�����g�g��g�	%F�k��U]��%������t��A��g@銘�ma�į�3+����h��X>�g^�N�D�S����2��t��͙{&���?P�ח.�Е�_[]<L�ͯ����Q]�4kf]�$�3�Z�&�t҉���l�tR@�uY�Ä���d]�g3i���!-�nY����E�S�PxJH9�iS3��h[sJ�}2r�*��4�\��l�
�ky���c8V˔IzV�>�-��ȑ�L���P�d��s��N�Ȩ�:!>�4 .ؽkz>���f\��bK���*T3���1ԇ	���(�^��dL{@�������i��9��?I}O��AmST�k	�jX��l�^��K����[Gd��`���I���L��ρ(&��:W�X�Ϲ�h3�d�d�b����Q�j8F�6P�_��o#цұq���~t)2ݲ��,���Ct(���hj�:*�V� i6���Ē+ݙ�i������r�B6��4��Z�r��N0&-Z|����{�5��<FR���2:���ݣ��ߚT�������B��?��jC�5��^R��ɼvo{����՟�bl�n�yzYp�H���=��n"��.������� �8�7}e]���(��KX�x�N�2d��y�k���-��ml�%�,p�P�� B�tp�3��M�u,��T$o��"���ڭ6��'6����1���[�O�)@2C�YI���i H�����ΣFcK����������E�m��=��5N�<�&y�c�,]uD��-ZnZ}�F��A��q��/����ÈX'����@b��9�	�SR��Q��N�F0��$��t�����0���<;�K��M�
�P�D&U��~�v�H��Gٛ�`a�W�
��/z�ٰ���+h���Ε�/�ڡ���%0�+r�w�gWօؖ�0ђf���p:�����vb;ZL�&t�[#��MP�A��b����P~w�&h�	'� ���'+�I���T|{�5h2)N�I\�}:%��h���j�˺��Dv���1W���ӏW���2�I�L���a� _�V�שJˇEh*f�R��Jr���U��到g�&�I�x��|
 "��2����x��w ����?�w'�ޔ%�q�D�I]4]��&et��𖇡n�#R�/������o�t�7��T��\	%I�S��)3-�-�p�4��s��|��.o�%���f~�k�}���aP34�Һ���ȋ�d�7�t
��*4�>t6F��Nm
��;;_d��V*>�j�wXRq�5��m�r+��d�}r��LWG!�CJޥ��ͮc���l���oKsY�_���H<B��g}�7�\���(�K����,0�O�V�N@G�C�0��|�ࢴ�ڷ��Gɋ!�AbI�H��4��^��/D9���G� e��$(��h�"��X�>�[=�܃�����,Z4�1���S�z-zѴ�ĶrW��G�l�R�сy�~�W^%& �G/�u���l�~�?��v�"�X�����"xX�)�Y��ӝ���(�T�ǃ�1ch0ԒǱ8UH��
� ��s�=ۻm��Y��&������L�'q��gޘ�͹Y��cf�ʷ*x�bri$)c6���P��1�1�uu�$�j1Tú�����é�cx���{P�lN�`jTo��?4�@�I�s���Kzh�OR�$s�A��0Ʀ
��bb�+6/�X� �rL��(��ʇ���,��<�0�����⶚�N.0�H0�9u����W*�G��G�^���:�@�S���d-�S�2�
����uR��AV���U��6z@VH�r��P�Ŀ��6�jK_��@G�<�c�k��-l��^�3է�PH-,&��r��RH�c<��?��W���$[���K�V��+Od��\�f"����<�����׌�}�`Ü���j�A ")��C���Z����>�X#@C[�f�@���qb����L�D �[�]\�T#@�<C�DM�6 &�P���r� b�����)��+<C���3�k��Ү��`)��D��k�0rǤ��_��.{#�%��i��~�X~ Q9�mA�L�mq�}2�t�#�mZ� -q6|F�d_N��t*E��	q��Ė�h�;�y]�����g�P���}�Q���ic��Y�%?���u��A��5��Z�bՙ���L�-���y��қ
���@��xG��Xcm�<l�kKw�i�f8	��[n��f�I,���cʱ�7&q��V�@�F��[+���) {�C�ҭ� ��x5��s�#5�;��W���&��a���:��J��b/"5/�cє�J����l�I}3���s5ߧO�� o��eLŽ�]X(�]�=���9���>1�g���_�pV3�M���V�w�6��1בٹ8������M��Z�����|����a[6jUP�dt�8St����ּ�o�y�DYmG�Rպ8��^�Fb�TI�>�� �٘�Ơ��=t���������U����2�%oӋih�PM��*���tH�J��^�!�� �|�z�z��F�[<|Il�l�;޳eN2;�&�.�
c�ߢ?-�$#�@�px���a0��LC_:��@��H�\�(w��TR����6�"ը���p\*9���2~�bs�d�-�>�$�r_������ϥX����C� ew��6@���>NJPAD������&u/e��� C� }2]a8�j��6m���]�T�ԧ1:A�	�T�=���3�t�YH�l474��E���,.��5�G��.q�.Gr�Бq��$ #��r�X�BEE-��DU���+�q��v�uJ�<Yl=� ��p|�*&Ш���R�C��쳖�!jy�⠷���)}����c�x�wT��7�&��V�����ABhp�+0�65|߳㔮�D�c�]�����pO<@�QNR*�^r��f�ei�j\P�Y�Ջ��A,jd����b��m�����O\Ma�p�ӛ���9{�'c�p���n.�B}�){k�Z�^���::Y�Nʄ��-���~*95p�rOS����E��_�����T�IŲ��;ls��n���N�	l���~�!��;��3��/�!��ί�5� ߷��D�B�<K���'7�z�F�+e[��X���a���~L�2�k����në���X?�g�ָ��be~��2>�Y?/iC�$��Թ������X_f��f
�*���O�ІhLċ�'�q5K՚Z�x�Z�F+J�h	�f�`wf�d9�����Ȇ��*��u \�^I��A1�>9<A��e��}2�J���*a��3���q}���t�Qu�a�˶'l˾�:չ�Ffժ��j���pC)o���M	g�r��L��{z�,GuH"�P�
2�F��yG�[n6���~�!
��%5G�hD��d�IYūL�	Dy�\����G�Ħ�4��o��y�
���5z� gA�Z����p�����Qxwb1�P\�&�6��L�ƻ�\�!�+������G���������RIQCW�[�KӶ/A[����S�T��gQ����D�� ʷQc�vڀ`-U;D��=�XF�F 9�ޢn�?%�`o��K�Q5*G�I��l�6X��40��x���#��P-�Q)���W�_�F�C!��k��-m�l,�#$��ć�I���������x��xi�X��4����*�ac?����g!o����X[fTCQ'�����jj�<�(��"���Y�4u& �A����W
0,��嗥�����2:�ܑ���e��:5���D\�{R��v��0���,�1��P�����7����dOG0R�Ա���S�&Н#�U�.Kx��f�6�,��mp������
�T?�Iy��c���qJ6��JVJo��I�S�E}��۲�}��L6^�,#���w��ڸH���4��[��-B*GQ8�	�鍡M*\�م�=|�Ĵ$�j2(5B�@��2g�lZ�VV`�o*����I�z�<B�L��6�N�e���
��n���*��΅`�<��mw����x����X"݊����!4 G�o�P@��6�Pz����c����F�t���G������47z�F��{ ��@�aH&	��$K�� �
�;#�W�>�fx���Z��c�/���`�Q�V�ź3m�sNW���3�D)FA�!�[����K#E��k� Cٵ��D,�>�@���q@5��r��
Q�U����՜��Q=J��:1����TK!�%���^:����v�JJe