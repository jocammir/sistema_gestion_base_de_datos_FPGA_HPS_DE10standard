��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%������Z��B��Z����eS��D���Kg��
A�N�(�a��Q�n��U��N!8ߎ`ۼ<-:[�t1 �m��PN��߭J�]�V3E@m���nf��,rﲴ��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0����c"�JU��_���>D�s�N�	}j��̥6���-���x�4���L�3�(f�NqF�Ґ���X ǤP"9r��Xr�E�$1V&�����0����u��n�\"�ѾB��i�$,�L��y��'�����G�1�@��ˀ��
���qy�+6�І��L�/�Ý���ˀA���Kv&0�g���/������>�j�|(���^��҈�d���&<��!��L_Dx^Y,�r9MT3��T^GrV!���5�����.󫐙dmW!��	��$eсb�f���U�ü��wk�u�y��D�b,Z���*{��C���g�����Cけ:����Ǯ�-Dƒ4�W�
� 	�o�i\�b\�;^]/�)XЯ�^:?AQ�"@�g����.
���%Z�Ԙ���%�sA�p@���MO t���!:�&7��5��~a#�*]nk��j�4���{��.�J��F��U&h���b�s�:'C5'�Q� �m01��s�ib�Eɽ�:��OE�]Jz�v���W?(���j�b��yΟ�3�D��D�`p!�j��5J��h�%,� A��H��l���=KX*�P�k���'S���� F����������Y����T�?W��f��7�?���ȡ�0������X�x���Ț�Q<��Z��ei[v�_<����C��Y8��t7��p�(�T�U�.R�x��d�(^|v.+��e�x��Tک}��dtңN���A��������(��~kx	��mOSK�-�C*?�IN��)�U�yK����tk3ܙ� -f��
b��d�� �Z+��RM��WX�;����2�ĸ��K������9���`��j&XA�*�VU����>�o�ը/3R�R9�?K�Aju�V�s�  kX�Å��ɱ�"��	��C�g��2P�����Id`�R�>�0���MD�Q�����8�9����u��&���7�N�|�E{:��7�v�
��!7���T�nZ����b�6ˊ&j�%f��O;�0(�|��<���T?R����	��d	2M��kD�2`�Ҹ�	���bt,E�]T��lU�e�7Q������;��	q�fS����2p�[���z�s��}��1C����3��;������ookC`I���
�F�Yj��Tp�R5�+I�uq�e�
��s�gf�3S5}��]�O9�H<���M��D�0Ӟ-s�}�jk\ѿU9i���^ɰ���ZE2C�f�����N#�	E	�m%'Z\T�R���$Zͅ����jO(5�D���:�YP������yk!ژru�ua� G9f����7�/���xL��n�����S�d���k�HBQ3�Z�f)߈���r�R������Xi���yoՈ.�a�ss�4g�i�?��;9z��->��kr)��r1�SuGH벻A?���\�%>O٦�rb���$8y��A��?X������*5d���n�7�-n�(���S4r�W�Ex��z���g%C8�$��&)�Oq��8�L�q˚:�?YCN�9Ͱ���+"�{���/�g�}�W�-��9��i���`��LZ�J<XT�Жyh����x�b\O�����p�g
���ۂ��b�	zt��9�nb�=̮S��U��t- ��t����w뭰��C�]I( =?�	��7m�1�/��^�F<�W�������;��DI�g|�a�I@j(�0�d݊7�>@����PE�X�G��@��e�>��ĬI�8�"!�Q�6���iu����8�B����-���^�Re=y������)�X���k^�B\�s���W����I�Z֘G=5�X��!X�r��h?fOԱwؿ?����>a�4�d}rѼ��B����x'=`L����>LULo6�=�[u��/��Aw���:vBohzt��I�b���ӣ����J���J6-U̢��t�_�W�;�Ԡ{��ݛ�^I��1��$h���}�l���Bܜ����CPE-�����{^5'��OC{Y�Ɖ���Z}ɫ)����y
D���>z�Ѐ���d�:�9p���9n�l�����-Q�G�N� �5�ɡqB��[��<�a��CE<g_�#��z��q�,�\�Z%�9�5%���,{�dt$��/�pxV�D�=���Ap ���� �η��p����˻-�ďc`g�J�[���e�f���}+#3?-ͅ��5A����JئA�4�	N8�\.D���&�����_�ʏ/r���\�{���8U�	ލ�K���<�Q1_���u��x��y)�M~8���'����x�z��9�y�G�v'�.b	U夌�R�ҕ�u  ��[�K��H�i���4�'���*#�pd>p�f�D+�|ܡR�CЙ�����^l���,i�r�B��o0��/�ś�	o3�#�]�����=j-W��Ÿ�<~P?�SQP�@k�4\��6S�f����������a���7skn=N�E��Q' �o�_����d�@�7M�� ��?�G�ONG6�v�rtOy�4��ϙ��Kӊd�{�WbPg�����t�PC0��0Ȃ\�� �)��S�I�B���}1*`���S��(��֣-�����j����ԻW��k��W�,͜+ص5-�N~�[�a^)�r!������%'5芬Ph���1ϴ`��?-}I���J/೫����}$j��Q|��?`�z��<�禧��V[���>JO
��W�_;�}d�l\^�]W���pZ1�c_�b��#�z�ގ�δD���+ J�����-�@�|�1h  ��j܌wSJ>g�(���Ť�i�jzl���z+{5�J��8E�蜈6�5/���Yy}�y��hr�h�|����]�1'>��3��h&�Z��� [�;��,b@z���P�=U�
�1^B@���P7��[R,3��|��W�b�� �R�fk�b{�=�i��Xr���lt�p���<<�y$c֮�
di�M�a�!��Bq����5����y{��FY�NrVulǃ�.i#{p76	�����n �v"i�@�U����l���RER46�bX7�a�ޘ����E�� �V���\�+d[��jN9X<?�k� G~̴�\�>�W�r�iuQ�p�S��_ח`IՏމm��	����X�b���Ӫt�6ÿp�r=�����1m�s�G������]S���Qk�Z B��H.��7��³�Z-��OK�(2�"7����������`�|���ʠ�2�5��Ɏ;��ln.� �7D�l��/��_�-��X�%Q��{�+
h=���K/���T�s1t#���#�4yP�����u�9��S4�6�ˈ�A;�\�H�fr �Y8_�)�H��X��c	�@<MJ���%%0�BO��	N����e ��C���E*����A�(EYI��҂{B���I����xS؛yf�wۅ]}o��[����L���.Ǖ�����]q�v�5 ���>;���2��fn(p�Cr���CW�d���X������sBLI)�O�*(zBA�O(����TdW��u���Ѯm�.m�G�O���I�o*
�~��df�Ɨ{��-�]!V���i{�p����+�rу!Qu�����Зk>����c�
�o�3V�X�!n��>���H/zxk���IH k����q��цq:^%�϶��@~�]��w�{�4�����"\�~+)��c�^�gn,Ԭ�uB�C�]Y�Y�7���|�M��c���mO������K��2?
F$̵���~��<��,�-݈�jPл�3�d�5-��[s�R�S ��9��l�t2{	ʴg�@XeRġ�J]	d|�t'EZ\�Q�$Fq�9j-��(^jZ��p��F��:f����M\-0w�4V����#�o���EN}��eΦ%}aNY��#'�*'�b��|�J%�t��R�W@dKD�+�
����\�K0����*�Ѫ�Rہ�����^Ɍ��m��C[bPh�r��"H�AE�A����P���;{i��s䚐��.�φ������+��#j"�BPE�?���.1;'_]x�%p��l�����`�~����Z�_����*�ݠ�5�T�;z�����E����e@�a�k缓�7��N��AG9���=�N�]y5��{5���q'#m����P�h^���u��*m��uz[�SXhu��w�q�ɂ�;�N �&R�躬O������bjh(��N@J��#��&-�9>�;����2#��k��Ѽk�t`$n ��~���tt���uN����*�&S�iF�N$�S1o'Ss�����^�~��>���	�	�����l"��hL������~sb����M�Q�nlJ����K�(r�"H�ې��&��M##�X���Ta��՘���-�duB����K�!cPJ��󬃺���x�x}��חH"��dϧ����9�-����[`׽�z@8���O?��Ī,w��+����[��a��{]V�(o����ˬoE��w�+�K>�Y���$��7��<�K�"��[��p-�`��)!I�#�*���Y{��u�ۯ־�,�5R�9�۴�',�q?�V��x�_��ڒ�Iٽ�U����b�|�Kh���ؠ�o�Ҟ Tu'B��zO�K[��'�4��q�n"���(1�L��w���FY��-���f{5��nx��%0\	ì�j�}FV�ɿ�"���9)腞.��o���%y��v���L������-�z��v{O��r��q<�� N�pMˇ�6k	}�����Nخ�������ͬ�rzn�<<�G{gzM��7��L��+�ᠣ ކB=-� ��G*��8�iqOhOg���|�_Y�1����"�x۔� �#�Y.��jϡ,�	���N���m)��3��!���|��)jD��r��_����5�f^��dB��(�
��3K�tD��L�>��1���AMG�]��	�"�W�������S��������vK$1���ݰQ��@FJ�󩤹!��Ȭ���o0蘛�$jg�ly>Y��i�梟��D]�dnT��"5�ݴ�}��� +��d<u�rL+e���&�[8�)v8M�U��vy�#�yi2�E����O�Ib񶟪v���-��>� ��՝�2��2İї�td)��0nB=�X����?x����m��Pu��Q�{S"!r���դht���#�v�}7�V�����eN�h��o�l��`qBc�JW˃&%Y��Yp>���#!Ɂ��+����ڠֳ�ԛ�6ÚP����c��v�B����bJ�o�/��W�r�����y��*٠�^i�LwY!�%�Zӏ�������\�v���q��.P�܈��9ʋ�s�Â�R�<qֹ��1ÀjD���&���!��A.�S�S!�,P�	S���P@sl��j<�sdM�5�v��h�8n��5/�id+ր��=v�3�=�g��r��Ш��ۨ�Ӂ �kS��Ek.1�E8�N���F/9 B�"�'Z��g��EC���`�i���Ht���R#6I���v�d�G������/pg���[���}� 1��ƿZ.���tk������'�hd�u��q*�n[Ҕ�=ÙB���ϣ�BS�]�UK).��t�F��{ݬB��^?o �����s`�XFpR'�:�9��Zn;�G�Q	ɪ�I�,)ɷ��h�r��8`q�wx|�t��g��Uk/�*0�Dlۤ'��'ހ�
7c�+3�V�k<R��$�OǶ������z��m��/���z?�W*g>����:çdm+���Y�`t����d�H��{A�9��g(�{
m��ËY�3���o��b�v�zTͰ�j6%V4j���[��u��+ɘ7�նCy�E�
��+��k�[{�{H��vݭU�/�M���)"��}�>MU��u#�s^5*��f+�@����ͻ  �����
O6��X�9��_�����֍[�i��'e�]�K��e3��7ςsVYcB��I�3����Q�B��}.r�a򕂪���ʞ|�����3Q��/����)[��Q�+xG�sA`{�}z!J%�T7&2�������e7��Β-��~��@�w�]��*�A̳X�/��
FyB����Y5��ToT��0����Lfw.��J���u��vE��~]"��� D|��u�A�T
\�^F��^&Ot	J=G:"�����!������>�ZR�e!��Ɖ�b^���U�5x�$�\{0[:a��_6��W_��E7��;�1aq<~�j�Aܻ�k�^��f�Z��wzۦ	�?G���͹��O �h�"�'��JSY1� ����r��&�g���WꇾS\Sl���A>~��|��{���/�aNFD���f�e`���$u��R�0����F��QG�wk��.����w�� ����Ԡ^��([m��x�?vuI���*��*�G�@�4�!��y�<'��&���v�HPFa�-�KZ7!��,��uo��l`��R��������m0N�8N7-�K�u�����K����J�=�pgMn\/rT*
'G's��6*$��#-jeD�;�]�]AS�}����2�Ьѿ6�j�R4݃zk��W�����pw��� �z����i�ҽ��+w�odDC��� ��C�7
y�5�zz�,�	���d��xc�y��4��J/�������p��~���i�m��p��vW}�B_���䜍�6�@f�T|����9y=���K�������s��pb���.���d$��s
2�E9@A��c|~��D�ub�o"��E{��`�Q
$�q�}�����wi���r-�ل	�Z4W�B��lჶ��Ӎ�a���4~�$�)�0Z+y?�mcG(	����F&�~�����[a���l�VN?Q��������㔔F�=�GH�K�-��o?@��Kb�~]�o�I��&Ǭ�ȷO��b�ǀD0�� t��q�����da�vE��D�c�B�@��/��6"@��	�o}��܎v3�	Z�bdE1�)ꪪ��>24��ƦHƠ����H��*Q�5\��3��}��@��r1O�aKȀ�>���^��_1���+���D��v�%׆u`�%Nf%�w��D3/'�Q��F�8�0?eů�$+/e��w�$e�a>��E�����3[�􅈋w�h��3�Xܸ
�Jx�{ǚ����ȂN���	3Aׯ��2O�:�����Zs�ܚCN�0�j\��0�;���Igk�[���#x�k ���0ۗ�Z�z��2�v�"�^����9K]v�[=�;Re�hc���h���'��+>���Kk] �t�=�x�STB����(�ޑ �����V�-		稢�ɥ��zX6��e�EsD�����ċ��e��ay6��J9\���c�(J�T��@��eR���/�0���2�~��m�DF�f�0�{���K@]�?s���%&X>�G�������̿�$��o>���ܧ@���=I��ǻ��*���_�>�ԡ��TD9W��Cx���Cda��v+��$��1����� �XO.�F�"��E-��3E�a��9�F�#�}�l,��
%����J����cf��_�'Ѽ�s�����~;�	����@p�~xu��]V^���u��[9�R�W=�ߤ<�dȪ��h����c��O����a���(�I
-z� ����%�ڗ�ߏ�{ &o/)�Ƈ$�M�Ǭy�q�H��/Kֶ�?�XφPO�L܍�0W�Gh
"j;T��gbe]@L��֟�O1���Ms�䝔eӸ=�v r �|.Z@`�z�f� 5�N�k�l�%��{R����@K9`6��X7]d1�.٫� �+`��5j�/a�%�^���x,�H���=M!�O����2=^fg������"ŔX1ǭ1�)%�HM<e�.6�6�ż����u�K����,�RG�(�k)d���q���g�
�1d�]q?��z�,�`f9����oޏA츶֋���Ac��LH�����U�����]�!I���}��S��yN*����}�R�h�nW�J#�NE�ƛ�a�&���bOB� ��,��+K��?���H�O��b�G��:K��"{�-{�����r5�� ��2��B*Jp=�a��Dmʻ �V���h��R\�x鎩ˋ=:�K�������=�+woQk�	4rߨj����s%Sx4i���tA�Ŧ�S�&����5P�q9T��o舱\l���*wg������P1���m|1I�#�!����e�O���5j���� �����gg��{��
�M����J���6/�B-d�͎�b TXx�mbY��Xx���lm�%��N濭3#y�2`���7��T��|I�l�l�h&c�F�$/�0���x{Э���H3�~XX��ZQ�ӊ����}i��Z�}���#��a���� �t��R�؋�vڍ�V�D0,Q 0GH��[�n�EL�۬x�v��M[ꢌ�u2�qի��l���$�&�r�^f	��ٿ���k�♝�]窏�<?��{�:K���:WK74�A��9U���\�!iDg_�ﱩ��R��In]����2 q�R8�-j@$���=r4���<9G�����ڦ�z���+굟TGؿ�Sz�ס��J5���Y�h�.�Ä�����<�j4 �f�!lz��-=�Z��0��c����������[ΚX:<�7��??���+$M�8�3�ʔ��2=��sk��]�qT�/+6Z_��^������Q#�M��>l����=�X#J�Z6)zoՃ	�}5#�-E	5�I��M��q��`@�N��[ě�h�Щ�Cw	C<��F�Q�N��0�l��&��I%���@ئ�Q$)�26�ZK=�{��!�ԉs� T�}1�m��n�S���GB\F��!�tg�el�n>���-Y��q���^�Yy�'��f�x#ח^UR����s������+ʹ�Y_l}X�H���A�_����3�D�[_�.�-I�?6L�%G�c��v�b�wnӖ�ۣ�Q��|���+P �ߧ9��q��Z=�S	�\]e�wI�>b25�,�m�g�Ԧ�WE�8W Y���VV:�*"�!?�zDŞ���1�/55��,H0��G��?M+�g�L�Hg!��`ن�,����}������F��b>:����Qx˨�ԉH�e�.bS�Ώǻ��#�%ݖ���o�Z���u��1e�q�������2��7�H��!Pvty=E�t~�$M�1�f>W����R�M���V(dH��@*p�O���W.͌��Ӡ�:�s(|�u�?A授�����*���i��	���3�'�3ނ����@΂Wi֮p䋺���[��%�i�Q�u�z���h7�Kd�~ߍ�z��r���A/�F⓷�
x���l#LykY����ٰ�\�[�C���1�	n��wPa�o��Ϸ?ґ5�G��6�+��L����W�P�;�mH��h������k}�t��[�C2��K�ѽ�����<����
Ѯ<kY���)���h��.�-+ya����G'g3�VB}��Ǯ�=�J�� cE%�f���ƛb�E��بG���_Ђj�4�Ӛ@����~v)��NV��aVzs]y�MNaDc1-L4��@X?��ɓ�n2e�� U���v^��:�4��*ݍ7���u�G�*x��И?�q�����ل�Y�{�7;��]&���t����W*�4�+ձ�Ȣ43\q�E��s��b�����@��a���'D3�oa�+�Ŭ�� �[�PV*��'�{�c�ۈ���tB��br����d�~�'�%�T��nQk(A� d�s�t�ը#��!̎�O���rwG�g:�:Y�����pl&�J��J��i�8=}�M(yߢ���Nz��Э�$46:�}g��7VJ݀<KKA9j�X�GA�CpX�mo�N�f�'R��C���|҇z5:U��A�n����
�� �%����	*6Ø�����g�t s�E6��I9]���ۿ��(�;�A{Ԋ6_�n<fg��_����mxj���Z�I�W��C�� �)cD���s�f��'��H-��� D�cs(��Ӻ��H+Q���X��K�f�|噽�#�e���� ��ޕ�{��IJ#]c'���ޒ���|ؿ7b��o�ja�q�9q��\�d=k�5��\��XA1C�*ǡ����dv��xCC9l�����'P7$����H�ʁ ��^d~5]�x~!Y���*hل+�4�����X�&Lh�D���."� �����fW�浩3���z�Cz�A�"�R h
l��7���)�_�Lff�(��_��)���H����Q쀷�,�Y ���u��QWW�en4\��Z:O��nW�)[��:R�YG��<�SEjT F-�rC���/��D�y(�vJ�o�RX�	<��k	T�K��\T;y	Y�9z(����L�E2��:�&�N[�J�Dѹ�`k���;�Gd��f�9B>~�"��� ��^�x	��29͑��v�_IG^���G���a9+Q��ZŢs���O�O#/�w
�����g�#�v��S��_�^#�	c����+�,ӻE���`����Hs�I�?`�C�R����݉���\"|͑��,^����HKл`A朗"��-�.|t�D�!�$|?xW�~�����5=lI��K�H�'��3�W�>�4U�i��=/X)c�X2�^&O���&xnI���\E[#�lڛ���{�Ì��,lmVUH����A����4�p�<W�c*s,��!��,��40>�6��?�,�n�.��_�V#59��%E/	Lj�?�G��$}x;��$6	�o�*�o7��~=��:f1hކ%�TR�i�k�Ò�`�g����+�gVr(@Ar'p��ji8MKz�]�'��t.3���c�<������-�7�b��ev��� Q5��j�Y!m�X�rf����U�\����`�V;���Xf���N���W����@|{�sM���o��� B�� ��#n@�)���/�v7�IHȌ���N�K$���ⵤL�|��2t=s�i���5S>v�Y�=�u�/?�˩���ʖ�.���
��ZM�
���P�𯱽� 6?:�����ě�� \��%)�u��S�����a�C��}��iw�!�j��9�2ܯT�U&]���-�uta@��vb7�b��W��~������+�mO��"���5}�L|�2r�aYv�������U~�0��As;w�ă5H�9������m�!ik��8�WZ����;(��e�b����u
m�s�����3�龞.|���S���a�7�WZw��2�����H;`�٩?0������(�GR�Y,��3/�y?�Kb!�x���]�7n�v��Ƅ$ܹ�.�t��f���w�v4po���\~�g7z�]��"g�.4%���ˌ��#s�5�y��1�}g;�U���#��|̋z��o�Zo-T[���e~������,> ��?�S�prqm�{G�}�������YӅ��{�X�����;+�5PP�q���9MoK��(�D�K��l�2�f~c��l���%*m0FH>�
8|�-�!�H�wፇ̛�d��#�Z�[~P�vx������u�ma��Po�#P��+$R�#�Z�"���5�Θ)<�@j�$aF^����ғ�,�g�h�����Kv��\�������ֺcÎ�m��u���4Ά�v�B�Lu*|��`�Bm��Luِ�
�<�����jz扸��#�-s�D1�0�:�#�]�_-o-�Ǥ��Ut�`��v��5@Uov������ }�$c��3�nle.���v&�	F�4��[߆��
�5yg���KQ���QA�a/`0Ƽ�@�f���N�W����bv�D�A���T�I��Μ�H�߶��� �Λ�{�ݏ�O)慴��%m%��.�a�Gޞ��X+bVｹQ�zA��� ���{N*L��l��u�/��|�8t���`D�5	^	GUf���s�Dܷ���F?��'ۅwCejI�o��/�W�/x���[s�Q� �����Ld.����.���U(I��c�MZ�����7�eF�������;�w�ߵ��yd�=���е���a7P����쎝ϩ��B&@O��y�h�/غK!�82-���;�\�Ձ!Ro�9���JJ����@x�>u�,/�>GHη��AF(oC���	�|���Z�pB�4��E֌S�-����UC��f���xLO��s�Q/�_\�&G������Z��ZV�����!1�>ꈞ;�*����B���0}KeqS���o�
�-����ED7���f7cU�Z�b�Y�Ԟ�%+�lyް�A}	��L� ��şO_�;�)�<�'@\"��C���F�E�����pb'������Tѕd��N��}���5k��ց8��X2����p����\
0=���ˍ�B^0Y�LJ.qRBHV�|C���C�N���)��Bn)}����F%-~�ˏ��F��&�� �K�W^V�4�s��eU���Iw�-�y�i�������}�vy�����Ta�C���x���'S�o���d��S���Dr��L������ςvu���#�l��sT��uz��q��`�[ڟ6e'�,ʚ�aw���y��z��/>$��ΘD۹m�M̈�iZD&��@#�8�BQIt0d�����SOXv+�a�o�����ibǰ��Ԫԇ�j���2/,�`Ra+c���yTHU�c*!�N�ᦡ�A��B�t��F�2��6��z<�Xdx �����o���>����(f�ub�e�����"x��$��2����Z�6f�ƨ�B-LFy�6��m���]i/�!rM�d�J�[�I0fC�@8�lUG����I9Y��L�W�I��:N�����ػ�n�O����v�+$�*�f���)fCw	� �:��jF���O_�/ľ�ۀ2(��q�l�Vn-{qeZA�Z~��[?V��^޴̱���A�bb��^�ڸPk�����D���/Km������V���z�P��gY��mg�)��
����rA�;�o�d�,��:��FO�l�~T	�$����l��
�HP�s�Wj}(��4$}��#(ۢ�ڶ�"L����Gf��j]�2��3p;L�t�}��w����6�%�R�8љL�(i�H
SN<�0x�@y�O�5� �t���ؿ�fy�����Xn$݁X�
�����dAy�! �|R!�m�YX�3���-;Ҭ�T�`|D����������Z"�o#3��TE ���101�\��x⺡%4��9:cݒ=L:��!+"}(.��Y��0�N���]���{�u�l�\%���EN�tڏ
�p!�ڿ4��Qf��3��g��'k2S���Vn?�/�e��s�r��(O˚,������Ӧ��+R�zR�� '��$B��T����a&��O��< ��v�Kr�5�@����0�"o����I�7��\�}6S2��]3n��Op҇~�Y.�_��-�y$~y��DWy���|f*�R�C��^�0��!�_~5=��v;5�e�m�J��;����;q+(���DզG�˴��h���6����������RW�;ĲdՔ�'x;��p�J��R�Xj^F�w`���NՏ�j��>E�kl�����8�O�NY�x	�R�ż�\%�ͨ��C\�$���[o3�D.�����e��/�|x���S**���kD��;@�/�K	�
[�l�G��F����x�:L@�𷓇��t�Dw �����I�������ZGN�	jh
b���O�yV��8
2�"���y׏�"|6Ƶ'Ղ��':$��y�$ �ݗ#a�����0PmdH�������D��q�|�ʘ ���2��g�ݵh��N�a���J�ɣ��`��F�Q9PYKm�<���Zg�d��t���
�`#r^��4��z��ɴ���F���o,��o�c�x��}yq*�����Z�UU���O+��W����+�8t�h�Yzi�׬,�/�-:-�p��S�[.�@�[;XA�Ȉ=������%^^���1K��68��t_$�n������^V����3�K���xz��1���� '�X\�.�j��.*�0i�[�i�V��;��)F�y���Ɯ�&���������(&�Y��da�:�6�]�@�&e�E�;���r�F�!!�Sau�MӥG��_L���O�{ "�4':p�; n����p�� ��"z��Z�8$"9��壯[��s�z�iD7��0�O�-cmĘ��}�B�"�����~�]Z��S֓�_ݱ:S�&�L*!�B�è,�/s�����f�M�H��8��ï��{����iz�0Z�Ƥ�a_∮s�=S��+�=���mc#�r�ٱFٷ�մI�|�O��&��"�
�-P�s_��W����ƾTc/�2��3:Ý�{+��L�.�5�0�aa�@o��Q��H�_o��G���r��x���kf��4#aZ	>���䆆�k�ewA�\�����7��.k+��*/+X�]G{�U�>iUt���l6��ʬ��*��i�8��\���,z^��eS맠q����G����~8�ф�O E���l�����֤YO���^a𻽡����6�v�Ԅ���"�$3K�3��Nh��H[!{��uC1���L�$�@>��F�<4��?��~��cc:�2����^��բE����0^9�Z��}#�c3L�lk�G�	b�`q���Y�a���_�|;k:ea��_<(ɖB�U3x:
�T{��Ҿ��8�&:��=fKe��<�^� ��SMe��{�B/�l�I��������kn��̨����ZOՁ�P���l��o�	1�W��T�j<`M]�[� �Pj�wڦg��Hb`�T`����9e$>5vq��O\�ij�]l�1ҹ�~:�b�g�c@�n�c 9츼'����#�q%�!�P��JE�ɜ��K��r�oꪓ2�X�"���L�U������~�ӓ_���A �T�T狧UA�M�p�j�?�p��'����T����-��أ�m��t�� ��ծ�EE=xj�2-�|@`k=��s�T���k�R5��p/��3G�J�'JH�g�8H���|�[�mfvݖ�a��N�]�ВQ2���8������kn�Jm�nc^�0���$���e�({���q+��%�:+:��)�F��\w�س7�"�y���� ]��3[�}+H�yb*����~�� X���
<��$�Hج@+�R�kɥi,�a�g+{_���?���v�!=���u��'����@'��!���1Ȋ󫐟������

u��0���$9D�!�԰1bm�s�d�}i��k�M�%�ӷ\����l/7� �o�x��J����S�U��Gk6�{g�(�7uV�[�>���� ��F��v�qoȺ�,�	Ϊ�_���)��d�}������2J�Ċ���.O��[�'��1�;L��8���B�ԗ`��i�"������'��I��ӂX</��Ag��Z%#�c���Cw}M�?�q�û�����p���x� �0|�l��^JA㷩4P��g-�0�|b�,��Ǫ��k��^? f
��^��v���%��.R�ˊ��+P�������w��@6���5�Ԍ0E6pu����3���A�w�������r3�,��#�����'��X2x�������~P'��u��8�4N�$?��1稐�.��@W}�39��$ݾ�Rj����M�\��z��Vã�2:� u"��ʳUE��?-#K���I��"�o���lMyu��Ge�/e�bׯ%v�˩�&�Ҍ4�X�<3�:ki ���)�刾j����{)�w�98.�9��#SV:^u��"d� ��d�Ԯ����?�E���c^&��DC��4�jf�-v[4!��߈&v$7�[��v�?�ݲ<sc�ح��Z�bʃ���5��8�Q�d6��D�E|Ѩf��y�X�'P�y���n�O��D���f���5�ۅ2��iK(�ʔT�M���.[+±�a~��ہ�ڊ��=ao�=Ε�f���e$����2|w������INƶ^��tH;UgG��q��/��2.!�q	N���H���i��J��v�f��U���aZ��	�؊P��"�]W۱��<�_��>G�0�ӫ��n�k��K����P�ō覚^�O�D��n���4ĸ�^;�DU�����^b.|��V�ɯ$h�?��֯��R�'u�X�J,쾸�P�p"���{9�i.����҆�ҽ	6,�5Q+?1�yLu�E�Ѡ���,
".����ߐ���-:��`��Xjv���t�|��tp܊P$I�l8���:�L��3n�W����l�G�q�x�ع�
�s�Q���)�ڙ��U�	���7t�N�&t��)N����%.' _m�ň���d�J/\j�ݡx.S���I�6���0E���^-i]����ԯ�)�L9	[��lLoLj��:!�5WO��� �7=U�tX�v7�|l��1�XJ�2���ͯ���FL_�O����Xi�gƗ}X7�� as�F�Ǌ�����2�n����M1K,�o�!{y̍be����� ��48�M<=�A��Cu2����U�����Ap/�wrQ���i�c�s���⅏~v�P<�R�f|�%��[i��ZHXaw	�A��DV��|��ݑ&���1<�yX����O�z�)W����_T�g!�;��M1�h�P-��Fe�/䟯sR�����*�����@!�Ft�(4�$�O�'b��[��G5w��OK�/���N�/3-��)��Qt���M�x7=5=��E����X~r=��0��	�hUp�"��)��>!���]g�5}U�%TPc��M�܊����i�L�/�k�.̅�i�c�r�w?r6��S�	�~�茶����*-JK�F5����Q�q�MY��
":���]Y$Mb��)ځ�'XSe�϶���/D%r�!�C�-SX���D*��6�dk��u��U���D)��/�I��2�	��3�B�Z?I��\ّ��KL�6���r�j�f�>�~׏�������S]���~�#�$
5xLVE傦�ۈ��.3#O@��O��û�. K��Ngd]�:f�ThTl_V �1W�=>�ۆ���cMr ���=:��WC�9�vvk�ƚ�/��#�
+y��cޓ���Y+���!rq0�-p�r��E�w"5O!~��|�|.��o�>$���ӢP*�Ɓ_��1���lp௺��F�Z {U�S�-�w�5��� _�����]Oy'����y��v��}��=��Qu_Pn�Ǫ`��(���<򦉛"	r8B�4jFM�����e"���Dw��%�����>'4��	���n��!$�HΈ�]�c�I����	��T
���V)�5?g�Pԉ���"�8K�w���IN���Hڻ�%�
���a��<�z%tЄ'�1s$4Y\��cRr��#�.�4��1o�:�vkRWUv�3�X�!�`p#ݼ�J[�l�Hf.R�\p���X���� ��6$����Y�֐�����ɛ̮Z�LbQ5�b�{��\M;��}�|-k��ؒ�:�Ϻ,1���k����7S���Z��<��<�l�=I���3�ƧX�r��X4Nc��JQF��蜥 #�A��a�F�V �{�6���$6�Y��O�s���5b`�9���}�cC����r�dBצ6U�< L�&1Pv.��R��A�Ҁ�c�q�W1�;����鰖/�&-+j����		�v�!�w9b]"~��1!(0��v*����[ÞKs(Ui�w�Y^j�Ƅ�����7�q'�]�/���H�~���"#�/7������	�-�%�k.�z�4�|V�h�*�g%Z 1�e��ڦ��D��v���1&L$���vu�8��c^��;J�_Fdq""!�2z�Z���Q��LUI�U�`��R�2�	 /Ḋ%��Z�M���.2it-��f�4�c����q��D#�*�����)FSR�:1�}�#plKB#�Z->P�41��x0���Y�U�½A����ʖqR�kRzģk�pE=��hn`��i{̥ǠS�*h_�]�$bsS�7�Y�k?�h��$��&]�\v�x�ͼ�O�cSc)�]�����4�o���੆q_���<@q��f�5�s���ID�ܚe�1��"Ⰵ
6���[u���e�#ǁ�*�e��[1�@����̒�Ԁ
�V�i}�OE뼹-Ր$ϸf��f'��\����S�T�?W{ F}��+��y��_��'f/Ȱ������u6I�?���i�Blx5���裇3����I��m�x�6��a+t&��T'�~Jd1���J�~ݯ����p��畡��`�5��8��
;�Lf�=^?U �uC怯��t�+���j�y����|G��(���V\���d�o���V�m_���OM�ZX)��yj�
�p��W�]}.[V��z7���%+P<Jz��su�Qy �ΣJ����-���'������G�`���g��u�[b��F7sH�f!t��O��OЭ;e���㫡����!�E�>�o�?��t��n��fj��?Ua`\둮��ا?X�e�l�&s8S��ԡv�^*je�4x�x���b6z��g���-��M����5����G�����E=ݤ�5��XY.��g/i�ɏ��t~�Y8E.���b�P�0A#q�A�ﲹ�_ъy؛dq3)Z`�0l2�P�Wn�I #��.�{�mKJ�t������H�IT����V~��p���O�'�_�P��u)0lyh�k�?y�s�1������Z���2��;O���s�VQT�Rv���g}Qeq�����N[���n���©���1�����gn?�kN@%�M�f/J	���F���P�/@�<8ϊ�ĉQ\ `�u���Vv_�"v�w_�{Y|}��`}J�����F�	|X�Blǜ4��,y�������P�hnx�bۍ���(^`!��f1.Uy�+*9�C�E�� ;2
��=�rP\�Kh���o?��yO�
f<ج"�s�G��!1i�0�;�t@ {ұV�K�2'�kş�A�EG~��rIry:z�m���%��Pv���o&;�p����z虃Z��o�n�+�³���@¨3�K��}��E���BU��n%�M��&�����uD&
?�A���-�̆�M�YiFz����/���V?i��!3��	���ր�=.\U���D�p�yw�.
�ã�Yv�h
o�{T��r�^�Ѥ�Gt(���n̛ZS�����q�U���bK��Ux�k������یu+L��:�RΉ�<�r�~)�	�� g/��.^Sa���)���N�����W\��w�k�Yy�[���921m?GxѕQ�'�Hb�.j?S� ��p��P��A0�-�z-L�ߨ��ՕX`�0���� �J���	4]���������5@�u?��r�D��%��Įҥ|e�@,\rGTk���q!��=t�I4Tr�A����5� =�'�(���R�
����0D�p��#/��m��#tN�pW�br�@Y��9���`�_ȹ͂���`��kS�o��Qb�_��A�N�3hNB}Ƞ\s}H|�;�3�I�����[A+V��=��M6WZ#�<Sϻe"�mo�=ab� ����g5��V�5R�/��)�M�s\�`�%e�)��a��!�2v���{-nf :`�����	�>����� })���g�E�߽�)>�&'��T�n��Y�RE�x)��S
�|OR�.qڅѲC��8㩚��m���v"F�*��}�t,*�1���pg���`Hy}���a�Dk��٪)�8���nM�ŠD�b��;^�l6ʮ��,T�8Bڽ@��@�����[�}� ����)~X�k�m�|A��$���!�`��	E�+�탐�L^���uy�D�x�@7߽gT��\c�_���J~��e[<�YO�kt�\D�!}�s��L$nCrֱ3�ym({[�pK�M���#���=J>8-BhJR[�X�g��34�LRj��BH��]u1��u<v�g�*�w�Y���N�P�_K��˘�rLU�>�Ы}�6{joUp����"��}B��ivE�Ŀ��g��zg�с�P<�)����F|����P_NB�A�X�l!v��n��fI��[�dli�Z�z辱C9����r2�]�<8;��`0����Ei�{�ҩ�M%c����r�2����^���넞F�*>5��0$��� �F/�0,K�)E~���w����1+/�S���DE��{?���Jg������`�!��&��b�p����!�ۣm��3�Ns>��o�u)�{?h�g$�]��y��s��|�b��`�
���*!S�&�VG������S۴�Rs�;W��l���Ҭ|R�@���A(_#��;�ez"�[���b{-��.,z-C��(���\�*�����^��'{!���	_��֮�4����}� H���.k��͢��@��,�9���D�jq�S��Q@}F��H2S=� _B�!��؈�:D�.?����NQ;S���e1B��6�����Y`?��P*?i�a��b�tj?"�P-�����GhY�a��"��~��+���2�����.Y����.��c�#�X;*����FoS��U�Wc
ZR���Wl� f�eI�8��4w��L�f�*]��2CM�)L�O�,�%V���3�����n�V`D�~8?б`F9���t����ԓh���_��":Bz0����]�/;��0.�g �
��ޑ�(��َ����B,�COB��Mp�����[��a�d�"��E�R��^�U�ue+"�Vc[2(jF�w���%|��[�,�Au�^��sߺ3<����@��A����_,�NY ��zs��5�!O���OP$Pj��ŵW#>��!��<Z�1�� s���r�s�@v6�N�Q�4�ߡy4���UĪ���/��TX����Y4�``�2l������c���o���&6U��l�">n�\W�%w��<�/\Ń��C�d�z~>��
�(��10\l�O�ƨ΂��=T=�����[���*�0���)����[+X϶�9_�k����jY0����-�;�!�S�V��'��_`�5.m����f�Rt��	�{��i�j�$�nr�z-fa�Ui���w?LR-��m䬦�S�j/T<�z8�?g�TMN<�]gD����o��(�Q� h�U���g��d��Y���HO�F�r�}l�Pv�y�>=t��grϴ�TCK�vNb�E�H��7_�J�u�-v����Ϫ�+�ۂ������N�D��i(��9��/m�7[�6�K��z ea���x��*�
�X	��?XU�~�b|Gh����S��2ȋg�8�J����?A��<�� V�<�DJ�Lf�������jW��@	팱_���Z�H+�
�q�BZ�, K{:O�*��/���v�I�I�9�G�`ϗ�]�Ki��9��ǣ��l3sҘ�LU�`Pj�<�N��E���߫�W`K3���Ld�慺�EX O0�ݕ�h�XJ��L�D$�6��3�?Q�v����S[��t�p$�X�e����ᘡC`+��[�7�1,!�*l����s�� �DS�E�\�%��ݲl�Y���*�2o����BE�X��)�~ؗ	�hs>�Rf\3��0�FK�z�~�GhG�6>Wn�M�����8�u��b�{]�*Y2dѪ�������g�z���X���#���拉�I�M�o��,�]�8L�<q�o�}݁ҫ0���F*V�l&QA�$�Np`�i��N�aX}N֊T��*Ji��uʒ:r� 3���npxYhF�����B��ڽ@}���[x�_��x�Mtw�w~��
�/ �qv�6��G�`(�)i�2б�e#$A�)f�]��� �Q���0�nR_T1^?V�[K�r�5+�Ռ���p���>�V � '�E�	b�`��1,Y�^�#�����HPMV����[�Yvȿʭs.ݝ���!����z)
)���ܯ=��Y��3w)�l�%0����!��nxA"�Z΋_ojt}Q�N�] ��o���X��;MN\�;H�~��9i%��}+��j�i�U=cM<!oD�RsO5�o�W�Hw�m
�̚n��3�+���[���h�����	;�DV
^c����OW�2���jů�I�&�S��98I�����%%�|�
Ò���#��*v�y���.E;̎�Y哧{��)1����U���T�q<�^{������.Z�����>����ܹY/������O''`j��y����f�;��_�9u|�s��,�Y4U|f;V�����ͻ�����o����!�ha�Ͷ�����+�b���_L�&��y���a�%v�W�(8p�_S�~�0�bE��9&��kV0��g9�ƚ�����0ܙ�I#����³��C�b�a67���b�z�Ӭ��k�L�i2Ms/D�	
ҹ,k6�,�(�!�y	3��Ѐj@���9�u�]���%M����-h��Ŭ	A��Ze-F��^�P�m7h�mz��J1r�u�r,��vbM�S�5��u��y^���%PT���C �!5k� �r��ߋ�cr��S�%鿝U����)bS�&�3|]�֡�NB�]\�ia��a���Z:����N����36ukr�n�����P�ba6��
F�ߙ����\�-�g�a���ߣ�	�P�E�����QFR�T�;4���?���YⅯS���Q��m��b�����Bdc#>*/�8�g�,iD����=_m�;�W\��7A��ƨ(\e�A�z�[t5��֛b;�'���f�pk���Vw�s&I&U0���q��hC�ڈ��"�'�w�v���kv���=#޷]!$:Z�O+a�lc�7k7���ߺ�4j�\k�s�D@�5�yM��ؚ�p���.v�u59��B�i�����	��n!)��-oޚ�~:��L8ނ��Ҝ����Z*����"�q�)���2�.� �p�`�s J��­�Y�����Ŷ�����C�gN�"H#��@�zw���'ZOB��[�@�أ� ��fSCA��YbnF�:G#h��흺�,,��p�"�cj؊�y����rgÚ����rr���h���)3a�=�.���iW7�����4�� �c �Ž�)�ߝx��wP����X��BDQ&�%s���7��6Y/
ꍿ=�[�?��C�_�1Kk���#Z	��T�C:�ש���A�Hm�8��I�NL;3�d������Ц����� ٝ����n!�+�S��J�MHM����N2(İ���a��o�0ɼ-����6�9��@~�)�p=9N�MvY�.%B^qɲ=�;˟2�*�cѿz�'c��;m�{�pFhO�Qo��Vj��-:�ј��ك1$>R��*|�Q&���Ε�H���ߞ�5 ?G,�]��j�2��s�.*���Jde��cx��e�N��pߛ� �b�����8�vį�`q�~`:UnuHoB�Z<6b�a����Iz��]��13�k�)�8���y\����i�͍�H�e�J�n�ͷYJ�K+�F l�jZ�H���a�&�'L�GE���d��'����!TH'8����E���%\�� ��qV�hǲ?�lE%k˱e�$��YU����=����6qe�3$���jI��Wɚ��x��3w�i�م*�v�����4l��Όszވ��j�-�TG+�4y�(�YmN'�hr|% �\�4��,�Hu׍vH�C>5i��E/�^�X�芜��X}4$�d�IAk_�P�|��V"귚�sy�Ѕ����ڭ�}����{����FА_��yrz��@s������Q
A�W��6�/wL��hϛ��"���������)��L�L-$�{bA��F���Y žV��,4>���P�Uo
?.k�T�ۉ�j,�\�~��\azJxu:��<�_���Y���{]C�ᛉ�6mYj$�>��8�H�X����&=�z�i����sHMؖ+$�ժ��&�$��\>���a$�ʳ���wJP��(t�h�'�O-����ǝ���T f��H�b��ueK�k%v)�kwm����K��(��ʲ��a��8��46�Xd6�yc�h}��b:0ku_�������}�Ɠ���yٽf(�P���H���sn��'���OybU%�|}���O���._�& ��%�0>셄�Ts��)�\�� ��uR��d�!"���&h��#ꆐ̐�Lm��N����?<�W���r򺋀A^�?�UN^�*Jj�D���LYе�6Ї���Nt�����`n���2�CU}�{t�d�%LeK�'I�����Ң��,�+M��� >�c'��qnqL��@�Ġ@����ӏ�n�cj�Ԩ��&���ߔ��{����8��?�4��\P��P<��͙�a��>:G�x,�}�s�KƬ ?�xx�l�)�JF��e`���� Zs�g�`'$���7k�%
��O�����?�,L��J�j�;�֞S���cD~�,qܦO�c�R1h�I	�ΆA�_�?�|y�n�ة�m��GX��,+�%yHE�k�g��]�k ��>W�g�����%���rqB������o�#^!�_����ʩi8����4��cw�����6��������S�f��i�ʸȢ� ��S鬈�#�&������S�$_	7vZ���7��*TbY���-ť��7�B ����Ni�����ѪZ���,�~v�q���˚��c�����'K�9m[`�n�[�3�����t��nZ�6뙒�����h�| �rWwϿ�ʒ1g��	����	���o:�-x-5-��T:�5�H���6)f�Α�,^�J�}�&ml=^{z�H��0@1��Ϋ�n��0����j�k`�Ȑ	�r[o��zN�ƒμ;����iJv�Fm�|��J�x)��ԩZ�h����!�S��M��ܳo)m������yWa�!���4s NL�]\�$�V}���N���k^"e2)�'J�_hn��H}�k��j��x�!�7���� ���L�7$wk���q؀�
��5|�&
n��ȇMx�u�j�Y� ؈���5�����^Rz���~�-���F3"��:�9�xqTڙ�7���X<R^G_p8վ.�Y�&������g5ěE=��BzN}��x8kG��� FLa����-�&=�(�oX���-�$��&�v�&�G��{�tţ�����+��c-`�- :���?�����"�q1Ɏ�,���[D�a���$W��:n��.�yV/�d�wSZ�B-:Y9�.��%���L���9}�/�[�YI *����!�qgY���F�E��n�E�-�er���o�B 7��'�ؾ?ܻ1��,I8���ٸ�����=�dDKhK�7T�I������p�$=Xv8�w��M3�VQ��41������=b'���J	��9��+�YKl{���*)��u���Ӕ1�F8,3���Fc�5I��hM��uL��&.DEz��L9�G�gᩋ�4���|�/�_�q[���`�Q���A`�B
l�A���Xw~4фY�R�)��G����k%��=�0[�Os�>P��Z%V|\��ףkL*�}�5f��5WsͿ��nR���6����a���ˈ�M����4�C�V`|N��,���ьS�5Z\vfݝ�(u���P�(�H�s�/�w��o��ʸ�"q�Xzkhh�)~)g5$�y�=uԠ�D� ��PW����!�{��P���fǀp���'JK�gA"�%���<�m,�L���=3�gx�}�H|nx}�p��1���Lآj��Ha�uh%F]�z����?������W��c"�@���I���=1QHX�'�{�ޏ�W�Y��K(E�y���#�34[���c�g�?<Z_3f�>z��~�E���0Py�Y3�o]���2�K�lzh�T���4�����;2m���D�
@^=Ѷ^,E��i����U�ϓ"ă[0-Tu8K������B@����oQ�dm�Z�N�����D_�3�a:>��Y��=���eSvDt�O`<��`"3��It��Is��N�� e�9�!@�����ٚh�R������t�l>O��H���9��='��?K^�Kv�*���`��P45�d}"pZ�4!j0��R�7*Zq����ج��v*��~B�@<b*�d�8��K����׳�&��.���ܫ%�8�ӹ�[��Lfu}��8�%AG���U��(4��zP �ײxcL-�!�����Cޮ�,�5�\�k�;k���k�g�5����
5+���m����KG&f�W�*���gm4Ð��=9Lc��^���~w��-vV��`�2
|2`��ic��"��و,g�^��F	��4�6��2�p�P$�C��S�I��f��)#JD�/��}~�$��L��B��Ɨ7��5�+��
���'��[���Y_cT鴝d��i����sU-I(�j����)����Z<���$«L�`��{���B��-���B�w��XD���3-S���Ѣ,�\���ղ
�Ve\��" ��$-�ۯ�wۼ��I�[���1���P[?6QZs5uv�A����UHז.zaN�D�J��XM獧�,��f8XNC���'�7���P�\-ĶI��ُ�\��qZ��i�@��^z��9�A�&���nA��ʵ��03/��QD&{k��]���'�p�!�6?��ut|���Vh@E(�	�����0�K۪��0��2]�3z�C��#4��9>y�t����Fg9�oÿ�Z�m>���&�u3�>wB�?l�r���ܒ��`5��J�2=��Tu��+!52="/��q"���\U��GF�f.A{c��D0b0��9��ÿ��P�>�̵��=d6?&�����*�0�hO}]���,��3qb^�~����9�
������c<����R%���}��ǳ	���q b�m���w�hP}Ȇ%�\"�Ǔ�("�Hg]�Ӷ�@������w���Mɩ��C��;�`
������<�܁G���Q �`͌g��3�pn�F��w��d�zI\ޯ����a�i�I溯�(������5�|�Y魽�y篎�j�sZ>��C�A�*��XG���#$�ò(i8�z!z��98:3�w�Kʡi�
��h
���`f���Rӑ���[	��)*�}�$�~#9�ŵu�8��y��;�Ƃcej�8�P d��ԒtA4��H��g2��[%A��Y�Q�T�����=�Ӣ&�8�Y4�3�ҽ�qkQ��N�ُ<�֡���83X/5uWI���SI�s��!:���1*8C�*8�λ�������lXY��j��~@T��Iy������坖TK'.��bo뒫��^��Kz�@���A�rc��;WB���Bh�;�l�0�fJQ���4M���@ҵy%���z����Uyf��z-S�Qc�b\�	�7u(�0e:��Y������s\Ċf��.E�����z�O[��VYv�{wzd����of¾��4�;�B���p�����a��	��%5�Z�&�ۏ�%�D��' U�\�ظF�����8T���&-��QO��w�u�T*?��V�D=c�r��c��#�~���h�k͜�PKw�P�ߜ[cъ^{6M(kR��_�N�H4�>��pK�Y��VpYS3�agi]\e�R�~�� ��¾�V9RI�/��Aﶦ!�k����Q��� �6�A��[a�
�:����◛�즦<�b�f�!��3*
 �U&*C͈��#��$Y�b����Br� N~�]��0� �»{B�� w��d<���.Oɾ)�� ���/�ri�4���u5\Քi�»[ܥXZ���{ �%�ؚ\z-�9k0\�_��3qM���M��~�傠x+{~��c����d���L��@�5ep��4YgA�x$yPVF��*�݌^��E��ן���x�~x,�;�.�J�D>`�,�J4���urA���$1��Mh��T���2n����{��Y��E��!�&�ӝ� ҫ&sPփ��C�a�� ���3��e�*F��v��p!ܹrɚ��$��
v̠�[�G���:#!����o;�J5"�v�� ��X!��X/�Q�*��W	yi�_}&5�@�,�MWc�z�=���,��kׯ8^��nԬ���錕�ie@s/T��/���k�Iq��f>g��ɛ�Y�@��	T
}%��`�N
���q�POw���~L�b�ZD�_k��*�|�߫.`���Qښ�x;���Z��Ra&�ڬ� N�$�������r5L�>1yU������f&���?�{���'�F0@)�S���s�^Q^��T$l�6�"i���ri��`o�b��e:1S~#����������FH#�#[F3b/ p�r�d���)�WсAUp��2u���f�b;�T��ј����
B���;��y�Ͱ�(�����0's����@��:a�<���`���0��M��i�ChD����p�����3��Y��v�g~���
��Ǳ��}y]<ܘ��5�ͬ�X��`����M�\C%"�y SQ��63i��A��Ӡ6N�d�#h��]�� �3Ut�=������O4��Cw�GH�HS�����S�N%3#�����]�`ƚ�ъ���§�I�N�}���# 3�&�a�r���s��$dfN�^dk��2�+�-���h�iiua�O�����rҲA�߃VB�V�:��׵�JGC����'U�ҌM�R��f���n��ne4��|���Z�����d&���k�F�RF�(Za��q��S�0��rMG�@\�����v���m�3�L��J��Y�Z5��+�a"D�����mܳ��~_��4��$3ƿSV��@�Oox���q�������OX�����TI]+�����GJ!���4�X�S��j��@��;���(ak��{���⏉IW'�ݹ��$9����Y.�u���P�z�.�w�4t�!���L/W6>���y�߆�j0��|A}tٛ����c�?L��	D�	{Tۛ���΁k�XC��CX�a�ֻ�+�	��,����~1]�#����ywY�rIn��O_��m��u�6���^f�G��Is����dv X(7�ߣ���E���D�J��D�4;�![�0�`�p�cK��T�c����]�(:���0�c���S�<w�R�iQ�L�����J�[9�D�ֈs�p DU��jޘK������M��M17�A�xr~סn��i$ʲMCS����hhxn�V�0Єn��k8�&�o:����b�i�n1���i��Y�+��0�2�g�ĺq0sˣ��(��4�%_���I<�C����%I��<|�f�-�P�+5�V�@ f�|��� S#������{���A�u�G�����@� ���b���x��`n���*�7����\�9L�Y
������N��������K������������Ho��i��p��$��{�T���&�@J.���a�l�Aڏ�{�^�|�����~��ѩ�2(����u])���HEY���Ɏ�D2��:4��d\�4��/a�k.\�:WŤ�"�85���斉Ԧڜ�J�T�;q�sX�H�bq�s��ɩ��Y�y���r]M��v!y���۾D &O��H����h�ZJ��Σr�QՄy���yp]2Ʀ�٤�"�2iy��]�*��o>"6L�^%co�{-$��+�bs�:���wD�u��uy���G�#P���Ŋ����d�Auv��_��� �_�r��8m
�
��j�I�<*��~ý��
<�u�&r�ؒ>a5�J-ں�c�+�*�7���d.S-rƙz��C�c��f���J����)@��8^�L-<x7�Ȏ����L��T3��85�]J�J�a��Eamh��"􀄚.8LKhȩ�
+�iN��Y�gY=�R����6���Q�� alj��iDIU�o��?�jM>oJi�=P�6��ݑ���4��V<꽛�V�p��G����_�ߌ��6�Q����x(��1�39@�z��uZ��F�lD����� �ӰB��\Ƽ����|��`T�|��?:l���������J&�
�N�H���T�EzrK�y׏*�x����a��S�f ����厬�~C����=��Ak
bY�T�����D��
��Zo�9�~�a���a8*�G>���f�b�m=�����P2k督zn���ߝ��a��vշ��0"#��t�/C G0	�^�?��Z�9aqS�&��{Ɂ�B�q?(�V=%j{��l0����������t����Cӯ���9D�#r�:z��7m	u�u��i�^���wX��Hl��ƿľ����"�}��	��QN ��猄
 ��=)��4.�(/ͭ#�P�G�r <���Л�w���"~hd�CE������1#��a;������.%�Y��,����p��>�h��銦<��!�״�s+�)��/I+"^�	����Sh�W@'tnJ�YLJ9�S���q�'S�z��h�r��;��!'�k)����3�~�E�Q�G�:!���Մ������{�E9�Vx�_�q�p�2:!I|r����pX9��Ќ<)��ɘ�r=c��?�gz�
E@`�[9��/��@/���@�<	���8��su�� ���ԗ��_����� �Ǔq@�1HJ>�&L~1B�"��uii�*� ×��>�J�APj���r`�K�_r������h�M�:&4���o�)0�Q{gHc��zU]}�_�6j
4%}���a�H�0��(��E��F�^�1�U�U��b�s܊,L%_5�dv���l1W�a�&{I��S��
1	 bS���na��m34�󬗶�L�h���J��`.����7�}0���Ɵ��
�=���&p\a?7
��R�����lk�^���i�J*e"-��^M��D�c���HH�� y�&:�e�^إ�W���y���:u�PÅ,ƈ�<����=���͸gO)hHX�g�u�]�Z۟s�q�¯0�����f`��ګ㚬 `_q��L�sO����L4R�^IQ����n���r�b�P�����
���Il��λ�L[r.S����������ݹ�%ݿ8�̻+	�[����|Yi�=uf1�{Vח�K����>�z����,�9Ӿ���d|q�$�5�Y�/��ۨ�=��B����M�q��ۚ�E꼸̆�-�Z;y�bm���X�����
ۉ��&|�P���*5H�'N��7��݁l?ħyzq���k�m�Y�P S��M�=� k������2e����n�|?�۷LȻ��ߋ� <4$j!�D#�Z8����E:�[žKW�@�D��E^�z�JBVq����SeM��x��AlZ�ZI_��2Cl=�D��{W<cc�J�7HB�(_ ��X�G������:~��~��h�V!l��$X��3} �����VA�b[�Z���b�Ok���� l�XIJ�Io�sw|�+�N{��%p�3���fDR�w��b��z�
�3*M�1��2}^s�b<���� �ާ�Ԣ[ ��=7����Qb��S!�~���f��F�-���߳�������Z��u�BΊ�nx�]��]�3	�W)�$U�	�'�Aߵ�s� Ï�v��?�7�)�z0H�9|K�%�B;E!������m0���+�#;��Ղ&��W�"�������
��y���o:���
T5Δ�&.�'��LW�i�O]�qۉ�fS�_?�[�4�ď�'Q�u}�ߵ��ܫ䐔y�R���(�^�J�B�tk`n�k�����RM��Yz�ЪH�2-���e%��sO��������z�l���=(eu�N�5�&	���:� �A>��ċ�qG��������q:5�aQW鿭����\���r��oj�g�v�Kt�M������$��E�0V��	��/��e�7Dmh��O��7��`QO6���#nx_&�I�wΜ��3�/��;����qot�ez�x2-�&���� a�Ԣ��Ҽ�Y���3&��/���ڷm#Z�sI��>�i|�͏�GD'@�}����2w�a`t�<�D��AQ=���̓@Ȕحn?�DϽ�i�nlBv��;��5H-F|�.�TY|��g~P%�3h-M������=�K���Ti�8�� ��L�oI�956�rwa�ή����1&�QQ��ş�$�?���Cm��eƧ���A�����=�������yg���ˏ{y�]VG�n�
���//Dߠ�E8�k�U����n]_>�Š��o�d:�QM_j4-���@-�W�)_逸���	VE�j��[�>̐*�pdd.�-Q.�gg60bк`�Ts�|�o˝j@G_�Jf�!���<���2��ěvt���ȫ��e��k`�׳��7}Vw�X}y��;�uU���婿��m�}�3��o�os,k�勚���%(�V:�� ��c����Z�9��r:vxfW���TT�P����|����7`:���r�?]�i������c�i)!"4B5�d��&�z�\��yz�Q-?�����0��rmx��n���l+nL`�~� !���M`|��<�Y��2
ۀ:Ӭ��E�4��
^㲌�(�J�la�_�8ǅ&l���Lt��U��Mz�ߍE]yM��!Kf�a̽��s�x��3�V|R����8���|�r�yb�;���#E�� �D��|�ٌ
.�oZ���o��b�l�`C��Ji��BX�*�=YN�W��gdW�� �=&�yw��d,�.ZxGh�[�s���q�MPoU|�O��
v�BC����hi���$Z}|��	���I�#�&�FC�}J����������5	����]��_& ��c�P��xS�;k����M�u6���L��p"������Ɯ������Na��6GΏi��PD5���P?�����Fp)�6�I�)��Be'�M#B�룔=�q�D�iGr'BbB��~A��R�$�Iʕ�wBMhȝ�[�L7���y@�7`�d�X�XٞڮPHS!�C�eiۊ9����p����;-T�df���G�G�Rܸ�E� .��I�hL����mճ\%;�W���?7�䬱 ��6%?�}����/P��	�F$e۝��yy���5D�l�<O�lNVG�F���mm`�]�!����]Bۧ��5y0g`=K�X�l�bxo��_dt��2e[h�Gs��}�
1+j��-��D?$`i�Xxui/'���u��0 �n�\R��&&��{�t�����,E�_��8B��U$^�S7-�"�k0KU��RS�T�qt�=|���}�P�A4��G����ka�OfFI�66���4�/@��"�ݶwN�7v��;��'��q�b�&8�S>�.�L�ѣ��dC�������R
W;�,��"tY�r�<}b�Lg?G���H�۳}�����tëv�C���2�oq�c��&�ql�u9ӈ��o/r�dSð�`=Q���">����޷��R��Y:n94aq��FI��Y�~��p
e�^��L�|��/vW��e�]LcS�_#�>;!q�d-%�mAC�?:9y*��L�j�P�i"y��8����!DiO�&�Ѷ�����ż$j��;���X�f��0x� ��5ɻ�;��e?�˦a��~�+�� �/NA��A�*3J���;|t`��ق�<�S,~�����������RV�u�N���w̰0�˸UQ���ql��X�iz��H�B�Y7x���J�B"5eZ�e6�%pr���z�ZS.AR�5i֕��z�1#�a��ѫ]���57�(��ә6�>���>A�oe+'E�<%�`�����<�`��X�G��l� �yMԻ�}��1���l`5Q�(���1����7�3�O�'�_���z�ҿ�����+_�[ �ʏ�	���lD@TN�6cT�<�lO>��ۏ<ĂyJ��.x�/p��^R�ڣ�\��0�A��/	ߣ*D�=s_i�kٯϏ9r�8��H%����hi�3"����ۤUAK�G���y:�	�J�x��Tf�B"�X�肉��'����H�/p3Df�LW��ד�~_E.�E|+��C+�7��8����$赦��Z�KQ��6�2������Qs.Ȓ6��:B���:�U����1��u���ap\�@�,(��=-�kv�h^B��B+Cc22�n&�$�B�q�.`�/k�NI$ɽ���-��	@7�vĆ�b("�X*ux��e����4��2��8q�k��/��mu�e��r�5z �{;]�0�]��}˵}m���~�����>�<�*D�&�	C4��o�'l��#%C��,�9�7"J�!Zjϴ]��0@WIk%�u����M'$8l�D%t��Ʌx�����}�/�h7Щ
�
��<-�M�j+�l�|)�p���Û M�%M����A���=d.�~��M��N��t����ot��:iB�� ǫ��kL碡!?�h�|e������8�bG���(�I=Sv��/��+��moA<��fKx�{�����.��y�< �a�{&xI���l��&'mnzGPn��~�~��@k7��Ң�����.`�i�g��NW�|ɉ�1���M�����6�8������P�,j�f#���z�9乡��gZ`���D;+��h$#r��h�C��Y�n�F��Z�Y�-��w�!~��*d�S�@4��z
:-��v �p9��˪�ĀNݒhW�q�-{p�
_�(�3?)V�zr8g_�Gio�vK�&ڢ�|?S*�6�^�/��z����f��Z ��w�
��`.�3����� ի:H{��z��4[�W�E��5RR��6�+�z��j3���SȁmT�d=%C����>i��h��m"����x�-����r�|7!����U>:��Ÿ|d��u:.^���GU�U�e���^��C�w�1DZ�+Q�������z���w������r}���d���^�`R�����H4�ZJ�Bŏ�!����e�X�S��+� Hz��Ape����#�րd!W�fR�Q}3��*����bc"	�-ۢ��t|t�u.��'��ܾw#������F�?z�
u����
	?���U;��u�uJ���	��ԝ']�=�>dG'{�WOkB��;��wY̅�#e��@K�|���v#��������<2�.A7�c���cHTV �mn�� �m���d"�u9BK�.�U�(?�Nβ�i�u�2u�&"�-�[���{dgj���ڊZ�?[�	�T?�������.��9z�Kd�$a�?X�6���JTN'�� �H*B��o���1�~�v���[��Ƴ����C���������	lh
���?�#ї��V�O�\2� ĢtS�s�O'ښG�:�	O��uY�����������O�Q��`Op ����S�;�k�4��Ӹ.W��J���~;�Ac`K�T k���̾"��'t���ݭ��'Ôr�ɿ�u1~����z���_A�h�&/{I/��n�q�p.S��-�p�cK�N�M��� ���*�8|M��	$�0]�7w�$%w�x">�����5U���^������&�Ija�=s�p���!�����Oo^u���O�?��p:6[��]���,K~\�����1e1ޒ;�����k�>�� �zxM�6��n$��SG=R@��}q�Q�� �z�S�����(��j.��J%ً�]��|x ����Y��3�*�(��N�N��ᢍ!Z�3+,��4	p�O^J[\o�g��d�G�/`�L�AR�֤��l(�@��cl��[%&n+����2�,�M�V��X\u��~,������ �PP]D�t#4t��W%0�'�9ݲ$��F���愽>�q`�6�/�U��K8'����m���K�a����C��Z��Ɍ�mO�*��*l�@��E2_��M�H��qs�S>"������C+D=�OR��yK�t�J��R�u.��g/K�s|a�p�lū�O��r]򣖗�"���E+�f��Gt*����{�}�`��ĭ_5T�8�77tҵ����,�U���$�5��;��F�ܦ�:'����z���s��<��������u/��S���}���Llw%̓�@��#�� ���9��1&���ɣ�յ��'I90��N���ʂb�q����6Ze�?�~�S�w�����WLU��V��|�	��(�W ���)��2�;:淪?Y����W#5}R��&�
�$��w��9J��Q���˓�N���@A.�Ƶ��Iy�$⻓ܨW�[:��i�g�\b���Ok�l�m,�8>	�5���Q�(.�_5�W�F"�Rnh5Ӳ	��ZU������b�	m�оr��p2m��VYc����D߷2�N�fB��Z��T��k�"�<-HQPZ@��Cn�
tPh�F3�F���JY�Ik�U8��=ɿKnۺ�6+�#�̡�.o[9/UzYRy�I6��!A>�2��N�?��?������TCF}�߹��LT%������3�I�������e5F�.�����ndhT7Es�Еf�F!f�����xJm�Q�����Sz	�:Xr1�2�ޏ�n.6$N�:�� �ݕz�GM;���90 #�`���a�YU�:�U��\')@4�c���s�l�y���]�L�
�K�<�O���Ǫ�Dȸ/~/9/�#����u�U�c`[�#�����d6��q?�q�}�q�(�JX'ȧ�b+uS��R���J@�X�@(�kQ�U�|+=�3���M��!㶸���F$h�}qM*m�,k?�^M�+��J��u=E�t	B��^f�t6�7�E1��Y]&�#~3ѓ��@��A�G�#ٵW��]�������VE�1�w�1�*�gҩư�_���q��lXo4�\}����e�w:��/J��U)Uĸ��A	7��yu��0ג�����.�FY��0��s��݋u�q�!����!_���Ds�Qs��	��{�SK���>�#Ia�+]�
��;�|����|��!��.p���)��ۄjԴѴ�@-»P�j@��KV[��_d���.�.w�6=״k�t��Z�K;l�H�%ϰ���l}��j?Ō�¹�������ORJZ>Q~D����6��E:�l�u�9GN�Ϙ%��3&�C��qdv�W�pL���;��x�N�%c����s&�������ط���n����J�^�V�c���PՅԾ���sG��v�po
ľ��5�"���!*�W��0�q�s�4[坒&$�r/O0�7z	���*g�29�7�ܳ7ik_l���b~g]���Z6���k6�1�k���uq�f	Z���ef%؉/U�A�u����b�
=|+����i.�,x��<VK;c_�i�9+�5��~W��bG����{����-�1|�/�?�����H��Ñ8Yn]�w���y\<h�dz���_P������6���O,pL���'���3�<EӼG�/�m��� p�5�57�_�B�^����hN�6���7a�3��.��*��<�mŖ@��+�y�][|Y�������i���t����#��'s��i��,u`�?����qg�d�G^�>����r��ZM]��Bش�s\�S���WV	�'�wW�x��	���1W_�=��>"\s^u��>3��x�i&T�?�|-��9�1�:��"���A)RYe*���s�\�1F}����޲�,>JG0�7T�����V�0,%}k#�Ch��k��n�_(�C%:7��q