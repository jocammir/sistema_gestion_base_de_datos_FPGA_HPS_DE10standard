��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0����_���3���eĭ)|u��XXp�>h��m�g ��.vdZ�XEP��/���e[�`�Fx8��3�DѲ�y���������=���2�UB��:�vK�w����o�0�?#�N\�lX!�9
�!;Hh���r>���a��?��L?��#Z9�+00��([rŒB��f��]��ÿ~������6�s�?��7H�2��YPS|�_�{�n�^��x��6܎e�G��^=	�3���kb��i�M'��e�"�� �N.{fO����f�}	1rat�U�k����Y�
0�&_�
kS�+�0$${�+b+�f�B�q�s5�����ʋ���|'��j��Ê�Y�G���^Kjy�hV���L|D��T~�o���W���`f�n��yVUS���������b�-7�� TB����<����p1�v��߲>���2X���]�[�;��&"��/6��}��мſ��C�(�,#�S��Xo�l�z8t��ri����;qr�g�x�R�����U�f.�A7^R(0�L0��S�Hp�Y�z]>�c+X������.h��S^�M)2ڥ��Q��k
���Y����#G�V2�X�B(���P�T�Q�	M�ͻ���Ű�G�i[�uƺ��Q���O����\�)%!:� ���U(���!�v�Sh��{�	t]�R�M�-c��`I�P؁=�}��hӀ�Y����+��{��,�{�N<T)Q����ja��	i��U���90C�2C�&��;V��|��4�c�}s��}�!I��w��L�`:j���ךw��K��RG�<>�q��S��@�JM��n\	����o�/�kae��":IHU;���}1j�����E��+���;A��oQDm���#O��
�o�)J&�S`��yc����c��6��T���^�l/�#r�܊�{��÷�]{��v�)8#����ޡ_���G�9�5��d~�j��.>���Ƨ����)����g7-�����l��l�1��
3汉�͸슾o�!�#2hG�?n�E�М���-5p�]j�i���*�<�p�H�[.)����b麗��ӆ �U��A�����;B\�����a;���?��H�$���ӀD�	�z��R�K?͏�1c'���l�Λ*'�e�©;�!R��ʜ�WsCP(%N$��]y|�>�MX��9�d���S`�fA���B?��jcj�֢�~2ާiL�	  �O�5��1����,],�s����Ҕ�\��\Z����3ɖ���A8)��; M6X��x���9�C��XE<!� ������;��s"d	��LJK춼�f#��� �EN<u�xv.��̘>����<|ׂ;�j��RZM����:�,hM������F�~>����G�w������=7��T����n�qJe%�����UX��ឤ>��)��]���U􁯸i��[Ą3A�NymSǃ!�S���%M��An��2��H�3��Af���g�&����2��b^��Ӓ���T�̸� �و9�48gA(�W��l���f���5��8�ڲ�I�4�H�V�L�/e���Z�oD"��L��h-	�`��� Y�{�F#��e��]�Gc��&{zS�T]c����e _���/ �{* 3#�
j�"��|��jp"ü!��[֩�Q�[���[�T³ҳ�C;�~3�&���y)�m��S\���3���f7!��~��1�थ�wpv��En}�BW�q�L �%5H-`�W��=�?!ɗzgf �$CFk L�vZU`�*o'�L�>J��b��b�J�m�Ɠ;j�a�DT�6�}M#�f�����N�� ��������e��;J�#�lM�3��.ޡy@���ӽ�"P<9�)����G��mj���4$w�'��N�~�u%݉�
Z_vi̓����/�.�%��!!�������lC���[|�H�������W�F�-�҂x�+�qH
ؤ�t����5����k���JPJU�����҅�u�93�l-��N�O�ں� ���Իj�h�rŅs�hQ����0��AR���<4b⧷I/���ƒ�,_�J��]z�uӥ��L[-�;Ă�@�q�O�p8񹘀	T���9�}S4�KI(� ZH<�$��؜?�e�B�k�DºQ|���8T��vb�1��P�R�ɐ�2��o�� CƧ��F��0��j�~(ir����
t�F�x)�����a�j�W����S��������U�I��k����i�ob�_���O�7	�M���(\�o�������zK;�։��$8[�ea�
4\]bŃ�ׅ͘ �%��u��%1q%�o+��}��B�c`�4q�A�^�oy�Hڛr��ӯ��C�KyD�#�!>΋�ap�����굝���>+�����y=�����N1�Mu�|5��Q��1����5����ױ��^,.1���3!M#�H���ϵ��a5`�)�*Bt�A���p�iư��t��PJ&h1�>�Es\q�Yt�~i�`I/��A���h9��03(6nȽ<$e��L�H=]���kR�U0�S��@�8oPJٴ;�I���U����]��dt�^�2\�,r�Q�+~Z�7�YWNL���'�m�D�:/�T�Ǫsl,?��;\"�sk+h�y$�8�-��h=6�N�����qu��K�ħv`�yh<�>�s�Mg�ЗE��OU!tPUnQ��&Y/��E�����~�H)�a��W���K~=c�P@OCC��]27���}���R���f�ؿ^��Q�S�'eշ���Kk��}�z�YJ\�p�a� ��9c��1!@����f�=e��a�=Qn6P�D�s��7
�˟�O�N�����<�������-�q!�x�R�]Q����N��s��`g�wq��VSc������Qyw!�(� �^�n�LE~ײ����t�2��V����tL=�g�K�] ԅL#e��F����� �G|�4�-jw�O
���M��z��q��A��}vũ��[�ThM�0	�=�)rQw��rٓ���5��IV�7�༞11n��jz沿����p�ZN����Z�I�=���56�,tR�Đ;�́��($��#	�:��N��y�*^�%7$�Ψ����=����O�hڃ�_���tP�d�� ?��&��j9a��)q�Z�	h�h�Z�%w_5XH�#�d�ÄG���"���1Ã@d\z������w�7qF��T��^�صu-��v�;��bB�I�,���]1{�t�8tFHW;��<��=7n2�>]�-ߍ�5\�s���Y��/_�)��8�٬�V��9J]�a�l�&P�$��p�J���F�8��&�	
�2o3��n����5aI{�~�Q���}'��Y/�AAg����`�ܦ����>'me�d|���G3�%߹����}�^�F���o�P�Q�aFTШН����7WC=��~���s.�=����]n�s1��xL�G1&=�	Mj�DD�\ԣ��_�<K��^�9T��pLqYQ�_�xUt�A�r�(` 9�������{�VM�$iU���2�IP��y|M��92�Q�1@v�lC�.-'��ޏ��u�S��	�y�.x-��I��-�>bv�r��x(�O��k	N� ��R���������������׉�ֻ� ��/غԿ|��ĕgm5 �Bd���_�m~uGƏ�67?c���\�y�6�P6�5�&骝%x���+���Zs�H�Ӂ#�su�u��:J.�L+YK�.\���3k�89�9�*����twƟ��F�o��{�ۙ`�y��Z�b�G)?��e��"U�	�& �_g�����R'Hf��
;��s�U�Cv��9�WპP|dVB&h9�����rH����^���m�:/��v<&l�2�f�pFR��-w�LS��*�$:I����� +/�uUV��ۡe|���`�k9%�>�!��G�?��"�"����g(�єz�J���d�56�<�xȧ�f�G�]���OקLK�Zv���hl8+O��[����}��7�$6��5�g� �-x�[π�����b^���#�T�j�C�x�"�U����7=�� �'���:-S��}"3e�������a{j:��b,�j:��w.���� )��1n!  O�'
���{��K�s(p.���>` e�Zr�~ؾ0쫦�^�+e!XW�p� �Q���g9��\<G<L"�q��p�:wqD�]���B�1��F�8!�>R�0p��d��ki������sX���k� �/	ȵ{��5Z7!n�L������u��M��|-�c���.3p�ʑE��k.Z�J^��H>�8�c�
p#e�t� Ӱ@,ح�G8��ӊ�l�MQU�����ed�dW,�j�`�!��o&&�S�5S�W�3i��Dkf�t��K#Np���('�W`��$l9˛�{����S����p[+�T3�Nf�2��/!jh��#��e��-���(�N	=I�����t�%[���-�O1��NDO^ Y�rI���n-��.���U��,G�8&@�9���,Fk#V6n�@���\l-Zp������"�(&d��6|��T$x��6)�lK�PS���<��lK���2��9)������;�P�,����b!	~O[A��@=��#9�[~�̬:F�L��R`{�����C�)h�	�jģ-W��9�����o��f�HG~c�"p���/=c�2��'���VA��8+�N^�&��~�߀�����l�U�"`m0���K{�!��B�;ąjqb��dy�h�/"�j>v®�P��#�����5^��7�ȕ�y�W
N����|����\<"�V}|kk~��;ٕ@?����*��pa0���y���g��7�����W��[�!������_{�B��Ȉ{	��`���%�%I��5'�z9��l�?$�,f�u�:)}�:z'����!�z��/p,\V�){�6j-!����zb����x�iMM�|I�"ʃ������ef�V�lČS1P|{��UJ�޾�W�������_U�s���&�#�=�#�NԬ�&��%�c-�G�Q�iHL�J
������&/��e'#Y5��#�G�����#�|���HQny*��+]�}��p�N���GS,�ҋ�tNQ�_x��W�B�^��<CHu��%�0�Ze@�C`�> �@?.WȲ`�`��!u�AI��3��W�s�g��bjd�62ԹQ_i�
�ƶ�%�ǲ����Z#R��˘Kx�кo�[�Dv�^���R�ߕ�t�����%�F�#�b\Wj,��G�K�� �)�6�P�WO�4X��P�Sd��j�e*J�-3��K��L��)���lI��:�LJ$��S���aɩ�8
���"�1�Xߏ
w�����j^�F�ē�^g__��A֤-��T��˵��[N��%w��ڈ�n{���22�m�W�i�q�qq����[�/��c�?0e3�JJ�@eɶ��	}��w>�g�N���!}�76�~�
����/;��$�M3����$;��.GF�Ēh��uA���{'#IU'�5��z��a�̬uq�e��,3�����x���v��f��ׂV�n-�ζ�s�t����e� ��\����à(��{7;��w�N�B�.b���H%VY�)�c�{g��×8�Իz��~�ѻdI��x���-*����8��sۗ9��k����s�Ӫf���
�����aH�3S�S>j���́IΦ�k��3�OG	�|��?/ 4½>�NR�V	�)�A�$yf����ؑ�w��Tv���~�U.���2]���f����=݈� �w�F@�^梃"��F�Y�*�K�"��j=���<���mh�&��UM�"�����c��m��lOC�0�Y�&����8)�&��,���}N`����ˢ۶t�J�]�Qb0�b��U]X�uɂao&��aT/��t���>hev��rf<M��i���l�>�oCi3b3w�,0�Z�/����N�����������{����0^O��ւp�KIA�T���?A���((B"Eʧ6C������q�̍���?X���gY�s!����X�zb��W$w�ɡ�[f�W'���:;�a�F|���^���	�]�0��̔a��A�a_���
�D����:��D>��S"��4�GFɛ�0D��	�L'�I�C�^7p<�#�+���.4��ى"e�]A��]���`	"�e����_2�@��w��M nK��Y�G+�9ד�P�o�z7�٘ /K �_�%;���}����a��D��]��S���l�h��f�����K�7�.�Y�<��|O�~N���p��A�\
5I�(�>�ֹ�=q£�3,�aÝa�si[8#�Kvgf���;�fj�J>�tlK����jٵVވ+��o"P�/�ָ+��ǡ�I�;e�y����6���x~�Y�Y�!�l�8���T�9ۘk�)����B�T%�����I�8�I4�	1�r
�tp�jeg�����K����I�Z�y��W�{<
[�@��dM͞����t~U�94��ͳ�R�#<�]w09<�XB�3���|B�(�e��Udދ�p��xɌ�v��Я�3��VI��.�,��BG�6
�௉��u������Ã��� �Х�z�B����9��&YX�����D�g�����Qu��	v0o�2��Np���g��x�!���(��w�*Tk�Y~FT�@z��'F��7��D��,o��<���D�Cn���6��_���\D���xu������V��p���v��]r�zu6�y,�{�%G/�:�
��f� C�/��L��op�Jl��������-�����?p4�:�jM����Vyq0K"#^�5�rM����)̸��κ��a�m1����n�Y�7d�F�#��utj��ۋ��%C�>v�Bp��Cg?th���N�Oc�xx�F�����?�L���CV(������E��N��'7����/���`�>I�(t1W$�E�"Ci�4C�be��sr�5�:����7���T���V%��"�������P!�h��,�+��%�S�T6'�UQK e��!�4�M�$�M�?����#���+*�3��"��ydF��ňnR&����l���,�Y�W|�w��`�%IM�ıiR�=�n"��Al�j{`IY��Ǜ )��h3�����p�䭽^�z�s��1�)�ls1I�I:W�e�ގ��u�� ����7rj����'H�zq/,�b��e�/�M���VZx-K��8
#�	���κW����	�N�&��v�'�\��I`��XUr���b��T����y�Y�����(Z'.
��,��V�_��N������~,1��k��)-줚�>@(�G`Sa|P{k�3�Ȫ<�;LϚ��m!q9t��E�Ô0����a:!S�0#���]��Щ���,�<W� ���H&�垮��� ��ke0�=1���Ϙ���j��q��ß�?��P�و������Z�z�xo��G�0�s��@���U|�y:��H)c<�d��pԴb���'�~��?m�ҌG]pOd�n`�'�+Rf>�fm��u�<v��Q��l�
���W�8`��!y�XK3u��l�J߷�p����У��4�N*u�Њ�p� �����W��G����������w��
_4�PC�0ٝ��Y��ų����\�Z�`&D�Ty���z0�rب& 8�ԝ�}Ͷ(��)f@�3[�Ȉ"���S:O�Yҽ>����0��0>p��	-A��
b_:�<���é�p���N~F���r�ǀK����oJ�l�]�'�E_Z_U�7����h '�
�^|�HP�s_-!V����� +�|�>M6<���,���\�sQDf���i-���>'�:��-a�ȓA��w�YܨfO�|��Qݞ�Ё8�D�J~]���������?A)TF��٦h��2P{++q�O~��%v����?�(�����g�Ko���e�:���)
���qR��%ɥ�$���#SM4:)��q���'��񮴍��_hn�K�*-����[�@��2Ta��� ��֒���S�E�:��N���5�X�0u��,���9����6H�b�tz��/�	�L�.ge�ή���h<+���%�����}��:�Ϥ[vmx,���ŕp�W�Ć^je���^��榲
]?)-�I;����?(����$�	���Nܻ1�Xz����5��r��($dT�Kv����+�7�oAA� 
�=7�3�O�b��S�ꮘ@L%	$���v��A����BI? �3M�Ԟ����hmƌN5�����ۈ5�F)3`[Y>d�F�ciT*�<%�8ċ�(/���7if&#)�4Κ.�vU�r�̈́�],��%5PՁ�\|���݀��q��~�E=5�7����cZ��W�_�Bh���D��0Y�GĊ��a�u��O3� ���an���N�lX���A~�����7��EX,ȍ�8�{6m�@یv��,���a��ؐ�I�U�S���k䝎�:׭��Ў���O�]���R�^꽈5+���Vw'�^;���9��~Qo�t/A!�O�R��k�����$x�7���r��K%i"�cT����Ey`,�%��ֈSs��(����w饄�\�����N��C7����;�T��|\#y3��jX�F�{��<��� J_�	#SU��[�ä%�8a�x:v#Ȍ	�>~�}*��R��Z]5/�簮���(-bTt�<�U⽃uMR��QA�_:�� /Q�pm�,m��|~h0�\�ă�-�rp�{R��D��찞ж��3E��[���?� ̋5Ja�jM���@&�V	a�����~ˊ���d��Ty�����Wۻ0�EĖ`�!g��C�c:�G�Pݙ��GM9i.��Hxٜ���5��t�����2���K�ڠi#��0�A�X�Ε�b�C�K�&�K�_���
���Rͬ�8%I��?Z7�d����LVf�ωh*�wU�x�%p�fGV���oW�O"�9��N�C$��$���v���8���i�Y��n:�3�p�_�1=���Y��V��$�+���{�f�"��b�}*d]��Nq��U�`�1l b��ѽy�!W^a�[[�Pa �=��	�S����`��*�_^��{�Д���
�A�)�1
*n�HHVm�Z ��S��AU@�9��Y�]�|=1#[�v��NS(P�
ɲ���Fʧ�@<T����q��v���ߟ6��(i�AF��n���A�{7����c��"C�)�2�s���i���~��z�ջ�W�D�A�����܄���ԙ������a�܊� w�!O~�����6��r�~�:�~��5T�0KH���ؾ����PX���ɠ�(O�GU��@(\V�>�ί���+�e�X+p7�0�j�1�>� ����z�}�,��S7?���""�%�9�*�J���~��UiZ���R��G�� �B���!��+�̚�0�Pe�U������,I�.mV����g����!:���Q�WJV���<�u�DG�we�6aH�p��v���C�
ͫ�3�+)r�N�|���%r��g�K`�<��;z����+�W��ǌ�A0I�^w�b�p�t��ډ�!�9U|c;Z�'����y��e��})�1*EMs�|��@��=\>aF�\=%="��$3Я��7���H�^��E��� Ոz������i�8O��:������x]�1�hx�8�����ߏ�x�͚�J
�Sv�x�f�tFOgL�K'3�h����۱� _�p-swk)����qh[0^�M�m#c��SeT�5F��A��Kf`���g_�P��]��"�|��^u��a�ʴ�@f6�-�{����
��h��>8Jy�!��9�rd�E��Q�/��\���{mF�ŐEZ{W���$Uۀ��m��f0r�1�af_�b�E+PG�7�W�c�����2B2V�:�Crk�s�U(��Ֆ,��[���UIFd���X�"������3�ά_�v���MpNlԳRL��3Y�FMo��D �b�O[U�d}W*Y6����*���.<�����4�4�WJ������g�����E��%���p<T߸J��C�������DLXZX��mŁ�Ļݩ5�����?:��<Go�C����gwȕ�u����ʁN����X��l�v�7�:rOũ!��2�8WM�$u~�FYDix���3�]�lB��y_�G8]�^z]%#��`����_���yr�C�oN����������1
�aEw�5褳;����A���̜)k�B����w���ħΕ ��g�T>ޫ�@>2�Q���>ڽ"���v��C�y{�]�	�\t�A�O���f��26-,C\a�Q�@�g��؉����S�|���2��2Dl
2{'��߹s�,/O�^tq>��mC`�u��4H�E�3��S>ցG(>&M���w*٩ꌹԆʸ�w�S�,�Y���)K��*40߿	����\���$Fe��	Zq�s�&�
.9��G)�
qU!�_��Ӂ����}��2~
�ay�E�a��TJ"���G��^�$? �T�Ĺ�I����˪i斆�����,7k���������ǭ�����(�J�嫃��u����d�Z��ށ���D+�h�zNI�Z]?�T������n!r�
��-=�w�D��.�tf��R]$�n�	�}��'�]=׌V[�Շ��>a��N#���s��Tf�9�	�/"��\j��C*J���K�S�$>����ٵG���2�#<l�9��n���{Fؔ�Vm�_˚���_e4'�#P�K�~b]�:W;'��p;�p� 4�C��`������Rz7XF�8TC� �S�\i��e���g�NJI���d�(r��H@y�\��"(��1HM�(�X��B�hb}��Q��J�*=��=/nWvf�z�'o�\�y��γ�l�Xm�0%������H��tcE�E9㡚Q�"~^���V�)�f�#)X��6c����ZoyT]��?�n��� ��d#���3Y4��|g X�41�T�D��mzXd��(:5Yk�%"�� �%�6��I��Wr�\��4���&�~��+r�& �ű]?�7���^O�"�T�b�����/��UCK�b;��ҿ�{�*(��	���}Z�k�#�"��Qf ���=`��)���޽�N둣��W�9%�O~r&Ϡ�~Z:6C���G��r��7'\��ں$�2��x��^�x���a9�w��2(��uQ��/?�-��҇����vY w�\LPz��SD�D��a�wi����<�A;�,�Z �7[����!��j޷r��L�hC�Jx��H� �ү��� ������oG2B�h�v��F�wX_k����Օ� �eq�휜��g�z;Ҳ�])�1s���c�-[`���,�VӸ�;��Y��T�c�q�#���!b� �n�m��B��#�T��%$�t$���&�����G8��`	��Js�`�8_����ı���,�\Ϊ7���/�μ�`##���P�և:�M�B�PK@��l&:���H��z
��c��צ=kE Q���pa�5F�˹�Sg�~G��Z\wd�Fx.��s|��~K0���2����*ec�-Z�]�/F�3����]��A��wu�~�<h�2{e x��M�����/ɪ�6t]��,
�o3�WU�^s���4A R��5��"�/X�h������t��p����3�c�3.#Fos�q|iZ��N�E+{�c��!3^�4��l����^˦����_#,N�r�E	)�!k/���d�"_���t
�j�7�7l�l�ֈ���B�Fե8����i�O� ��gb=�<q <����W�ƂZgԫ�~�	�OM1�����ݼ�U����{&�]�%���A���nʻ� ��CHnM@<�p|�g[�l����wU��G��+
��م�0�f�=���9�����9�V�9������N�C��V,Z9O�<� {U�0#*�M�	�<�޽�I�P��Y���	IYȧխ��f_���M�"?5���9�q%4e���K�������?;�V�D��b-�U�J��+0�L�!"9�T���4ƥ�k�L.%V�UW�����O����Y�tlq�� �1�2��o��ۆOL����3�>C�i���ٔ��?#��:G�q,r5q��6���S�2-CFi2ϋ�ޡE��+§��*|��ޝJa�6�q�	uލr�tR�z���Ǜ~�_��tv�z�=���K0T Z���|ņr�oq��um�v�z{7��:��H;MLV��z,;9󴗁%+痂AI�i�黣�� ����c��IF�`��b^�P."��KI�e��F�k����Q< �sy��+�R� ������Hh�G3�حk�������Ϭ�8ۿ3��Ӄq��Jn�:U9F�b�4��u�@�V�=�s�wɃ㡡�~�8�K8��t얉����˽��;2�[���Io��7���6��ZX�Y���	5LՇ�� ��n����}���ܬ��#��W�E������9�^�9i���n%i���X�O3X���Ҫ)��D�(�7:�w�c��2�d�����`%\��<6x�D[����G���y�ę�D���K�?_+<�X�a�'� +��0���3�iH��9ƜOz�uMd��x��X��;����I�#�A_��&�V_��ۺt/����8_$�r��`A3(0�+�뙊��c��;�o����6���NP�S�q܇�#$*A7=�诸Ѧ�����6�q`�Z��K������`@�x����=�M�Q�T	�2�^МT`.�,$�a��"9T&$ �n�1.���wt��s.b^M\Yb�t2R{�)��@j�� %�|�q%GDN_>G��[@f�Q���Fn�Ќ���䯰V����LBN��n��Q��YpC�[mgm"�TA�/�J���-k鶞�ݨY�w�G'��F���Q�E�ږqyhK(��-fS��+�ⅉ�4&�:m��F}j�t��%�&"����4-|�(�WV0��WՇz�����t@渨c�c�B�"��.����Z�;.������gU_��|:���	j5V	��3���D���#U+�U���w���MN�@j��P��'�B�����*L(���>�uvm�������ͪ���	߮��fuh����S�����K"dx�k��z_Ki����$T��:ïu/�d���Jjx�a<:X͸���x��~�4:�If���Jb�o�}E������^y��-���wB$.`M�����0 �u��E��c�E�R�=��4��i��^�;��W� ������/Y#J�R,�*#(;��r�O��Xr����]���<p������L�hT�J%����<����l��/,yg�?,]���u���J��7���z��E`O��D
 L).�  �S��c^L�� B��n'c^���rߗK��}��ɐ���Ǯb)����ɜ�{c
w����uR�˓����)�Vܷ�X���횦��#�f%J5�[�Snd(ȋ;��օg��ͷɽp���I�Im�D���-�T1��Yv#����EHQi>��R? w�j+E��r�m�[j��;D"ui��`�jFt��	-�ΰ��[�����&S�s��z�W̶�A;���(-CF��Ro:0,�dZ�f�0~����S���e�غ;�߿�Ǹ�Ю��?b+�l��@?��b�!�'i�z6w�-�����`���)�u@�ut�EJ�c-W�p���j%����f�@Tޝ]���D��{��Tᰈ�S\t׌k��5����,P�lE\Ы�ZuM����Z��[�����P!�'	��?>���ÿ%�O�C�#��x�E���6簧1 ��.f�tǎ���D��.fm� �i8�8���{��Z�]���99FR��H-���-/ku)ە��7m�M��=���0	H�Si��F[ɰr��;��]7�:�^>"��%
�+�� �x�� �a�YU��Z_��{&��9�R���^�C=�$F��%��'�-��m��1{�h�j'cC�QP��f�=P,�/ϝ��kq[�7��ahE}1��@��s�����K��7��.n��	���� �!B�����"�rk+��{I�Q����:k�;�P\�c�G!D�'aH�> r�ܽ���,��ެN������q<>��:)*��Ÿ�YO�^�k>0�9���G~�줬�������S*_����;yZ
�¶�)���>���d�U�#3�6�%�����>)-E�ش���K��+������l5���n�m	�b���|��o-p�Y`����gZ?/�����6tSꖔT`)�|��Z�ǦI���H��ى|("�X_���dV�7i�^]x�����f�!�N#�����1զ�8C��(�WZ�MΚL������ɽ	�z!���X���87E����Mз�A��k�?r�&�X߫��-�fȴh�o��T���[*^�0J=�)b��=+�x*7ͷ��_����t`F�;vP��~._\�2�Q�C��WS5��&q߰�5)}E��`iϾ���@Ǒ��Eϥ�����wɀG%��_x�Jΰ$�2_�2��-�<�J��(��9�c@�f'�w%D�ꡠ�\�J!�&'O�0n�K��h�T�L1L��_a��Tt�N�t�|�˚���l��f��0�ě�M��;3쑧$/��I!�39�<�^^�K�Z��6����/���"����bl4�4upj��HG��2)��gr�ϰ����T���kl'4�jcae_t
���cϚE�,�?�v)��
��+�K��J�WvԮVz�XMI �u� �U�\��k�C���`�Y��a�q�dNr��>3k�W��"|�{���*�P�uT�[�LXЙ�������}@�&E.�ZH�FKᮨa��r�$�F"�%�#N/�7�+b�?ߴ#��,{U!��X�[I* �'t:�&��@�7�j@�T�x]�C��=����Dō��Z:��-8�I�+���x>���U��4�i����<W�x8.�d�-MV|e��m�ll�L���e��Y$ۚ)1��
>�4�إ9�v���j~_w:EL�x�M�h��z�q�Z�6��bK�|����x}�ܼ�!��D���e�|9��E����s��w�������Q��0DBp\���I�29�<�����;� d���=O?�o.j���t�/l�wB�d�gj|����&W/��G�({���Q��kضޢ��̘��@;ޠ�o�\���hE�L幯�IL�� X�8����� �6?"sxn˃�.�2OՔ��;6�t� a�1̍m�>&[)C�c�H���^B^�;d��duӧ�:28fy�����ê�Li�]�h�^���0�i�$��l 8��g:�_�|�[����=��lE
ف'�*ZjM�/{����#�b `��8���<���y�ʹ� �Vw��,tCAm��&�u���A��t�%�5��k��+U�j%��y@C��
>h2CG����e�>)b'K�x�I2c8|���[;�oz,׵N�c�T�O��}���
��L��̀bA)�j6���r��mZ�������%l�z,�I�l�(�,3�1�R�(g��?�vx�*L����O�U�}�h���7|�:�ta�n6M��x��Vgݦ��W�q���f�퇡��LQ\/#J���H)�(e��=�a�K5zK��ث�Y��ܵ�#���kɗ�]m��^�\�T�D��]%�����9.IRpZ�2�ϧ��� � ���3~�h�@��v���(�v� NM��Ad���W��}e5+�B���,CR��N�_�'_Z_@O�G�jW�w]��|`�� #c
�f���R�2I�	2c@ͣ��w8����+�i���xZ�$�6HV<��Sd���.y�$!(:���QW1]�VsΩ�;��bQ�5��ݤ��b*r��ܖB�� �4�"�2#�$\v�m���o���[���j��[��U�%:$����m#^�� +��)��Z��Uo��*�6�;�۠�o߶9e<~jWBf˫"�*�W�lRq��a����m�$'��ǽc�uV�E�Wf�~����dp�3Z�+�z�"ʵj�<\L�Cܖ �MM���I�%�b�Kxl�EMI�b����R,�:NoN��.Q��݅.��	8@\F��e��BS���7� ����g��(�-��\�b0�r��KS
�0U�mYC
��
�s���Ӧ�d�r�-K�:7f�#��-_����E*��q}G��*���� �n�p��$KG� X�i`����t��>�L���$DR��Q�`��d&
�9ю�S�6�M�%ӥ��L�J*��#td���5�Pǂu�"�l
C��񷀝R^L��X$Szw����q����8���H��o|��xZt15����d����C�,Zot�x�o`�؜�$k�sQ���;�e��dvt���wD�fdg�_�>@όఔ���Ŀ(ʵ	�o�6�#�fV�ګw��J
�_`��M0� �w����xn5�t��J��Մ�Iq�z���Cc4�_�}|�؆��G����pM��.�}�>�J�
 �����ͭ�x$�n]]���(��\My&���'� �gǐk��QH5���8�ŭ RA��0�~�(R����W�I���R�ո�l)VU�Һ]����L��i�v����FT�5�����i(X�k�i�nA�y�)"�������u�G�JC;��O(�D���dey�AE*� j<bGܤmju�/�����$zzlr���Qd�LjI!ˁ�!��xҼ�Cu�0?�ԔA�(�qqه�5���[eۄ�]��8*/Xe�������E�!��[-��}`Fӥ�C
��B�E��V����Tp��q?:�A�օ���\Ԇ�?:ֳߏ U� }�	+�zNϧ������OѠ�j����� �bO��`{Q��)Z�X���	4�Q�!ǀ�{�X-+��((Gq��}�;~���H��#��x�e��e���]T��Rٸ4�m��n�)�S����ZX�2�� ��['6g(�LD�k���&p�Y�w�> <A먆1:'b�}F�gk�N���KШQ�H;`'Y!��ӄ6���.��\���<v��J�Yr�����am��7�C�_Z>�$�Gx3];�Z�]qXL외��U:E��$�$ru�_��g��6I�K��N�T@�H,k�1QI<XT�M��G���Ct_rp��պ��'P��e�w, �WPپAH&�1��})��ei��7`�Đ�wNhգ�ÿ�-�?B
7 Z%;�b��P��phf�c���j�TG2L�84�	A����	~����ш���2?U���W����L�r��]e�tV���V]��ݑ;���Z��e��jq�k�~�s~V�PR�luU�0އ���
�q}^\�V;L�
�\(�\T�%Ԩ�E+ ��o�X���h�Z�@�k!�s���v)_�,?1P2�i>�.CN�Z*A��t�v�1�o���Q�%���sٿ8q���}��lv�#<���(2]����b��ߏ�.*#j���`vx�{}cz�q,cS����e�HE�_�8��4�%�v�t�7� �Pvצ3�aF\������W�83��D�V�k?�1��RvM��́ \�f|�����:5V �E�a�#�.���'A�x�G�N����qO�U	g���u(k���XOT�YWN�\�q�ʺG/�$��e�Y?�	��V;^Itߏ�H����Cf_���S5���1r�O�߶�O���C���=O�P��7������Z`ܾ���sޭ�:��F�Z�8}�)J�
��d����f��ub����RQ]�̱�������酏�M��,�%�*��r7 ��{kc�S��p��VVf�I��T�:��K)'���o �����z�5 $0!��u�����i���@�,����)��l��P�:H�����~Q �'���p�g���:��1�l?������EW�XZq}�?��b��M��l �3ߧr��Ƙ�/��[��)P-��#�;�%�k����z�?X�{���׹���%Q���*��D3M
[/-��U�B5��mp�
X:�,# ��7��R^�c���V����J�k��q�Q�¥�|i߱��m�_��z�lr����Jo@e�б[�������!�ܓ�-���X�9�*ݘx(�}��w˗c�)/bq��r�-I�R6�4s�=����#
K������F��'O���R��b-�yl�MX�S��~�%��~��(u>v�� � �pNI+��Z?K,�Ԇ��iB`S�ew��>>?�:�&J�%'O �Edg�:bǔ�$�z�2��s߈�n�?��d�|.;���H�5��ѿ�C�p`��&@�6r$7�X.���O�NHw,��n@�鑼:��	��
d1�P48�3���iIV�vR%��ǽ^���mx-�K��$
T	5I;:����7��A���50�s�r��&.���h��p�����Լ���A�DEM�Q*K0#G,��ѮL���M�ߗ�[ǡ C.+k�ߴ�'e���v6��5���u�B)>�\����=�HA�*��3�PH>1w�پ!���Qf��{�I徐��ꟾ�j�H��8��eD�n�z���_0�Z��A�����z�R]�����`P��2���Ð�US��mr���/Ĉ}��6�b/�2r3�ݸ"pO���
��FK~���l�9�iT��W���]W`v�9��&�G`6�/�!c_z<�l��ԳӬ�=��?f%]�zz�ّJ�0	�*���b|�>K˛*Ym���u���g��۾����k����"зm�N����e��j�[9�<  �q/S�~�eĐJ�_<lv�-�ʊ��(AV��~���F_F$�Ꮲ��3�>1Qv�,����vx�Z\�l��Ŧ�e�H����Ĵ�,9:C�*�Yҧz���ւ�;��l?��4��5!�j�is�)�f;��&F�oB24;<7`��;5u�Wgoj�X���x!j��I7�L��[�8V���ѕ���?�i�/����LRN"U1oz�7��T�Ī���L���ŝ��T[-����J�Y�Si]�<�&rĻl�hX>�!��A�K��sX3�-r ���j214*	#Da��O��6�&��K��Rj��n����Pd}��Zz*`[f�������Y,5;z�����->,q�ů�s� Jq�ӫ��ML����[�9�(�ɒΦ����ȗ�tkJ��|X(�ǿ�# �.D+o��6ԇ�ZC[�k�W�c���W+���-�a�2��/�Iƭf�>��~m������\��U:��|śMͪ���I�aV�X��C/EY�$ް9VY�P���|��6��k�$M�y���@R�Z����a ��S z/����盞5�����gA�1m��l7W�j�d;����-�.>(�f��/q&�k�PV�p΃p�厞0IA��zB���҃�x�3���|x��$�` N��0=�~N��^V��Q�˙7�e#:=y��I�N����/�Me_E����YM|��蘯g[�u��Q�btz5F���L �]E�2	&Í�I��!h������c"2Ŭy���=og��z�ac����Oc����.�(SӒe����٢E�B�i@�����e�����4P���)�5�sy����Α��3J��1*�H�Ab\B5�l�Y�.�JMtB�L���>�	-�]�����o�9�W4g��~�Y��X���J%#�1�}w:�p&�rx�Q��ȅ�
�
�����e0g�����r���H��(Ob"\Q׳��cN#��x�k�ޫ�e<<�"&�&�$�Q����
Lt�EԞ�|h�MF����{&o+3�߶h����z@�&?�:-ɀ�F�×�c1�!����zV�W�=~$���Hg� �@����­d���"�Zɡ�%�����-�/�� ��~��@��X#iO9���I�75�����I�����t��^g�ׄ��&����l@�N�ݹX�j�Q�ЁN��ަ^+g�s�vf_�uͽ%�őI�{���M
����Y&���N�vX<e�H���}��3��J�G3H�̅%����yop��o�	�
�9�	¸�סiV���f�Ğ�e'tH��|7@��]�]�_`ݴ�Psѿ��&�`0�%̆�<ͮSK���V����0��d*��4S������?��.#^Z�o�� ѭ]�Ф&b�㘻R�Ո@bK�y$���E_���O��j������[#��d3�����߽�|4z���h�Nl}�$ĳ
]�Q�