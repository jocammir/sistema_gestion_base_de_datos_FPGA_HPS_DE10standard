��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��Nڭ�	�����B�#Z���?�4�j��0�ΐz�A�y�[��I4�fB���_Ɛ���-����B���M'~��k,���'zf���]A�� -̭���ҧ���D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T幫$��7��`��$��l��[��.�X�R����W^�oG�o�Ø[jJ�޲.bj�6�ܕ�Iq��]�Ҽ�J�㢅����f׊�c/�}е	��~�ͱ�jA}=���O���f�V/%y��W<�!*+G�c!���@-a���X�����΀��1�v���lpM5�e�}U��
���[���z*")�~�^�m�w������ak{[�A�æh���d��++��0���?�5��C�$Q������b&��}]�3�{ۮ$��2���] /��s1�u�9�8S>��?��!�'�nv�n�3&� X2sPS��\ߐD�9a|o��LJ&�h�	���""��f�ajCↅ���@�<��5{��\cDVB�h7���w:V�����Ȣݘ^�)&���G݆mH��:O�W�:�T^)l6�f�c�<��7"�Jִj4��I(�Rd �^q^ ��!BZ�[�<��C�����!�D
Uan��՛�@�j��ʥ�"������3Wd�ƕ�Od�S���Ŵ- ���#�
�O���VO�2l����D0G �^�8 �`H��?�Cd���=t�c�7j̚b����O��^Y�D;��H��ȪCB,������~q?����O���}�_�tog	Q*��\����-26�ߩ�̾h�����H��w�1F�,O>\��:�����1Mmh��?YRNA�M�3"�n��MWW�
g�rit�1T�
tg� ]�d9��Y~�~�Nt+
��o<��-�oD���S�2���D�t"_�ƅ�BؙR�:�}���i�^��{�y���Ӷ�������ȇyg�n�
�]%�5Q� hS�8��Ա�"%�|ӻL�pp)�ӧ��l}�����e�ҨI��q�2ZJ n5����r���g����O��x�3̭G���Y�y_��П�+H�w̙5a� ��<��6ڙz�0�2�� 6���}�k�R4Y�\�{\��IY��q��c(���Z�r����-Fo��C��#����@�,~ ���14(����4s�'Ǣ�x��������e/�!��b��M�1zAߢ�a�W�.�ℜ���X��HD?��S{�&�/��'0�WJ�h�Q��}����D ��$Ȏ�Uۓx������r�D��e6Ջ�P"?o��q�8��'���~�2	m�`��-���! n���D	 ��g�A5��'כ�[N8J�Ƥ1O��p�qC�˃C̣C��`��
��?�`��B���mӈ����q@�+�S�	섗����q��C=DV8�FV_h��J�<2��B�3N$4�Ǡ]%��2��I�.�DFs�����@�K�K�MZ�3��ʜ	��8�Ӆ�&1z��xU������]�ASh� c ��V�Il��|>%\a����G�L��}�����A#"e���>FH.p!v���|r�'�=�3LZ��>�Ϟ�;���H�?Y3m=皶�⇹����\��1�X6z�}�b��=��w$'/ڎ��}kj��&�Ł�e�4��4�6�jSl#n4cB���MJ��V