��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0���C	�i��E�:r�&���<K��NBEX�+{�J�#Ys%`�{ہ��uh�u�|T��Yi�m~R�H�T�mg��#rd!�B^dQ�*���EFi��+;Y}$�".���$��`�"�ͧLR�cj���j.K����Mko;#E@�Xd�yfh����:���6�=l�⤆�q�����fR��Ȕ�Y�D��&t��x�>��c�n�!қ��0�u#w0�|2�(��kr��~N@����TΏ	>h<r��Y�����;�f�T���&P�qO���1�c���tZ��*m!�5�}A�MS�$D�T���,��=v���^�0���ۍ�跿����漪:�:�jU6�V<z�eu�8�'�fTh�L�l��Z2���t-��S�0\Zx��!����`O�#����A��S^j�IR�x�y�c�D%Ж���5%�	�X���6���ċ5I���wt)�ٳ1E�:	��w����KlMl�ҋ���錑u�P��@�V�0xa�6�q��=�*���y�����!�P��Q͞W�$\�l2,,"_���C/�:~yèj�0WJ��o����UY	���c��*K�g���@"��}ذ`J�&�]U��g t����R�GY3a�X�A��q� <My&��w$%�d]��ΨM}vX	HJ6Ȭ�!���6��O�cv2E`y7i����q�9��������tJ4J_/:�ʻ-�@Y�juh��Tf�&�XG�l�����3���y��H[3F0K��"9�v��S�XP*	�F]�L�V%��n�[%d(�\�=07��B!4,�������s����Z��<��98�o^ճ�.���V"Ջs��^�Ǳ����͇�-x��U9�����t�mn���,sS�VL&�/�ѻ���E�n�Ѹ��w�}un�||\�'�2C���-�B��(�aḬ66;k�{�����ڼ�d��2l�H���a�a������$���!k|�"nҽBHӰ���ԋbtK��8:��q��h�.��z���C�;A��4����7~LaWN��K:��+��Dޡ���趟���
Z%7��9�< k�|��9&`n�?m��[��ҿ<B�<ў�/O�ψP�i��4�Y��\��j{��=��̣�g�	�ۯ4�%�Z�=���=�s�2� �A�癭�!�=zNC[��|�U�I�尯cJ��U��9��d'dU��p�����L�b�i����,�u)�G	�w��ځ���x� ����n��I�a��I�k_b+1B��.���
��G)��]P:=Q`�6 -�Ĕ�T[�i�xcW���c���{���m�g�2���8,��\�d	g��O9a��_N`�$O��4�z�>��.�|�i�X��,4۸5h�A�ö�{4��J˚Lq�2Sҧ�D��5�/nV;d��}��-�*�Z�6!]xX"y#|�L���v6��m�V�Y�w����ָ���`
H&�j+<�_B�+K��;�Uį�$�NR7P=�$��g�J�<#]�Y\�\�O���h�AeW�DE�?[��S�8��:�T�d���g��ֶ5�q,�t)��#D�(S�A)P�A��'�b!�O_3y��9�e���1���I���'���L������������1��鼫Y�R^�`f����̾]E0EE��Օ��=gJIz%e�ɔ�1�6ҽ����gqP6*:�a���%Hs�����^I��o_��xC����'��&]���k\�*��[�̯ټ��
���\��_3DW�*��\~�E�~����Aɸ�UpB�	b���h*�i���Ktx�|L��l��'�rS������륢�.5A���w�) �t_�}�,T-��l�\�gE�����_Ν��o�����Fd&����!R�����Ln�x�(���S
�'�%�\��;���0�@��j&iO�>1�#�eP���z��=��o�=qL��u�,�d�b�z.�D�Sg��E R��j�hل��_C��6S�G���/������e�6}y'_߶@{�X�,��� �Qx��`W�.io#N�j槿�r��U�_T�|޼)$�kp}
�&�6^�c%YPw`�vh��@ٽ������V�� ����F˶����@�P�5�ܮ=�A���f|�t�@�؋�Wj,Ҋ�ey����}Z��n�w�'ʋ�� %Q���h*	�#��N.q�K�Yi��hV�hE�o]�6I;�6M�Q�X�ɤ�^�A��t��!8�`�W���'$GFK���6��ࠞ��iȇ܁v����f�Dj�"��mGן?Σx�n'���\q����\I�Se������WD _�>��� ��@}·m�W=��}��c*t�,� ?�gph���{���٢�'vmS�΍d���h���y�:�#��*$�p��
�{M.R��`��]k��v�öxWF����|3�O$i=�u5D�Aܯi��w�?�w�gő�/>Il���yNO���xЄ,fejom�B�	�+;1w+��9t^�2C@�� �[~�-�����rs�b���䚈�zkG�m7�khJ���&񗦍@�����Cj�}7�#~�3O��4-Rq	��E�kF��;ӮV��!p
@�����˜��`?��y$�<�rD#�3�y��NFC��K�����I�a�/��F-f��ȥ��	�b��0�O及�1C�y�2�F��{��$7�F�?��9/ꇄ:<j	����TI�+7� ���	�ol�N �H��߃����>.�o��eB1eyM+��h�<�	O��E��ذI�j�=-�~�aԮ�����'dsx��E����%t���ߞ�[mo�s,�m�A2�����΍��������D^�g�wU*��Kq�(S�v�NiV,�ǀ;+*�}�6\G�Xj9U�駵��٨3v�ƕ��ʹ�z{˝�ԏ �%#��ct�����y߳��X�)�I�ǀBg�V�aA�lS�>��D�enz�N�SOwȵ�S��2q����,PX�*���/%�}JpEt�_�x����f�_=%�W��廄fJO���Xo^��41�<�~Ƿ,��\���bҧ��,��ݭ�[Ʃ&3Nv2-ܷ��:z�L�޻�ؚ�(�C(��X�E�����Uf��N~3�sЫt��8�a�#%7_S3�ݪ���*��Z9�ëL��1�ɗ`�	� !�2�H�GB,�l�DL�Rp���8��EP������&(��9����>|����Y1���X�#Ǧ���ʙ�_��w>J�ȱ�u��װ9�l��ű;�;_��
턞m�!�2S�T:��B{*��-�Y|P����pU��V�٫�B�dB��z�(!/U���ݝ��$)
�ͼ�9��6�Br�Uul�4�����Z�P���L��+{�-:��-�C"��[�I	�o�L;v���X��b�&PGzN�w/w]u�e��M�$ PiI�����9^Gp���-�rn��y]��q�p�J�s����_�ı���f�s�X�vX�b�q�� �C����% ش�L'�X^��Ss�=��̨�o��5y�k�K��?>;�E�%T�D�������F#>�-�/q�3c؞���sK_A�oȵ%����F�Ы���f�������wS#�t$=~�/��֒p�_Yw�[�xyUS2p��n�'N�����O��ܲqy����'���MS�oʿ�*��5��d�7)z���d�[QJ����W��Wc0��%ko����� ׀�FQ�\=d�q�����X���҃�Z0�"��%ק��)Ej��M(D�e�Pn�9��Z�K%�EB�Y? .�/��L�L��_�6Aoo���C�� `+L�J����D�p��Q�%dg�ɀ���ܮ�q��挝H=�~��ޠG�L{� M�=M��T	�I@���4}L[�ZD
5 JH�,Aܸ��~��H�\|�~��y�E������PHO����`ĺAbs\D]��#c���~`������;�ߡ��=z�#[�\=��+����Q�¦�����>����*���n]��k��e�3���[�ѵ/f�_�q0{��5}bq�*T��O�)R��u�޿��2U�%��G�1oJ^Ysp$�>�&&�����'"��;���yj��Kr\�U;E
���X����M1�����Z�*:b�Ӂ�R��� gh���""D��S��53�!��*��(M�n���߮Ӓ��X�K"�:�/"��j=�}T;������Q�m��7�' +OCj�u���%���4����L�`��?$V��]�u���.Q�_z��B����=�'�[�ZGvzS�\xE�v�x�b��3�-���ن��E1�]�e�]P�j��	�� ���j�C{Ti��܅w�k���z�\��t����uu����B�JʆC��\>F(梌��#�z@�/~cn�!��r�o�� O��$
6mϐ+�����DYg(e����W%"$v�0PU��]�.Uԭ�uDw{隼�z�&���ٷ�R���4r�D����CWwAh�:����
�n/�?"�����[��h���J��tM�V7���)���ڏ���a6?���� �E�r���G�C L��ݻ�.gXa=�����^% ��F�����y�dm|��2|��nt'N�d�A���ƺ�a���H6ֶ�ҡ-:\�R5NR̆K�z.�㚉`�j=��PKXc��Z,��,=��I�vl ���@�8u�,R��@�i�;mW�,�[}�őd�����zc�������c4�He�����m���4~f<{���D�E�p��6���5{��A�	-��G�� <*Wcvژ=����&gC�~�z���
L
�1TU�;'��o�c�T'�{0y�6�����'�k&�l��f}j
�ER�ゲ����-� ۡ�\��RX�˂I���7Դ�eQ��mb�ɽ@!ޛ�j_���A�;P胈�9;�U;6���.����e����	Y|���%=c��`Ɇ3�ϨO�)tȇ	/�T ����~r������G�p?�����5Խ� ;��`�9fK��Z�u�
�q�#k����L�M_�H��5sc\b`��j�^�yԟp���y����Ǳ�v��%}��u�*V�� !����(�pح�Y���@�{���Ɠ��<�V�ܼ��g� DR|�&�Gȼ�������U�w�(g���i��p�ܙ`	� [!R�xgWmU�d�呑MW�k¥.am�J��:V�mF��۝{��í���<�wYm��s��g��S&��o�ܡ�G_��~ �w�&B3Y�֊���Zo$Jl͏�o2��0��f�
	�I�7���;�"���i)ب]�͟V[�Ǎ����J���J$ɛx��Xl��+�� +�̌��ǐY��p 9���=p�o87�u'7�r���I
�K�Q������z�V�`*x9ǻ�t���st�.s�X��g��q�B��=si�u��ůW*�҇�)�����o�u�P���Z�9Nl��}�tً��r₉�����9&s���2�ҧ���8�$��ĒL �K��ͳ*I�
��~�,t!q�H�j5���l�	b�Cu�E����x���i�1߅N�I��0g���gvpW�HtG;ol@̉3�9�3s�%���*}�wF�a�W����Xco����EpS~_�	g幂\Y;���}�����ߤ+ɋqZ�Me�MՃ��$����9�@��4p5R���̯Ǳ����!�ڋNC�@��i�ܹ��n��n]�>�|���Xr�\,ڗ�j8?oNk�(y�F�)9)1�GB�a9!����_�`�nc(�Vu�3�[~m���3�������DRQ��3�7`FJf�@=�'�[*��b�4jZ�5{�����'N��1릈b6u@y�"B8�t^���CrVU{�� XP 7e'W�+���_��(Di�7E�7���\tʓ�+w:_���1�L�3�[Ҏ�{�ua��??3*A�SW�����3�H�����=�/����a�K�]+�L)n��+�n�b���73����W���S�-��`M�򯜨��e�8�=ﺿ�����%��3�eB����8�ј�ݾ|ׇ_R "p�A�t�fԃ����6c�̹.CH0LOD��<��Uq�ŊWXt��Ol����(p�ĵ����pm;"̸��kra�, �Wg��-W��V����/��)�
b�cM�j�o��@�$��aK}�VMh�^~mNz�0�5��ɩ���{�R�2��!���]��Bdb�510,�$��F ���jֺ+�
XG����4�`��e���\_`�Ty�[��򈺌yh�x�f}>�f����-�_b52=·���5t�%�<�散{9B�=/�&���&�K��8P&X;����}U��fLS�
H�]F,k��Qމ����aa��F�)T,gV�M9���=�d��ˌ�S�B���a9i�ǿ�g��Hk s��l��ZmZ�����J��qt"��֑~7pP4��z�c����9�u�Y��<"t�����!�Ԡ���!A9po��;�슊�Q-����Q�i�q��g�W�ᐡ��8}�P�<1��9�+�:�ŇH>� �~tq�u;O������������#�35���ׄ�]u�iœ��Ys;�rM���|�H����>��v  'H�Y��Y�|7Ί��0�� v�,�5>R�Ab�;��g��d�{ͮ�qVR+�O�b)Ya��2�u?bfz��	�s�-ݼ�cӥ���ʷБ��N�}<2�p��40�6r�P*{�����d�
�gzӧ"v��'��*��C�cz�M&f׫���t���2[<����|?��E��E���C���N�:2�����퍪E[�Yd��c	py�1�.P�ԍ�I(�~(�}�����eiȥ#Z�j=�6�s�3	.��\�K��J����L��s{��5�����0�����=p�2�;��;�n�x��R�勠D �@;�:��o�>��x���f\g��u�L���Y=����)$����&1��߲=��{�`?g#�5t���-:S���ryo�X���8��|9�f��x�-��:�)\K;m�
{���5�E�eD�E���O�8�p%6ɇ�4ʆo|�N(��k�lZ�l��S�z�p���V�W"������*�O�ل�OX����Ѩ�>�KCg3v��6<wώ�π�<�i���(I�w���@��$Z�#>M$<g)��ۍ�F3�r]!I$�]oX�~�q}�$���+�*�6��g6��h�#[��=9�eG����4��G�O<�I~�F�=�L18�M<Uk�/�i>�<�$b�yGib���u�$��*9th8VxC�3t��@��ʓ���ڂ��sut䡸���ŝ�)-h���?����J�4Qؖ]�i�k�(������;�my��Fٟ�|���g���w��[�	^���8�`�@� 
U�H��xӕ��0H{����mp��{��y�w_Ŷ�YT���x�#��q�&(��S�&�>bF)9�#�'\`"%l*�N��`��&N�o�?�i`��0�)j�q���q��	*�k�pE(+h:�܀�����?�c�,1��g�����M���& ���[X�����6}�5��9��,FӾ����ng�-éB�p��QK%>�����ݶk7�_Yb��|���>���Gj���6��zh�ܨ�M �cv�p��OZ�ۈ�E��a�~�+�*iR�jEiAZ)/��q�W,��՟�+�ݰ�p�e]p?J�F/�*��P@%U���M�������h2��,�<w��G�Di����4lC�ߊ��\��)�Vs7�<�(|�,�p�[_���X�U �g��H3d�^�dwcZ�lL`���H�?b�7���y��ē��O�ii(8@v(Ej>�a��$fM�ܠ3�����Mg����p�C-G�Ƀ1Ww���ORm�b2)c�#Q�Ҵ�H�*��V���C�vlw6�a�	ƻ��+�IT`Պu�G��f��}%�0̧G!9~�Y)�����jq�E>��thTtt
}(ˇE(8g���DC�+|�~�oTϣ�kg�e�Vr!<:N�q��`��Z|pDog%>��Arؠ�����E��,"�xR3nK�P�ú�ˣ:���L���=��9��jv����Y�J���U��_Iǯ>�q���y0K�_��&Q���A=���|$�9�c����'8�)�?z�cO�ԉrbtH�����Uhy3�!��%��q�����!qt������c��Q�K�&��(�
H*>B/B��H�>Z��U�^���O~p��r>��Wi:�3�?�W�΍�u:�V�l9{��yJc�q���Qc^S�7���F���_�jF�B��"�q[g�ě�=��0��7���s���H��O�Q%2�J>S⾻� ��t�f�D$ܹ�#'&��Z��3�h��o�ht�5�"\5m�]h!������`47�8Eˀy�QVWV
u؟�@l��/���
N��^�$d!	!WnFL;�W�$4��_��ė���˘���t�CK�#@�p]�?�������	Xa�ٸ�io�SxQ�=!��Ew�T0V���%��U�ȟ�a�z��(�@�P�u�,�܍���	J�2U��L��Y(��@�p�nj ���8��9A�(�bH�/��L���q�|n~2�2��Mee-�DHH���t��	�M'��x�v�aIv��!�2�$�ե���a7$9�O��Hk�?'OVHq=������(:�c�*�/��iSt��z>�$�����K\nD�!�oP��kjEf)�7G��W!JU��Ỵ�d*���/s�n�Q>�f��8�'�Q�1uۗ����f|�Z#VO�|B��?����@�E-��ЪH��4�`�9�K*<&�g�`��"��u����B���U^�׉:����� ��1i.XFBr���}~��wWt̋�Ld�H��n#�J4D�A�A��-_���}FԴ����gFt����x�-��Jfc���ĉ5 `|G�Pv�������#����f���GC7��pՓ�9l��_���YCQ�{��Y.qVY6u3�E)�ز���}K�HĖ��s1v�e�@B9����{�H�Bv9�C X2%|g�?n`��&,���grOK�q6�c�k�r�`J*�y�M�ع�ړ
��MYGFp[K3$*GH6� ��:�2XSz>�/r)DO�?�I�S�'�s �.�;��~̽���8$�P��iA���t�H�qK3PN0�CY������a����~'���J�~U8�s� ��׺Z��3�Z1GZ���n��<�{��#,Ci��W_�,����L<������?v���kX:�SZ���m�������E�A��1)��Qߧ ��Q3R�YTqTH��4�ŊN�Y�����x�Wq� u?:�x���Qq�@7�DXtj�W o�����QGe����c�<��3��O˰jjZv���Ə	��RP�+��հ};�ܒ���b�-�z=8����AfI�ױ�[�bd:����E�,����N�=e����V��=,�.6ǎ�zQ�[z���?m��T�X@]�)�Z���kS\ֿ��[u���2�2/��* ����nw.�O�Խ넢��|k-�w]T)�D�~83F#1&X��%c��>�/J����%+|>L��ȕ��侴����{�w�v?Q���1��������*E�t����
,��+�q#�~N�D�!����ݞ��X�mX�;�3 �K���c����վ{�e�H��?�e� �N�pZw���VT�F�&�c�t��_X�E�nA)�'[��e��[.�����A���U��%QK�A:<&�ta%Vx�er�F�=��Cu��F��c�10����E�\(i��ꁬ���8���V�cz���m��Vj�D�ܲ˝b�_�IF��+��gƏ?����ux	xO��������̗ʊ�B���ܫ�Q���w����wE�i�:�D�\����*+zS'C�&�hH�B~Ňa���\��N��J%Bd�6��\�9aG����V'�s�?�ٗ#���"�@�/���}�b��JIV����OO�zX�N�Mf�$��T��2=	������X�*@�yJ�H�!wѐ���Q��K5��/�#W��}��ot�6�Y��1�K��}��F��lU��b��{)a�d�o΃2�PB�-б��҄5��@@&�$0KVl���]�hZ�_�Xʡ��Y���	S*�<�<��3��`����	�lIl0���.�x�%�J���aQ�����;�ӯZώ9�qlK��h�_UA6o��c���
���Є=�m ��� "��s��"ݘwqSa
u񟒈�][Tp����	�9Gh��+�H��=M�g	��Z+z�Wi��o��Y�G��?����X�/赞���,$��/���<V!&I]aU���x �h(x��)Fc�a�"�5��	C���Jnlo���T{�}#T���q�ߵ�3i)U�TVP��mX��(�/�ѭ�A=�#8��t��s�����$]�e:㴍����O@��[�B�9X��J�M�H4��#K|�$��o;K�ճ��g��,�m��7xx�I�����d�t}��`׾Y��UVI7�ʘ(淂�g��q��BTSl[s'�$�Z�K������t�H>��r|�[�#����/^ �߱!߃9�PP���~#��bХ3�+���%��`tA�Yv2WǏn��$>,�a~�O�&wi\C&U���B�E�!��X�6����������i��̻���4���'>�UR��(�<qǆou���&m�/�䣟�k�`ƯdCQ�J������xoD)xⷢv�單��k ��6�w�qT=6x�Kֈޠ:�x�3
o�($��0��S3v$��H�j�zHY�q���W�jV��W���2*Ō��o��LH-�8��L���+��Uͩs�5�[|ঝ�I8��FD�鹗��Y!C� ��V3$fL:�UƦ�/F�c��A���� Nv����v�9�%�4�?��޻��KE���ڛRMq�YxcM�>͘�X6_,L�m���Ys�?2��\I7$S�|j�|b�)8Kp����~�8M��ҝ���'k�נ��Q�ָS\��7=d���E_:DUa�ge�&��Ē��tX_���Iip�A`B(�m(����b:��xetpS~裺�+�G2��� �
�����13�&�`�ĕx�����T���kʨ�b��(����l���J<���ξ94)�|���!��>LV颁Q�\�I�֌�����}���p��e���,OF�	����d���g,E%0q�*0��ű"�S��Uߖ�����);����?�6pǬ�nB��ka9���X�8PLz��&I�.jH�?z�w�t~�W�h�ȋI0�|l�|���� TP�ą��Eך?�p#a���`�X��u,��3��t��԰�3�@Mc!���z{��9k �C�ţ��	1�Ӯ�5�6Ӗ � q�؅����FVK��&��m�)��(��L���Y����⮓p�O3}�v�V����'�Eͨf��K���~��!��c('�ŏ��E���'��.欠h?�/�d�;C�TV�*P���=�6�Ȕ��Pm�N�y�eK�R�� ���r�J)�(�F�VHW �[;����G��k�&V����?o����GQ(R��4��W�^ieX��a�f��Z֤�s�G�z�1�F#���X�����e9w�z�<Ck���z�g���s\v�j=���Z��4ׂ=_a>.��l2LwX�d��_��Aq�Ӏ��>���
��J�`����	��h�ɀ��}_����QT�e�g_W4��A������������J�]M#�A\O�g&<A�����]��N��<n���,T{u��Z�oϙ���MIt�-�K����;��&f)&D��������9�'JZ�&��<o�w�WI��
h�0?��!W0�L6w��ZЛI�J��5����P�#8�mw.D\�ƬQR���eNM%��yE�9�lZ{֗N��c4�b�G}��CW�#�~�0�����E��{�>)�K ��J��3�@a��5�vZQ��Mib�>�<��sԛS���e���<��B:Ŷ+�I=ún��-�{q0�Z�=U�6n����p=JO�1ulҎf�u1T_�r�M�z$���x�;0/:ǁE�H+�嶤�������ꊖ��g7���8�q��ؐ�P�JN� �q޴Vk�S@"��[ϔ�5,-0G��3��	oD����X�3��jv�<BDg�zM�^�\��I�f�R��^���$�J���]oy(��� ��GHGP��M�x�
NL#�������KX&;�]��'3G��Hu�o"4]jn?4�+	�4�����i`�YU4�Ǌ�ǪA#��~��������ʈ�<�IY�|U�x^g��]�H�9�� [�4E� ��QcCQB��*k��n�����f�4e�߶��-�P�+��L=�� ��4)A��B`�'�sr���_���cW�]{�c)f�OI�N�r|Ɣl�TT5�X*-evS���3����\���F�
�]�=E%t	�So�[Q����X�)n��],�d�����ݟ�-u�h��7�#�w�D�T_/iJD��S�k�~�E��޶�l+�蒔V�Nͬ��\d`��=O��Y���#���+���\˦(��#�rj�[�ӂ�F��Q@��B��(��n�@ (,JE����������cG�'���T�5Vk��*��y��g
َ�[�� Ej��9��Or{����6p�r9
�ٶg|�l^�#o����8�;'�����6��)Uf}B1N���.����z=]�W�/�Qw��Ć|�6�ǣ5<�L�/��*�t��p�EКP~�kS�����3Qq�y^�6�yU�U��c`�js��b�#����
�Y���#Ɨ/T������1\���bs����+Q-��T�Wn��P��U�ϗ�Bȑ|dks���ũ.9�i��5�� xv���'d��1�@^ղ�1�D;`��]����Ԥu�-��57*BW�u2�ʾ�	D1c�3��q\�L�¯߁��&� X�RZ�ݟ3T</㝵��F`�����#�5DG\I�OYh�T��Ng�F� ��/,G�SF�׼S��L,���3�����F�&/�N�X��aC�8/ W�B�6��Qs[��Q^�O��Ǹ-�\C]shW��F׍�~uL��J�:ڥ���Be@D'�qa1��+�.��irl��zd��L����;��+
���7-,@n�`'�lW�_��#���G+�FC���u#E��f� �s�歋��~.�*�>J�*�ݷ��[@q^�ݽ$U���=�g��,�h7BS@-G�����DE0�5C 2&3n)���O���D"�I]j����'qFؐa�������pc�+����=�O�t��~��Æ�@�}J_�a�6�{�b%�����5I�c[�@W[��]�W?dɰ�M{�51�#��=&3:Ag���ބ	+�HHd0�Ё�J	�%�<�DV��'T`�RE�ԉ�/'�,%\[δ��ح�����lw��p�=@�)�L!9'#�������ZɉB�����Bu�{��'Y�[�7UbS��\��:�ȑk>U�z�F;���a}ߡ@���������Έ� j�R5��DO?�iub�p��%j�n�yņ^��)��E_w}$��c�����������q^�e.�M�<:��	8��M�3.vZ�;<��47���x�Ъ)!�Y��k��by���)�+�:;b�3V�y����	I'��l����qȔ���.�d�ۘ�K���ڹd�����3����R��v9�lG:hX������#A���!E�3�dB#U)�����)���0n�S���5в@�Z'��H�Q�����B�1��&k�sfr�ɼ���Mt��l�2�l B@]��}� :}UH���ml��r��D�.l��?<������C9�욈�;��Ǿ�B�����a�+q�A�BHBk%�2t.�wO4�ca'�S�0S�ʎV���u�Ϗ��^T�|�UNU�a�l����P�,X��S]8���ᜯ�0�����?������|��~Z〿��]i�+UQ����q��4���H�,s^�N.���RY��u�a�t>����+|p�e�F0�7�,)����y�������㜓��J���_��!Ц���e�fP
%#4<�|@���ɜ>e��i T����!a�K�5
����bJ!�h���7���`�W�o@�4 ��2�;0�hz1}�w��S3 ��
� {��&F���t�b7�Â?"�ܫ���]�U��JP��������$I5�9�7��2����c�"����L!�E���ZN���\�Ռ�c&�����e��z���p��kV��SR�iݰ�����@�R�[e���s�ˁ)����F����7y�,��`F��D9�B��I��{b�Y�ؗ�K��� oX�/��L����ƇIܫlWj�	�f�P��5e���KBgȷ9��)�KJt�\��y���U���3�-Ԟ�i�����с��uMo{���3�����?�	]h%8��`t��= \���W�I���&����}u~���gV��ɪ��o��CJ�'>�z��(=�}!�R�#�ݹ!���	�p��(g��}�AH#'4��꜉n��7�|0
!a��؊���d3�U���'�.Z�orͣ)*V ,�� `���R= ���]�r#?*�%��ّ猟hA����	��lp�*U�<�'�����&��^�H4�]X�}-�T��M����Z|���R�:�����K'{��J �L�yiU<�GFR���L7���Hg�|�q9���`P%��I��{�(�UJ���� Y������w2��&3#�)6&0�Ww�Cs�'�vg����S��7.�pC_��T��M�BI�R#x(�5�n�W���(ր�=K	���O�T�����3��m�+
�3:��Cw�YTl}
���\}A����M�h����V�6!t�;}]�	� I��&c�b����P���Yʢ�DW>���֒��� ��`��wb?�룪��7����Wm欣��,�b�&AN����`���פ.�=�����6�i�^6�v����bv�&�j�����z	�%�s�U9FQf)8If��@= 'A������� ,��؇Hr{��@VJ.���}Ӷ�c6��"y���ѨyA?qU���?P�RG1!0��O<���Y���?r�k�6�XkM@�V8ǈ2���d���I���:�!�k�J�l���m���f�ס(�7\N��8�Գ�Ի�m��>��S:�Xy���܃11� [�$䏑�[��y&&��`qq!ڂ4NY�WD���*��s���l\��dIK'8ZAG��S?�9��]d�~�A/�����Ң��45W�Dɳf����K�'|�Tࠤ{��=!������J��ҚR� �?�q��&@yI��P���i ʏ�D0�Je1; /s�lP1�l�1@zӂ�M��6�Y��2I��4R]p4�3�^���	X�>��P�x�w9@'��qw'�� G91.g��*W�� <����ƁzHh�5�&CF�Z?'��2�Δ�=�Z+�[�2�WBS�+��oT�1��r+1�d�.G"×����2��(��S�	�H���!Ł�����DH�C�X
Ι��D��J����k��ϡ�=s�P+������?�lUPOH�QsR��,̢$�n8����B @�VT�jT���\�$p��!h���ʑJu���`�����
��m��OQT��M^����B�kd�W�Ft��+u��Tù������i���+�t�������N�	��j2nb9e}�KK.M��X.HX�X��v���	�f�A���>���3z}�g�~ 5!`����~�}���.����V��Gc�׼���2���l})�wRG�l�cf8�زs �����V�,�'��w��i�P��ރ��z(���O����sY�V�-��������R:k�_�.�[�"j3�8-����W�%��A��àZ�����F�b��z��l��Q�i��':o��LP0)�����ҷ�N[o7�QֈU�f�C�{A���¾�n��;����}�i�Ie��;~�}���c�1�� �J�2���{��B�@��;%����ݫ�9n[�苂�W|ÜD�U�k?���>畄���ӷ��� �{�@'��o t�Q[ڳ��JԨ�ˉ�g>�J�0�5��^�0[�wA��(�w��^���2�&� �F@�9t����`3�н�����a4e���C���}��]��˷�-ES§vjY�Yf��q��h�+��H�'�p'[�j߽�t��6�H�0&�a��/zۖ�l� �uvm����*����=fK��J�ȦC
����� Ε�1V%9�v�j�f%�0�f�����+���k�Ƽ�p݊׏��Ĥ�s�O�F$K�];�O��zHm�J��`r�YD���p��Xd��*���ޫ+����*A�Ϩ��/��b@�����ku��H�b �?���Ho�HJ�_���w��&:4�9��f�+����jH�.:�g��;���E�E�g#�M���@�;a~ ����Ac�W�0'/çu�,o��yS8흝��5�Z�ɉ�"��}� ���G:���8���e���ҍ;\a;cV	��m�3譡���5������=[���P6�0�V��U��S#������2�ϡ&�$椫l�eueȖ�6/"��\'��`(U�8q ́�M�u�{oy�"HUM⡶��6�<�m:o3����cL6�>��2�6T�����̛p�\�r��3�_��#��djX��szI�*￪ȝ)��l�2�(v�ui�mSZz���oޯEKJ��nl�j!�f�e�w^�w�"$kl�q������_�&�v����հ�0d�#�	1&���U�Ո:Sj&�vPA���@^&�mg�v�Xu��IwVδ^0��Q�/\ld	��l�0�@��w"d�U��1�yJ7��R�`��K�އ���(P`� �����,J��B�3��W�>�_�:����5� ƴ�O������~'������?�wS^$�js�{6BTQ(:1�S�K��ˇ>����B�����ojq����!�Q�'O8aDj�R�K<��y󯩭��'��s��b��ߠU�k��O�Y��T��!�Y8�"
8��އ�t�eȸk0������q�]~��5=�hW��`�/pK��ϐ�v\&}{�f{ZC����O-l}�hig��&X�K��x\络���!nF6-��(�݈����L��E ��I�\�*0��oj�ώ�]� .:������4����-G��d�ܞ�s�bd[N]U�t]t� ������ �H;�F�tӛ�������ѐP�
�N����z���$����;j�M|t�j�)J��3������]�G죨�'���=�R��My;�4k	�dΔ���#�X���&�nXز�_A�����y���6��s���gg����Э0���p���#�9L�߁Na�q0V�K]�����TB�6���&�jue�'X�=�	>2��6�!��W�ЯMj�v�P��.���O��<�~8-��wY:O�6&a7[�B\e�!���*�Tl�q����y�ٔ� �XU�U���"gy�®)*���B��sH�"��n�V4K�:��g�l������l�7�p>������M�,,D�8�$�Pl3����*Eҏ[*�B-�D�Y��;�w	B^^P�P��������qWX���_,�֣9bz��!S�X����cB��T�%�
NΖ ��!����AB���к`/�nR���<���U���̨cG���Ր8��`D�m`V��9�25nf�m��!�T��Ź��$�!���
��%�����H�����&�*��h�T� �:�Tb�A�mA=���q�I�{+@�1���΁ Ȥ
�Huy�Z*0o+��Y�5[��=���绘�j�yC��������V�q�W�Ov��om��8`��$��}k�± �n	nX�!t	5�V��U�D�B��l�`�S�W���W��]qx�#�sj�{�7�x�X�Fǉ�p+N"�a �Ex�jJ3������0R��V[����[�\�NZ�����5:XE7O:�i��ݫ}],���;���8�mV�ۙ���`f���}��`,r�cߡ�7k�!�pI���dS�P��4�GT̡p���s��:�0��^n�,c�4?��/�>g������E4$7�=G`)0]��*�v��I�w[�9�q酇�C��6_\��y?9���,`h��!��[G<ƪ'o��Cw>�h"�7C�K�Cl�$W!e�X��	��2��d��K�ؠ�7�� �[U}����^]��펴�r�*�k6|�f}`խ���X��-"h#u�nt1۴#nv87�˾q�C^r� L
ĕ�ʁUg�(���8�>T2��u�9"h���#���SyLKi"rE��Ku睧�����������z�:���䜿@z��d��e�GҰ��_0�|=��z�������L=u\�G��X1�E6�Z�"�{�
 ��<eR�`�M��G}�h��X�K��2x�oOWA���+N�𝇱pj�T7��!U`YX�S�ecg�m]���o�����K�^Cu��Rړ`�/��N��w��ßD)���{K>���,��Y�?���eIQx�Ut�Ͷ�����:��#KƽFR�Atm��&w24f��|�N<������yQ;��V��:�8k�[����)IW8hvπ�]dr2E��E�5�K�R�@VSQhg0�����ٕ zȂUQ��w0g�n��]�0�Y��bt�e�f��o��⏩1z�1�E�V%^�<������e����)��wqW0WәS�L�qB%�g��&VH���6����1���Rl�t�0r�0E�o@�Q���'�����,�<}��%|�	�z�>���^O�d��~Idѷ��A�����W]�gNu����7�[��5~=��t���,4��o����f&K�xX���
��8����$��0�S:r�<UU��
i2�x�������7u��ZNj]�0���N,�;�h��I�3�,�ݰȫ=�#�樱�&Da���K������i )u���bߢj$ۊ5�B�0����Α�&M�=�<"N�rϺ�,(�
�g��yEܳ��޽G�������c�'z�~z=�$[o��άZ$r���ņ�}{W�<c���6bf�1���|)s�����N���+D�){'�_���Pn�3���㴋b��
��J�uMaU�\wL�C�m{2�4�V��"�[&����&���4�Y�Ͳ~D#LՄ��,s�1���}6���)��^c�=�c����Ԃ��i�[�.���/qd����$��K΁���V�"U��ۼUJ���h�ʜ�:}I#=��7N�4	�BfX-y�ȡ�iD�m�WŲf�HAro#�}Y������MUA/-O���9��L&����O�U��]Ix�^̥��Q��_����c~�ai�X�K�������Ud�'�qk��`�V́t\Z�o�����'��H^O�[G>1�8���o��Ј �Q �@��uH���K/q�_#-}��̌�S������vND�#g�WM�~����ğZ�[=�8�(�	��k�1�
N��<�a<>��k�L2��mq�GX�.2d��K�����jt�n�f6��qjm��障C� ���l��+�����ĉ��=L}�Bk�Z�NV�98�ϱ��&K_T��t���iJ`�����Y���!HdB�g�(�5�d�6��Hx���÷�=2�^�]������
q�e�@6�[ېտi�J@�!��	���������-��&^����ْ92Ɯ��_vS��8�T���C��1u ��PL�nQk���M������>��Pj ��h�p�;U{uf��W%��\��ȭOJ �X��꘬2�	\!�D2�$��:�8eo�I_�y�G�yd��CJ,sҭY�S<����5T�8���u�B��I������b�1����%��7/�&�*�`�8�	W�n��Q���O|*��޶#��{q�ub����n=vN<#� d��]�a>�0y�͔o�je��	:*��;]��" Y�n:�?���'��r���XLr��IKq ?c�8<-|ƀ�+U�Q����5���̾Lq�tx^�D�t�^�KL`�Z�v�CL���<��p�h���cw�#�F'�O�j4�&�#4_2�H�D� cC��(��g�j��,�f���3c��I�ccZ7���31u	��i��d#���8�,�ÞT�覓���J��[�k�"x.�z���L�֨ǲ�F8�2%���-���|p�YlfW)3��=�}��4���z���Ce�a{�$��$�A'�[Y��u�6x� ��w�4h��Z�T>#�P�U�a?�*8?�g-P&sgHaR��Y7'�8���P��_�Et�	実���A*Ģ�
+b���^�����&��
��RJG�A<q��]CA	Hߌ��a�ԡ���-��w�=���� D���X���M��`*��]s�ģ ��1��Q�{��"�'��[��Q���~�c��˼>�a� M�.�\�M&[!�8����@����������Q���t��n�"a��άp���%q�jy��U�����vܨ�-1�|��o�����j�M���J�Q���K�[*��� {~LTWP�u7��F?*�oo�<���q��z�Fc���C���|�����%Sj�<D���ΦL�Μ%�n��a�Bb�D~W ���`G�dJI�uj��>q,�!��$�g+ ��q��M�� v��].�8Uc��W�ASF!�G��n&�R:j�˛��kȘ�� �a��p���ә���^��x��hzs��_Ĉg"��*�<����q%fY>V��%�c�z�\�}�cAPL��t/u�,D��{Җ4�E����+��D���j���S��|���UKW1>��K�W����}�h?��(��W���e�a4f�1��F)�[����=���[2CrqZ��h�b����AkGg0�Kn�w�	o(\�Z{)~��J˱��Qو(�b�Bu@���a�|�ݬw�5b�kA���e�?�p���a�d��=;8{L�;��m����u�����65�Q��2��az�$��x6�t��[:j��V7��\F�{���#Da�b��~yՓ�[�֭v�-Am���TϢ�y�qT�]A���-�:�Sۄ+������p%��'��!�o�!{a쥹�j	&���f�M1Wn޺!8� �pj�x[�x��+����)�=u*�0dG�N&���$.)�3+���ϙ�0ֺ�����qY4V9gv�����9+ ������]�y�w�il'޾���!I�
g��J��/�t���u֎k���	!��BVR�a,������$������c,W��y���w�ꉰGm�?�}�LER�Ղ�|\�i�ߐ7Rĵ�I?��	�����`v,N�%B>-�ԹaE���`�t�e_��������ԝ�K�}ܝ��D~�d(���( ,��=�:�bMgsن'cJ.9��C.E~D�ס-C��~�b�ł�?i������QR"�@���Ú�����U���e�I*]v��=���]���X'���礶QG�q��׮榑TZ(���qt5�Q�a��*�bs�2���42����*pg�~GB���$�XOe�O���<[ȷ._�)Q!Q|4��+��Q�_JR���Yt��l���M����@Q�f�h����̧u�E���>�M�*��{�ȿq�/( �m�M	prYg��A�?�����g��?;�ۗ�J�)�B�kx�����1%�|���l�<����F�i%H�oȇ������Q��Gh`��Og$�U����{{h�4�/�`U�/������Q��:� ��{[��vy�k^�����-���aW��AL,<'4�s���j7Ø$a�y�h��䄬�����!��x'S<|���/!q�o�s��}�z�7,�4�?Mz���C���4�ʮ$w��u��q��ŵ�6e9&�NH�"��M����A-��$�6�}�����*ul릨2�� F�1�Rp�ۃ��,a�5���e,�c&��0�a��V���^�������%
��FP t��RX��F�������lMD�}��VX�H�M����&��k!����@š�͵�F"�$ሻ���KE���2$5Qz`������C���U�nJl� ����%��Z��y�9beusøR]�u�*ҙ��
P�1��#�ix���Y6|<���L�m�2�R�̡R"} .SM����-�[�mOee:F5qõ	�v+.L�i�`�i%b�\�}��ARs9z�O8��Ǎ�4��zR�Z?�E���`kӲ�{�!U�BHlf�N?,���jj(�W{v�8�H��$@
�l�� շ�GVc#�z�ر|p��r6w:'�
}H��#;��6b�8&px�$Æ�Z4�R��;@C�{ &j��!��mD�J+� ���D7|�p�H��[[v��e�2�=�Q��ڿ�b5Ke���#rڐ�E�8y�S�-PT��j��fGU��B��Ҳd,jn�Z.���B��s��� E���ln�b}��~T���ĹZc\ݥ�O�6+����[�r��Dts*չX6%�8{�'�$����%�@8<_w��������-���v��GI0�� ���Mfw$s��}�
�Vw���^�];�]6ݲiH�9����>󀅝cFe�Q�[��BC���w�z}=7cZ����zn��Ja]}��dpw�%���������� �I��h�Mx��׾�~�u��5l0���;r�k��:��y6"�DƬ7���g$C'�4}@���Ob���bq�!�R�Tw2}:�n��c�Sg�k�?���:1�Q�����j�9�6�Q/�T��ru�?d�8Y��y��lZ�^�91�!&Y8�5J�8�\{	���q ��8[��[_��FE�^ԃm������''\�碬);F��_�BR��K�i�2��>�)�T�|4C��`:�����۶�By۞��*���p�퀨ڛ�1a��I_�C��O�Z��*9��Z��}�O3�Gk����o�5<2� �4o<��@�̰r�:e�G�$a�x� ��iS���w��HUI��6,����2tm [|Jw�nS����p#ɕ?C+�DE����[�w_��}��Zt{�?t�� �c�'䯂��"��j������/чJ@8����v��z�<�����:c�t]2����sS�.�:0�g�.*��~)�c�&�\a�Lx�_�pj-��Do�"TR�gT�.yL�>Q*���e�5wC�E�����Q��lz�,�x����q��)��k5/	��!����زܘA�d�G�n�X�__�މ�[�c��Eu��^�����C{�G(���ێ	L�]�vF��hEG��R��≹z-�!�u���P�k�W�
[%BS������8b�]*�I N ��J
%	�t������G�+!�L�E-�Bq��n�N崔�u�)i�i�Mݖd��v��զ����7`��C�EGk��v���0'j��[<(r1����s�rp2"��E�g}�g��j{�xϾ8�H�m�C�s��S�����`/Ғ`8��2A�1�i5�7����@�kVx��3��E<����&�_u6Y���zB,%���2�2�}3i��2�)�1!�?>ԦN�\�t�1֥��z�z����3�93}� ���3߇�-�����C�#�
7�\l6^V��ppR��obYjJ��~eԝ���N&rj�9��K����z��;��~8N{V2}h]�d^R~��+>'E�S�����+��t՜b�:��C.�Dꙩ�)st�s{$;"@M�;=1�tF���#��nK��Ty����ppa���V�����s����=��v]p+}ೃ��G�� ��Dp���3�{&#�\(�}�s�g����aH�C����&/Z�ƺ�#0�h�J"���C����G[e?�~�r�\VY��WΡ��V;'�*��1£���W,C�%���lm�������j�%Dl'+pO�#��i�*ʳ�JЊM��^�Q�S�jl �u�vޥh �kc�h�)��"�p��Ժ��ǁ�(W� 7c�e>c�G��Rd��c�D��_D4�?/&��=��O�Ѧ��(��)5-B�[�'cz��}�<�T�V���Z�8qB0�����O�=&��"	�.�gަ�T�ퟦ-�h��4h ����.���)t���g4��p�?ya��/�VZd���v�D��1s|q���߮�f���S.��^!��օ/�L��Lω�U�����J*@�dWjQ����o �[��Ɔ)�[�s�]n',�/DA�^ڛ4�ܛ^s�ХC�'o:dPA$S:F�C'P9Q&g��E?^�aO$���)������Ni�>'����Cb(�D�s.7���c#E��� gI�h���?"��	E��0N&)���<�
��7�H!��`rQc?g/?d��t;�C_a���Wª�c/��_�� pR[�v�`�,�jj�,[#��Hɫ��	~:�>���!^���Q����ԃN��"#��`5m�<���D��
����F�22�y���zcu�Ot�V~7���P� YJ��qqb(��ܯ|T��������f��M�ܰ��N8P|�"�~���W�S{`���MK���ks�Q&����m�֯�2!�����w��𸰑�F��xO��G)z-�vE���C��&T5,{܂}gC�=>���Ǭ�.�X���av޶�z_!�l6r��������3�E�&��!뷄wߢ��f� &��������������2�52�Of�|\����4/J��[�-a� ���_��#�^����֝�ս��9j�*=�m;a��g	�`�J!�r�*84)/�CܓFn��C{7���bd�6e����)�����t~L��d�r�
,�$J(�3	&f�>}��`��J���mD1��u���	W�G�1�> ��)ݒ���$?|OE��C�v�I�iZ��lͱ<ѧ��R�d7m*�@�l�H��u���f��3�����5R�8��U��z� �U�X9��ϐ�?aD�9�����k�v���nX�t9�_���`K��i��4�����Na�͕����xz�ZO�~t��Cp�V�
�rtH=w��l������/���4l]�ߜMg���-��+�7�-RA0�~�y7�{
��D����*ގ�������R����/�-cC���^F���j�a����oaé$I#+��*��.�̑��T�Lp;�b�%i�A꺱7�Y�zͪ��w��B��Օ��u�V�&T9��0��z�L}���������7Z���1�s��#�ð^�$����'�|q �58c+�e}?Q�8ʹ�}�v��LJ�%�+��މ:���c��K��J��5���ےS��xг��Z�P�!�Y�X�Z�^d��!�I��<P��0mlN�Ѵ�GRx���J1��ծ��B�z�s�(ct�
�:툜U�|�|���Bֽ۸ec���y��p�Q�q�	r��i�qv�H��D=Ѩ�x��م��u� Ȇ�Υe�T�Z��dT|]�J�_�j�1���#˸��!�;�?V}�BMNEG@N|���9��Oڢо���01�����WI�Q>��_�6֓'�κP�7����y�I##�N#�m�j���U������:RY�̴n=�$�O^SzO�C�:K�7�n2H�;��a �*�т�� #s��.�@�')&� �����9z8cw���,�Dn�;�]iT�����!���D�Ʌ��E�|�N����,�qg�#3ٿ�y�v�<-��4�,��z�Q*թ����q�5Zr��ݡ;:xl�a������x��*�PFP5��+ c��+�{xȽ$�o,�s�{�А���������ȄI�WץH���5���
��TC�ϑÉ����1ҥi��n��
�P,��5S�h�] <�sˀ��j�˓�Ŭ�!1	m����5��`������A��%�Eig�����%�T联d�����9�󏒑^2-P�ns���˧�:�jA|r>�bB�P��(l5�LYvԁ�um��	�{w�8R��,a�"���P\��&|�`J(众��JC�2���#�3wCWU��k��G�m��8����[���Ul��7�xnF�$�S�g�f>���,3����y*Y���љ~��g�r:��-��n���gqd*�{��hr@����Е>I=q�H���a�~��tp��H)��s# �ŕ��Xv�}�3�y�6b@�����F�Kq�\�N��d!Q���'sU����R�B�-�ES/L����8��"��	�7�##0"��O����j�5�8�w�ש��<�#�akK���bcZ��WFg���oӜרo�
�:�*`�`���u��&N�8�XRݳ$a#�����p�+m��k����y`6�rY���<n��Hf88|W֤-U=�ݶ�թ��ʼ�����}~8�W&����R�H��rVb�-�ހиM��h�Ӓ*����V`�� �`�׻���5���6#�zڐ|=㔒=�f��6�w�/�m*�i�a��.��k��Ny�T�m�MI���+�.�s=��0�@�./�Q��Θ��G����|���}�.�m�5p�vfa˪����|D���2���qݙ�Ȯ#倵���5H.���nG D�驨�%Ҧ:sj�c���G�8�0�Mr�H
���eu�]y,Oߗ��J���I�b�gSF��R�>V8r}��&Պ.�n��ENa�_�M�8����#kQ�-����C��\-�ܜ��$���m���Á7sw
�]�?~:�À��S���n��u{�䝯괹Ȳ��8`���7$g �}j�W���YG�k^�(�H @�"�}�5�8���
�'G�7`�$��U�X	� mW��	'�M��UBw��,%�GҬUa�9R$�R�£�O7����WN�BU�u�B E_ e�W��*v�]A6�\��p彣aj�k�V�.-`d'�#��Yb�5;� z�^锱:7��h��&!wS(nܤ�����3�����G�w9��� �����^S�������3��p�����S�!���m7�������4�ux?�e�"�d`3�~��͟��P�����h�R��/vWP{f�:�5����$�w��#�2��w��'�0߳n�L��w�ODiT�:
t�y�:���?7�m��=���Fc��=�)i�L���'M{v�C�5V�mn׉nB��F��k�\���f���������|�@)�V�c��[���$�#}�;@wB6 . �/�t=8�?�j�.��%��J�gc$�2.ʜ���<�+Nd��Quv�۰���; [>���,6|�	��9���.����*�y��L���=n�q�Ǿ]&��.[ ������d7����I�q�'�!�bV /k*���a�\bY����J̧�N�^��E��x��ٳ��#a-���t��,�r�=3�n��#�;	�@��M!@e��U+ �]��Ys�Wٛ(��߼h��7-�O+E�g�S��/#�f���{y�T�_�6�4�Z>;�e�dT/�"*�=e�=����x����#��]%} �EK�Oʮ��PG����X�.j�2�j�UW������*�]2�sZz�^�=X�_�τZJ�)�j�R����e��_,�xD.o����ޘh.,����E$S;�#Q���^�f �hE�keĮ3g�V�l����<֯�}i\�m�*�)R��p��8,��� [-:�vm>U�d@��֜�[=:�ŴՐſ��2�N��u��?k�����ik�n5�`�K��(ԣ[�ĳN�8����e�� Д_':}vm@���O�xH��}���� ���L��$Bs^u5�C�%Y[���Ox����׫Җ4��炏�*��ʹ�Zs�Ƹ�X��o���l������g�ѹ�ٔ������c�5�{E�W��#(GN�y�n��g��L� �m�����	�����'�ph����?&���m���[��a��9�!<w�F�&����a}����t/6n����y��)������Yhf�e�}��U�?���E�a!'F�{?W$r��t!�{lB�HX=&d�У���w)e%倯��{���R!7�uu�����c�&�D-�,���s�� tpaܲ�l9�-�M����׀!P5�$��t�c$ȡ��Y�-���܀Zd�o�Z�lN"s�څ�9x/k{�b����hEr�6v:m�r`�S���=ωv!?���VCI,�X��76���<SG��X����='���s�Q�g�OT�y��5w�Z�kW���;�3�q�J�_����S��P�5�x�v{~�L�h�����ap�R��p��ѩ��E*��ueMC6DqϹ ��k��\����i�ˈD>F�]��a�#�e��)�.�p���?vtg����ZAl����7�u?68I1�2j�i�.,��r�t�:0�-�v[�C<o�¬ =`5of-��P�O3h-�K#r�io2>��x���|
F�����}�Is��
 �����'����(j
펇xV5ܠ�I?A�R�	����79�%	�38y���Cju��[���k�]�+�����C��43K
|��W3Z|����"���0�<4�Ǉu�$���U�+V=�En��I��sz1�\؞�e����E�Q"�0���E�y"��a�೦. OA���尌;�'��^��ixHa���?-h�	#�u�I;�ybÜ�[«'p3<2��'�9����߹aƶ�SG���:�v��ܟ�&鄤��*	xAFx�y�5#lԵ�K��P�K����|�2\���(�'mK��t�"�f�欈'[�O��]��W�c_��O���b����"_�D��^ X!��n�b�FL��i�B�M�!���
��?$#\����%W �\�3��ou�g�����1�S+�\���_��bKK_�ڞ7~K�ni��H�3�wA�����
��
Zb�xL<�d��%5&�*��h�v�����6�[��k�3��boNF�ג��"-�%q4om֮
0�`h-p}��ږ�Y��*�&�0ݚ�]���]�	�w`��OӦ�$~�e5���`p1�b�z��Ӧa�yе��s:��B�F�!��F��xy����'�V�\
�(�Z�N@ʚ�Ԍ��ז[̑KH���6�H^�2U�k�����$��׏�K�r�}�v�B�鈿'/�=�f+)��T�B�P��u�H�Z��=ElQ��HRf0�:�}�~u�'߀�*��%��d��ׇ��t�t�.���L��y�
I��3�^c	�Ǚ�xy;=5Y�F���B���mr򣒌C5}��F��<��A��h��}ƣ�B�8����;�Α�gy-�,����>Ť�X�IN���8��u�d�86_L�q�������9����ŖU>��G�jK�����|{u���_��g{�f��;��=!����|NZ1�e�o��pDg�*���]s�����^g����.�H]P��ܫ����*�?��0 1眞�	� `��Ղ��o]�9�����#N����q��DG�5�;���X��I���3ߏ�*��]�Т�HY�F$oU�ȥ���x�z�m'�#��X�[�f�`.�i.0�L}�0��>,�v�q��@��ױ�g7]�V�`�,��h��n
�p�{�����Ġ�o)X�E�{>����m�)pQp;�[:���8�<a�Vivq�}��x�cXi'|G�(]��\�kQ�E4c�*�v�l[��QMbwV�L(h0 v� v�pa�&Up�\��Μ��^�С�@�{{r��0�r䚨�����Z���E��50oa5��6�;����nT�ǘ�����J�S��z����w�>=�k�<H�=*bs��C�(I���ח������6�@�XQ8ڍ�i��9F$��pp�Q�*P���_��=u@5zo�3��2��F	S`�^�>]���U|���[\�Pѐ�xl��-�T�)�WzT�+�
'��n�������z䷡���&j�Q��2Nw����|�k�[�G/�=�Qj������h�G���%��޺w��Ƒb�yS5�����m�贸�]'��E���l�t�d]즭�|}�m3�<�+D��D e�{�ݴ�]<� �B��@X�kМ��]/�T��oܨ�g�@���|S���L������J�4��!L��{!t79�Ƹ��}OǓƬ������O��Y$":�b �w�V����
&)�R�Jp�1�����T�6����U�3;�c:%�����$eV�7Gɻ/����-k��n���qR�]T"-B!̬@Ͳ9�,������X�ۮ�2hX"���6��=U��5���mI�� ,~x3wIV��Q�T���n����%��1_��WΠ�DC�;.���9�vi�����d9�H�+�b�TA���j��X~����1��>v<�%�����9]-g=����j�$�Q�y:�_0a|�8�떚����lw��]��܉�C��jG��5�Ql׿X��D���z�n}�Ԙ�6�E}��qV��_�`^���������]s�j�?r�z`���Kq&�u�
0��ZTZ�lV	Z��ua�fp١�գg����@n���)c5��%b��捋��u�E��s��.�C� -q��@+aBĲ�>����x���O��#nx�1�s���"��t�S2�wS��B���1J�Nx�g$�.���M�O��w�ʑ�W'�nT|1H)�F�̧`���O�L{bά���)�����%�giץ!g��7���*����=8[O���Ϳ�q�!'��eH�P�y��E�;�\5�c�s�]���:҂=����S�w���
D����}B��ڱ��^D��e}�_�h��#��0x�����3��{kx�kq^� Ս9]=��-:e�38��aa�\�|?��j�Gp.)/z�,���b�o���SF��y�s�5j#�a���G�����F�HcU>©6z���� n_�SU�hX�/��_��b:Yg�0�3M?.���7��H�~��Ol>Uk(�R3goj�Q������8¬����O�-n9���<8�42)
��#�0Kh&����8�I�v�_��\���슃 +{;�#��Xn�h� �P�}8���
.�2jN�oe���h����=�ďrv�qd�aS?`��|�7�~��`���}�M��H=���u�����c��-��?a�b����u�5�A� ��0�����r��ml�	'�I���|f�B��x���������MB	4�{��չ�Y����6��Ե=��`Mh2Y���XoD]��ڹG�Q|p�y�G���M�oWgy�����,�U��f\C]*� Ŕ���@�"��sm���[���o��Y,���6<yl�����WmQ���ZY���U��U����<� /��񆹍l�{�$ݝ����!�CO�~�?����]��4$��,�66�n̄�|P�wv��8�-/T�� d�S;���`�؎�Z��XP�ŵ�t���B�N&�UZ��<ARX!�{������H|��∗qo�wĮw���9�X�������E��܃Ȉ��kW G����L�ܺ�v�
Q���
�TF���`DJ���P83�a���7�V8��Y���"��#(G\4&<��82Q���; I�C5$�e��߳����-������#k�t�7�^Yo�� F"���5#��ƽ�f��fgY乻�*�dM����x���C�RGD��7M����\!���D>�p9�l��k:q�,����C�C��4�-��#���C�!,E��Jv����F��Q��,����	n!y�9�z'3,��tl1U/���i�>1�c7�))�t'�R���p��Y��oSBw�|"�s�nZ~��i���:D;H]�d0%M�w#�'Z��4���&�C0��Z�^uO*!���PB�k�6�wR�i<��O/=�N�/<h:�O��;{�₂����ܛ��4�m��}
�_�Z���~��>����)PI�S�t:"=Q��p��������lo7�Υː���]+h�F8b�g�-}Y�'A-/��=�<� �������A0�g���ɐ��!#ś���qͥ�4�e�Z��v"��F/2�����L�4����P�GV �������!w[�@*�an[C쿽�L�#M��?n����|�'����]��x������Ϛ�����3>f��$0���3e���4� w�Z�w�\G׵�oE�ߞH�)��Ouֆ=�Im���s4�}�c2C1��f����L��ڜQ�8n��|�v@�Bf/Z��/�<�8����M�F�33������>P!��Ew�� �e���� P"�eAd�K����IDx�{X�ԒE$�����M��+}����[�>��ԉR+-_"���N��p}�R}��v�ƊQ���K���$�*�p�M����wC��|�U�ԓЮ.!�O�1�D[��~����m�ze���O���*�
���_�J�T���y#c_�t�Q�{cB�3�z����L�yK���#��!�@ok(a�i�Z$�sj����0�ǴJN���k���=���^�U�m·�`�.�37���m��B�qq\�f�1Oc9��\rF������Ұ�Nr��n�����_6����f��ɦ�m��m�ƨ��i���2� nI/���7�T��	𭣃�?/L�O���ÇsI�I��GT)sH?�I��=Jz�y������}�[	2`��M	V�bT�4��e�U~�ް�&N�I���� �_�,d�z{gy.B�T$\k�燽;���ď�����[A�\�t,?���#��p=��ǉl	gZ�,l���ɹ`A�h�L�;
C�Z�e�C��C(�Ӂ�����;5[L���$��<z���^��e0��ŝPU!:��iTOp�(��_��� z�m/v���<W�BM~�D2>YK{A��`v���Dʤ�G��>%���p�!A����4d��G%�()�V�Ό�\�f��VP+�&�n��xxߛ���'�	���4�թ��)�����Hf��JD�J�2�h�����9�6��I����>���ߏ�9�c��2����M��i
j��c2��Ud�XCϿ�_L"g����!+�@	��9��ʯ_2�����¬p?��>�Xc�GO������@`2���S��H,���=��Ʀ�@��4���K�-�C�ͮ��]�Ȋ�م�qwStI�2#��"��������oė�H�ko���e�D�:j����&�8�����ME1h/�w
�?�$�L_/^?u�s}�u���dڛ޶�Y0�r�mE�/�~��:�9�V$�ea�n�'���g$EQM �B�3D{���g�H,c�M]-��;�~\�#�F?����p�U��'�M�`"�l��ġ���S���4�<P?_��B���~ְ�0��H�#�z�ہ�׫�AT�E f�Yּ�i\�#
�5l�$��-t�)7�#)�Kb��#���|
:�
^��A� >@A*H�Eo����U���;np�EUhB;��.�4�c6��JdUv��;�lWǜA�9��3-.[`T�@'�6�"��2#�Hf���9