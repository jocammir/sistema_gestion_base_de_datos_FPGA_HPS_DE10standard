��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����{hi��7	G�����|��4/���YEs��Q��H�9e���ϒ��(��t�.�?�ѩ<�Փ�<�Evj���T�����B�ݰ7� ػ�3��p�����D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�D�c�;��ЄUO���?�G�����d����w��ܳ�5�@��=T�σCFV���C	��r���o��[��C)r�|Ϸ�A�4���b�� 8v$(�����vSw�D˔��I
!���Ӟ'8nJ]�A�q�Z�qK�m�q������ہ!.f����C������n������NPR�[���cF�]֏�U��_����ÍiD)l�h7�UƎ��a% \6���Q�7�������&��{�W��WsF�8�z���.(>.���|r1��51�4�U��1���(:(L�'�6���'	��ZS|��u_@�'D��T�Agu�t���Me����i��h�M��bU�_¯W��N+3� �0�W�έ��A�0�|{���&VT���
�+���I�ں6�� �K�<�k�tZ�	_T��Z,�ֆ�8�*�c����$�N2��+uɤe�c%D~�~~��1�ל�	���U�u��Ӣ�#˅���Kwx�
�V*0��újT)_+��Ua��.!\W�����&L�EX����Q��,��2�>�e6�7KZ�I�HlTl񻂑�x���l*vz�$�qR�r�5���O	��SΊ���޲�t	E\�e.�0�~2iw��Gw��b�һ�XT�{�n���$s>�v���5��Of��t&^AY�k�m;/Y4��K�#��h�Ӻ�.��[8�xֈ���">�V�0���^��t��}�	)�"�M�;�f�m9ҍ���/c�<b3g'��9��;pl!�ܩJ)ݴ؍���/�~d��<��r���A}�����u�n���?ˮ�;�
�I�|�r4����F�������)�{� a��J�*�
��봂bV���Q�*$,I�U3�`�q����R�:�a����,4u���^�*�2kxT7�"L���ľ����%e�&̫Q��6�@��4��h-� �;���8'5S�nl��/`hW��8�C� ��.�&l2[?����c1��c��� ˱���-���wN��3�aA�f�	� �d����cP�]$�Y�4��%g30���K�	��0��m ��،�z��4��XϏiɶC�1\&9ey�X۬c�E���Cp�S|�#po$������9mǍ��#�7Am���3�����`�ȁ�>���Z�ܦ�j�P�(�Cv���+ %�^��E���9�nL��ם��\	��ݕ�گ�����e:j�t�AN�;Қ�$_<��,�,�2G���Ͳы�[͸��A�쒟��G��:/đ3�#/+
%��6#)��B"�����6C�zezg��1������!I��o�)uE������R+��\�N�[����%���ԅ\B�0c�$��_�R�J2�w	`�R�U�%MZpƻ+9� �D��8A�m��;_�N��S.���y� %N놅��h)N �9^�[1�9'���k���ܤNVU�H�	Tg�J�nt3G�؁t��2���O�d���d�0�=#�l�e�w錍���&<F�����|�	G�G0���f�6��Q�(g�ZJ���ϗ �c6�-Z�7{|X],<8���l��5օ_mY�w�y;�cd�{�m%���U.=D�A�Gd��>�I��x�l��Y\ ��H@�z�r�Uo0�bDuM�0 �i�ˍK�m���wV���g�PT��Z(����-IQ��>2)��D�%F�<P+k�E ~M	�7�x����wBH����£�pk:ue�q;�>B�6�އ��S���i.!�foJ7���p'����Vm���y��ދ�I��^����Ƣ־��.!��  I�/�f�R����	��H^m@^����"�
i��v^kXlҟ���	r��<�J��Z���K���S6��"���3���ee����@�At�ư�~j����|*���M���v���A�U���H��zdHH,�#�7m0�-������"��q���&`nI��qڸ!�A�r6C�=L��8B ��[�>=p��¥��8_�A8��½�R��*en'F���z�ڟҀ�,�o�#��Q��S&&�4%����L�A\���V���n��Ǩ��|d �{]X]RMњ�n� ��[�ѳ�f�TpRݭ�Ө�+l;�x<u$�K$���׋��a-e#e��9_�����`	���j1J�*���ȏ�J�=�.e�pzD�n�Ei�Bύ��M��Q'��Z����� �s�oA���8���7h�R��>T�A�mGmM�)a=�=^�{��`1��2:*|���^����\qv8��4�2Z�w=(]��AE����;�@%i	HYx95hǴȄ��v�]y|�/T�^�J�<���U!�.阖�lmG��$�m���7,�J9���� ��O���]�	��Ј��AFg�;���^�E�c��-2l�~C��0�yI�~)��`�T��M��4Oz�AA��4�\ۃ&�����d&�yH�2w�uYM8�
�H<;M�O�����Kj����.>ֶ��XHf�N���b�@7��<B޳�3�MFXE�.zk)r�\P���W(|��ΐ6���e�E*��W�Sҧ��^�p����uA������6ČM�G����p�f`�S��@���=���{?IF�l��ՊS�#]���H������WW��x��g����ڟG����_��}Y���b��\~�8^ۆ�it�U�{��7<i�sU��%��>�����E��]'ؼF!�\�D��4�}/����i���	��I�z�N�ӊ���y6�$�#GL�J2��7 �~��p����l���c�9�'��Q�Wr�r���I� �z��ܮ1 ��� ��}{C(/���1���YQ�:h�ߪ[-�8��*���d٪&�Ȉ\�s6:��_���PLR)���3ͫ�;IT
{��9It_.եԃV$n'4�6�%_O��+�侌4��l�og�K�5�.�׮J���vq���N��懾h��A�i��o�����(v�h\;E���a
����6��K�Լ;��F�qp�<*6'ꍣ�)�;"]/W����������ԅW؜A��Sm��0�-��͹W]�����/��S�ghm�My6�������N����
�Dy6rA�FǢ����*+�91)b�2��l|� ����Č������K�\�}Ez��n\�Z�1�� f��ՙ�NV���"1�/@?��*����<�
��ʔB��pۥ��
%".��(�D��ȹ��*d��]�A����q�+?�X�N��L7�a�A�OO��ک�|���WN�S�$u�IFh�J�Z�I+XI/9�7dp�j.N��c�P�	Pk�4�Tى�}��Gb�P)~�:}��\?9-�t>�j5�4RGv�_�EՈS>)����^n�K=�[K5�o�|��ێw<�¡��ˊb�B{�������L	�L(~�B�68=�z�*9��)�瀕�Zd���=\�y� ,-,�&+��b��k��>sT��#��=�U�mg_��G�
C4��[���2�;����4�I�,�9N�mT�5Hz�\�=�u��X6�LQ �B���-�f�t�UZ�O���@}�	ڽ寜d\���W�Ɓ��J��b}wU |�>��G^i,!��_p��� ��3���s�\<�}����U"z�$䐢0��Bɳ�������=Y��-j7��iq9p�����5h����!,�-H�����c��+��am�>����X8C~�?�&�$�.R�Y���Cc�I�9���<���/�~�º�er�X�I������7�r5}��o�*[���{�d��'ZH�A�eki�
5��JU�=���M�2;!�2yw���L��-����(00�n--�x�2����۞���s[��}�Fl��[�7��32�*	$Ʒ��A�`���C�'�ag��y�;Γ���CKj�vU�ro^�&z�N3��'7����aHՏ��Q�J})j����ǄF�%ڸ�hfz��Ȗ˞(�f�h�b;�(�h��B�k:�j��D҇f�UU��c[�5�-��HG�y��<P��s>�"+C%�p"�d����W��l���_�`�;͐a}��O>b!�+h����d5E�>c	Ej�x�HMk��kۛ��q���5�`_�YO4BZ��^\N$p
0���bv8B2y���l}*w�\��}j��VQ�#��W;��yp�	Q;準P`-7�m��a(:0��#?Pyĺ��0Z�)��qo#1���;�VF_��Y��k�h��_'<�J��Q*-��N��fa.,�Ë�qኜ#��~������U��o�h�c�'C�o9s⒦
v��7)H��v�U��p�c#.~ �yh�As��ZRHg"y)��!�	w����M8����TC8s��?]d�oJ?����z��x�e�͈�����C�L0O��<"���7	���J-@Gh�3x6�O�%���ś̅N=���)�b��c]�V�ܿVsh!f����f��I�������vF\�(+nb��ʭB	�y�^%o\r����v��E����E�f�x)ws���hd���a�؜R#���F�?� :�%&wH��3%(&@��D�ߗ-�%cc�΂k	��},F�a��/O��{����:=��(ŸÌ�8�la%�+v6n6����^g�˚@Bg;{��Q;	����Fr[�w�
)1�������Q��oI��0#�V�]�,f���
#��/�b6��"3zQ�!�.G:r����}��G[����W�C�L/Xs�|�r�k*�ŋG�*JhQ��H�Ǩ��w�|�[n��רH�.K�"Ad�>�ޮ��1�i�4>�Ö	䧏4M�)c�"ߙkkz~.�`�4f�����8�����Ws��T�#�K���y�D�����]t0�Ῡ.ȏ����b��*7���g꺝��o18�_I���\�2k�
QwL�ȿ��mjS_�#�]�#In��~�3������#��Sg	���,�=d��M�1�,�T���|�6Ah��#n�5�Qr�e>F���!�+U�E��(�	U��WA���B����\Û�ږ���=�H����z���Ԯ�bA�n)����Qr0Y30�w)��C�O9��`g��f�#��O`5³o�C�-CU�|��9ц��j\�=���B�f:cڱw�]�������Mׇ���Ŝ2H��/_�c�Z���4�q��p�=Y�%{�亅gKbv8B����I�( ���T.?B����7�|�5�q�g�H	�	�e{6�Y���H4X�g�\�c�-X�����O�[���ux��l��������ש�����# ?;)��i�<��#�Z;
�����\������9��`n�l\���������F8*\��7�Z�=��i>ֻ�ʶϨ�I��ҽ����?�w5�� d���s"�X{�Nև�жVֻ�`@bTxW���q�X$��)�r;E&	�Y���ޘ�Cr�FR�xL�l�:����M���[M���� \�(��?u͡��"�+�8V��2jNr�,G'M�B��s��Q��º�أ�@@���B�/B�ڻ��	Ϧ�WpM!���r[���Z�.�ʀQ�ȬOK��#�x4��@�bj3n ��z����Zި�D�r�L�/#m�e\�5(#�ā4gc���7<sᲫ����(�g`��������7K�ʹC ��\}�35���C{���ȗL�ˌ��CA���]�.��,���fJE]�A�6�JC.LT�_��̅W��[j]U^��c-��O��!���"�Ks\K��v�1*ip���`f*���OgYB��~�"
+��(�(��1 ��~������Њ[6i8S�����ÁCy6x'���EHAE���]�G-��b�����1:(��&f݁�'4��VF悁���8R�o�4��f�(3aa���28]y�S2^��x�x���������}ϔ����mH�@!��%�1�m�v��o"�&�nBE��w�_�S�ox���_����F��e�5KB�7b�zEKYp���Q66T�z$���9�5+���md�?��ֵ%�>��mѻ��N�S^��|�a�Kg�A��������BÛ�S�
k�[K��y�h�{��ۓ@�*��Q���,TLҎmT���f�t)��������h�{C��14�|�<.��~�5"�
�}*��3����/A_�-��vEXUn{?� z�ݰ֫�"o2���"AE�$1�_�L�`
�	����f�X���]Z`�^+9@˹y��0p9�y��d�9j�3�<��J�%K����|  ����_$�M�����,1W�(��Q�:�ؐO�2��(�IL"}�.�˖�S�{�Q�`r��M�(�ё� ���0g�M�$f�W"���D�᎟<I�OTox |3��,c�(��q٩�`�B�¤&Ru�����;i��H����j�խl�ư�U�"i�?1]}��ڪ|�c��`8��Q�o/2���o�ð(�������EA�M��\����X.�Mƌ����ܸ^}y��� &{q|�i_xT�A/�n_E QP�K~�,�@{�嵔���P�g����#I_��������]��ls?��b������z����ގ��ǐ��8k6-�s�-]]��8g��߸b��Qhi����$��6;����ʅ�qC�J+HJ�U���z��������L��\��cڝx�ݑ�*[��=O�Sn����/�V�5��) �!����(2iX�g���Ubϕ/sU����R�z2<Ӧ�� �q$rMz�d�ː�0����c�Mp1k'��!�٪�����E�A�k���t�� ��_d2�P�2�Y_�ML&���,u�`�V�Í��+ 5����!V=�� ��%����2WW5'�쭸H�e��}�zQo'NP�>�Fg���X**|����b��xW�3pp$�O#�Yؒ���Q�|'J���=�\`�Sy���]�#Zd�|�jX���i���&��󅪹����U�'�W���S-�KNk��\��$A͕���;��������xv1�A�|2�0�9�Վf�h��|�C�&� �o�RZ
h<�y�s�d�cͶ}�8T�p�^�� ���.���gj}�s /�|`�J!ip�['�>��yǩ��Y�H��xp���a�Tv��	����:[6v�ϴ�<�!�p;7�#�hpt���g�)z9�,��43�	�	��¬��~dw-�o���`3�p�f7݅���s{�iM]I��8m��l���X+��蠦I�;!hd�~b��}h��;�f�y	a��g��-/�F�A�ά�#�3����$�����r�𵹾��}5��H��ԽG�P���kQ�����J���Z}���ŏ��ZaD
�&D��#ny�&[��րN���d��Q�A����������yGng�͈�*����:{Նg�kH�bk��s2��K&P���m��!j�M�QM�x�2�'m�y�k��{�,Pv�?9��#��,���POT%��DFiձ��9��!dTu�^�t�#���9s*�����$���5�S�컊�O$N3���X�dK�vJE�?��}��\#�L2?gЕ����S��B��o(�kE<O�bEy��	�+Vw��{��^G�m���dT.�=2�!�%kUm�?�r �Ǿ�eԄ�#	ʈi����F��4����ƺ[��*��H������C�i���"��I�.�R�`�1dG��A�թmՈ,Ǫ��R�drӾ��]�x��XU�B���r~X�����7	_��ҷ5ѓ����Je�`���M�~q��"k�����(�dͺ���� y�hS׌ǿ|~Oi�����uB�>�ҁ~P2�aՇ��ȥ- >
p:�|���J���eP�d"�<���YA#��Nw�	�O��:3� �0>i���1_c�,�ܛX=��������dd��~:	�-�~�g�yåj�>բ�q�)rѥb�r�L�<�V��m����T��M����C=��|r�Ǌq2ف�b�0�Gs3�f�h���\�<�#�� m���y*���+���`m)�{=�,#`�$g�;f�,��1���'7��L�u8�����:Z`��L�d2-��uع���3̙�-1�H�.�v��0>��VŮ�Yh~3r~h�n\��/m�Qgqt�ͯ}\/�|�/L���쏻Y�c8wt�~���@�����]�(�C���&���i?~��iPV��_������K�w��αw�+���+h�e�ё�Պ��`���ɩ����կ��E�:��NC��`x 	�&��0xE�Nb,���q��C,�?��	%1�J���j�I��.8�N�4\�dlrhL��i賶PS��֫=����R�eC��֞7nm_t��������foF:�d�|ݪxlbe^��>�]���fI?�
.�`��뱴<�}@��%m��I�1��'6q�F#�f_2��H��|���S�����ÙũE��С^� ����V�{'
xH�ӝ�H����{��Ŭr��/�Z�$R��ǯ�0�8,W�
��n}����bI��X� �Z�m��:��_-t��<���e�M����s��{z��$â{��WaH}��\øx�zUJ�0�ۂs}}��;b��3v3x�ҥ����_s�����b�'��HmKmMd�����`;��fT����B�<���4�E��ї�ɤ�)����Ŝ&����f�pDG����ӘY�o���b�?Q�h�|7U��&��ڈ��N�1}d�9)�Ь�i޹O���|�V�v���"�c�]��\g"[Z�q@A�y?^U*s�}�H{��S
g\�MO��̅X�i�ޟ?|�pbu�py�������,0����>�dDgUli�z�?�/���G�tu���}��>+�3g�jp�w.�����0���4��5BP_�OE��(�H�S2�M㾫�ݺ\������\}�R��+E��� ��?c�QO�����`]���žx��am/�_���=��̢�|7U:�;(" *\��͑�@	K{�O.n(�xc&o�;	���^��5����Q�"���W��MY����I=D�����5w��z�����P����J� �tPn�]�?a��R��7 #63p�0�H�av� <�#iݎ?��=��aY��.���C��������>n�1Bh��@��j�_:P*�?<��%$ZU�v���,/�vbAeR'�e��W��a|}�^��w��fu�"�&���;n�����Zo���r���s$^�B��m�y8I�+����̹P��	4(�f��M���1\��t�(${s����[��k���t{��j�d���ơ�/�V_�c���e
�,Q!�y�{^�Is�ő���J���괔x"�
eɮ  ŉB2�,ʯA�砪���q������	0��L<\�,����4��s�ux�do���"�-�L�֩�l�������7�m�2���#?QXV����_X�7��;�B�b@3E�4k&c��y1e���� ��C�m����#Me)��Lh���X�.�sCk��|������$b!�?��8���A�Л�޽^��jz���<�C��!��&��m�EՃ��١3��7Q`4�>�����?;�yA֡�m0)JT�Ea�l�<����E�����b,W�h����LSښO6�4΢�K�,�_'���t��&�)�B m #���VUL- fGZ�z�[Y������!b·����=�;��Ǹ�[&�s #�B�ޔ����{y��{��mu�I���ڼ2���?�w��i�T�Fl�d��pP�1`���~H͸�d��Q����"�F��/�c����Ց��i��r�(��^�z�8&tG�J�K]^iMm4�1b���L|�`
�5�xl����s�!W��$�M�h�Vh�< 
w�X�!kZ��7����a�ݨ�ɚ��-i�|���x��^K��P�1L�G
5���1���X�ǰ�'|?!{όT�-�1��c{�n�����3�7�)�'� ��o�f�\��&�O�~YR���y���GC���&4M�G�h��B߼�$��R���ܑ�e�*���)�����%Ȟ� cL�c7JI��_/bw>z����=,/���!$%*��j5F��Xc�����F�7΄��s/œ�t�I.�hwR�O��툟�1w
Ub���/���7�\c��s��_���;��|�M�G� ��b�A�LP��u��G p]��ྋi�U�L�U�t�n9��}��g�ОhE��+
����M�\ȑ�X�Z������u(.�%{8MC!�B='�-�W3r���[��yd�o���u�w͈
o���W�Qg�-������o<"�tGǮ�l���%�p(�
��IN`s[VV:%��2IUEyxm�qj��Md��5��c?� �����#LC�~K�	�^�$����C�4�Sl���Z˗�;8��\��SVN63�]��Fc�~�{���&|�0����7��F��aƖױ����!.�}gCo��t�/+8�F�T�K���X�!�g���qm:���ʳ"fm�鞺	U.�OF�����,� �"b���a�!���*;��t��r�lO�L��M8Ws�ٝ�P�!��ՇS��	{Ht}5�X�T�N�$����!I�n���*J���4a=�����]h�f܏�ڢ
䚣M�Xd���1�zA���Ur����_Ɂj��B^�4�d��*7$���;��4�=��.��>���X���IQRfh�g�R��tWR�N�rTB��Rz~\͸D�wm�qp��RDH�Nf�<rj�S׷�Q!{�W4I6��-U��QU&v9��r �' ���w��(L�";K������<��d��-��K�/� ��(�t��
��[�]�_��r���(w@�&��V���-1�XT�nմ�h^gn�DL���J���h��z���\cz�7�H��Z���.|����j%�o�HT!NpN�^*� ���p�M�����~=�T�=竮Yd�z�H>�X!��
/g�JM[zm3&D��uN#�aӠ��P�n��z���,����9�D ��Ľ~ׂ�&����d/<:c��np^���Q����c�H6�"�
��s6G�ľ`�Z����[���Vԗ�� ��/��8�_��۪
O��F�Y�f{v�\��n޳~"��R�B�}��cD�J2j��ҘD�Y0ٸH��C�Ċ��_`oM�N͒�!�'`�G�����OV�BK����(c��JTRq�� ��ߵ�]�8��ǩ�G�k�Iz�lE8���?F�}�����?�������0b�k��A�9[4�.kmׄ�8岌�f������xv��趿�.f$�N�@&R����x@^��nU!���S���?����K���g�}ݧMo ��u�~�������A�����,~��
��C����k=�����F(��ޛZ:]�;�ڐ�P�A�#�ab֌��u�E���Iߕ�ܱl�
�eB9@�QZ�\h��c̙��92l9��Rl�ҋ�m��H-������/��GwH�hr=*'/ڵ�l]�trv�����p��"L�3��@h:���d� KFP�([!%�8�X�c�M�(��<sݺ�1bB�Ez+w����n���t����d�����Jl�{��	���G��ּ
q&���`�X�9�����4ϐ�T �&�Q�/��6D�*�鉈�!��(Ur��r�EJ~,Y������kl��U7S�"=%�쳻g;�@������M����^u�o��P������<�5���Ԁ���J�Ns=�F����5%��K��O��1L�d��E2��"�`q������IP=� �W��餐�~θ�L�����.��sI���<\�����n�V
UW�l����rusB}�� �Uf+���V/翋��|Q�%C0{���(K;*?u�}5�V�=���v�[��P�3�D(���������n���A�B�S�k�ș3n0��/����B�l=^o���{�@�y��	�kg�m@,$�ܫk�i�V_��������ϲC|#H(IC����;���ɪm�=.50�(��z�#�jH��s����r�B%0#"g2��''F�W~餞*�M~҆��}2H۩|���30���en����C9��V'Lp^f'�@х\	���9��]��4x~��.��*ƆP_�R��tr�k��7\����녹ė��eC�ڲ�i��cS�����w��|�j�۔ʯC�\?� �{����D@��Z�zd1�W$�H�C_�t�S�u��2+7�
撎&���=_�X�������J���5%�\eM������:8�S�n��Q�D_��Sdc��/�l+�m���]g��ㅴ� N�!�ß�4�B|���yr��
k�f�+�;I�m:���Q��<^�[Ks�k�O��[��^�tdv�8�8jr��pPYmORF ��<�3h/p-���q(�htZ p�Z�dz�0���CLƢ3�����/$�W�T�T��` 'G'���¡"y;H�*��E<؜�MZ�	��=a�� {�@N��g_�$ս���yF�&n1���u�����|���\˛�ȮQ�i�uB�F4֐I��ǒ�uc��Mct鄍���4������p��_�ш�'�6�Me,��w1�Dj�$��B	��HD�fV��;Q4>�Y_ϩM�a콗l��?	9���'%���y(�2|Q��Q�_���=n�CsW���1&&�rp�l�T���ח�Ef�+J���� z>��!���j��'�ɦ!�fP���=fJc!�@�#��c?�5�+�}�/�p�u�q���>y%S�<�BD��oQEԱ_�G0��k�NU��~�fQ��(n
��@���`Ä:<���pգ'o)�� =Q�d��i�Q_�h�Ħ�B���=�Ϝ�bq�c�t3���B߆��~BoFڈ��+�4����f���k)u�Lz�K:f�� ��=g@E�6�?ra�'��3�H�^n���Z*�a�%kd�3o��Kf�wBN�f��^����_��v�]�%g���pK�@�v�:ڷ���� +�.گ��x0���~�Œշ`#ꕴ�6]�;-5��2��
�K��啥�!�+�;�n�6TZ*lrAA$Y�|9���v X��JpQ��i�h�]g&D�%��U%u�����!Jb�Z�I{�A�j���7u�<����It��|0��'�@��[0?c���xZ��˿��Y_:Q��7�F���w~�ݭ'��kY4'@�u� Z�S{c���yw̨����7��p�,o��t��`��&�m���;�sgd�5���A�e���X�.� �tT�2��v':ӈp�{�o>�}n��7���N�w
ba��/�N&*��O�1�k�:k��<��dz�����J��<Ram�S��6-|˗�9�ޥ]�5,�m��m�e"���:���}��dS)�f95��oaYW�J7ŀ�qS�5��W��� �X�~���#�P,h�"��x���ߖ.0
n�/����eظ_�)�i�,���j����l�,GF�ߪRA$w=b��͝#h�����mq�)�$��3T��	�I��A�kl����@��o������D�6�;Y��ҙ�m-�#�*S�I���|�i����j��4?BfN��9��+H��<�<�J�|����hXJЇgMҒ���5&}uQݍ�Nü��qA�H�.A�?��=�O�@[�[LBd-�)�xeCB�w*	TH�<e�1��Z��*L��NQ6f4|k�������k�n^O�ܽH�|�<Sy�����~W�k�H���-�թ�'�[9�[8G�Z<F�WpĦ�!+�h2��'	���0�^�&C��b������	��u��1��(�����Z]^�G��aF������y>:��l9�ٸOa�ũ:�f.��?8������kj��a�}a�kL{,m���ץ(hZ�^�W&���8��{��H�������k�9`�z��@vo����5���sd�L�D�:b�!2��&#ۣVD֙����޶���"���7�����\+�����y4E qԥ��=��Ӝ��"���.� /V�V�_��{�̫�8�:�k`ENi����/E��S1-D�X��5?F�F�Ϟ��4K�m�R 5��x�3�	�q,l#�ԁ����?����TD\�YA<��>�Ϥ6eއ^^;��T���`A9"A����O�x2����n��������5�=��H���#�&�&�d^7L�췳hio��zP�7b,i���H����AܨSuO��a�	�]�l�P���܀n�	q��9B��S�#:^0�'�F���^=�[�κ���[B��9Z�NmtT�FKEQ%K'#�GgEh;U�v%�O��9>4{q���_���^n�{�U�rT�p��E�g���շ������`���;Ќ��("��w�g"q�y
�T�;�&FN�����I~S���^G�4�L��{5��{���a��H�R�}�r~�L��}�K�C�J�Ē���'?[K��"#��;�К'W����n0��Xҕ5�uD
�Q<����5=��r���}�c&:�7�LΤ����}z}�-�e�!�"��٢[�i���7]A��)Kw�dƱ}��h��rc��5������5��!l�֚P��"m�(��}����x6�W������mv�h�0�	��:o���'홻����.&�g���k��I2�F�t?]O*f�ûztlx42�X�{����q4)(r(/�n8�0����*����	��Å�[\���iM|��nTǥ΋_1�QEl�g�s���S!�W���֝7lK�X?3��&G�	�����FH˯�:����0new̽��1)@�mJ��<�g�VD.X��.��c����GÞ_�0��iԖ��$���+}������ɸ�M�֪�ׯ�,��k���.u?r�����e�?AoP]Kv�{�AK^��u���>|�o���Ֆ�O�`w��C�`"�h�Y��HE�Nl�a����H�����w�I`�X�b ��h���-����ݨ��v������@r֧fA)�¡X�d������;�BV$���q([w�r��F��-Xv�F�X~�X���ߠ�����^��fh��)\9I.FaS�j�?��8���	-Mǐ�IS�7�̯xA�~QX��(�S ��z��<P���~�b�'��H�0VX_��3z���4��'����u�r� 8����\*<;�x��8%���m�q�QL��){W��U%�7Q��3S�(#��	�'�[i��ݵ'WhZr�&�ǹOF��	a��a�)@4!�(�]��ݯ��sR9h���$����}��������կ<��\w�a��e�"߃���m��hy�� ������dq�{���9W��E	'�M*��q-��9�����g�J\qa�au�iN�X�QŃ�G��9��,R�Ȳ!�]V���سl���@��<u�	 �C����]��@�"e�t�OB�)a�Z}���ʚW�8�ϧ,ZC�3�)نRs9�{:4&[�4������ ��'���r��^J�A ~�U���L�L�9c��S�
C�|v����9�`j>�[��>TA�X�?3�/t��#�f� �� '�!����y]_밼����I���/)"�C�I)��;�s�%��Bܿ��i��T�T����z�q�u�hz�(ް�����#}�u&�'�חQ�z����eׄOݜ�� $di!^&F������-y����I��$?;Nq�^"X�ŏ���,���Z��3Љm�����9c��b�7]����p[�hF����Z�,��ΰ�`<!���&���VTn~�8�u ��1.�-G�)�Sr�	$LR3F/x�b~D�đ^i]ۍ�A$����h�L���+R���f�)���}�F�% �e���%���S���N��Ǆ����C'Ǜc^�hg�CTC�X,��hBѓ��A��qz��F�=
��(�(�~�p��\���Ao������t�T���0�����,�?�퀸9���]5T���Ӂ���M�uF�0X�o���~5%l#)Jpk�N=N<��$:���v��"���O��Yr����`��댥��bRha�׭��Vqw9u��c��|k�Տ��sۙ��hM�Y�eeN��!�d�(b�ƺ{-�Gn� K��D�#�B���!p�2|�3W |�Ÿ�@Am0���	x�r�0rͬ6�੊�M��b���Y�qNQ)���!+gVq��L��:J�j��IM���B�Ē�O5!̰AB$}�T}��V�����`�V��Z���HBu�����c���9���Q�a��Y_�*�Sj��D����4-O#*p
���F���MS1{N֚��;&ٴ�������a�ΐ�@�%�Y"d9�h[�m�rO�0hټװ%ޠ����ys�A�À�'��g0D	0���@W����K�F~�x�T���,`�C�y17/�r���lK�y�X}\�-:��(��e( ͟q-���೒FwD��;aڰ��]��O9���%XY��"��H�g���߹�H��]F
%#fӺ����帗��Y�n[�g��V���Y$�Ó�Y+�]���Zq;{ܾ$Y���u�&a%r���< �F�^Y(���~�G�!#M�nb���"�2���(�m�}���`��ep�a�X���*�4�<��O�#Q�%�XaR9�X��#�rU��e��R�.�Daxq"��vv}��tz\�㫇8�N5�9�Mn�ﳹ�LkV�� m��4Z�������H&���6*��De�K�yk� ��~��V�u����#���TV�s�8S��>N��z��V>m.�s��UK��IV���E�T��yh���DR�FUü�=���9J?կ�?QƹepQ	8H�h��E��K�\-�o�^v���b�~V���D�'�/Ϊ�ߴA�BL�:r0�w�D,�Kv`���c��,��@�sb�����Y��LC^���=�@T&���X�b"�=[�M0���J�r�v���U��xL��Ȉmn�	���EYU�Qfܠ܆8tx�(�\�^�_�;.��HY|��J�nH�J�;��[�)���3'���pk��h��U��'�0��BR�>Z��	�
�q l�PӐ���RF��Y5{cZ�����˟aL\��@��@��rCkzE*��K��������|Z�G��(LT�k!v_K/L&�dU�r�
�(�G;~W������E���eJ����]�ؘ��*���m�쭿|�q.���cs��X�-��\똞��!L�ԻO��eh�dO�^S�FS|"�W�1�WĔ�]!���}�a��R��I���&�H��� �bZu�R!R�F'Q�=tI�30��5_a��n�ɸsj7w2�s�T��#�*�7	ab���($�(���a�zTVwT:T�1I��l��8�*����N��v�{���3��A1�	,�RZc}���Ô�<�O��yp�t�E<4�?z�	č��"��n\���εCcÝ�=�����}�|Fd�
`���X�:`�w�����6���߿��!�:���A�1b��\�L��c���Ƥ�[V�U���c6eF�F`��^~����>
FTC�'����4��ݜ.��R�|��W�T�[�E�Ж7�pS�1nf<C�}n��k�dxYv�h�`��ŴA�,è=��x��|a��5Ax�v!��-�Ʌ%E �M�v�w`�!�2}3�O[R>XG������"�CL��	-y�j���k�|���l��X���&OuaKء��sj��48�fP6ؗ8ۊx���?"�~m ͐m�X�n�L7_
]�)Kǽd,�f,6;I���{Hn@h��t����PG��G�M;p�9����9�� ��0yom)�'�l�*����W(��`�u��0l��h<K�U9o,�V��߅48_	�#�[�����y�0��O��'�4�.v�v��w���aY$�U�����U&YO9�����-:%O�X��<|���q���k��M>ø���om$����0���A@��������z�[��X�[{���ڤ�o�o��N����l��z�����@���5�^���_���'GW�4g#��\໤[V�k���a���2i7iz�K�#�7*ETM�_m^ZU�^�#{�$�)�
�$<�(�ٔ��G4�UY�&���D���N ��^R!����y$���r^o��	}}���(nD���Z�1���~�B,/8�-B���乇 M�f�����@ȕu4%�ࡧ�پ�p��%_}|�K(=Q@��͉���>�9���2_��>�g�*d�/������vL�<}�.Ѷ�N��f���� ����ޜ���N�ʨ�� ��H�,����[xqv�@��+4,Mի}I�.�餺����ȹ"�E	�J�G�ő�(N��*�w����&����)��q��깛,��+Y ��d��/Qg';|Q�VjS�檴���?s[�Iï�y����Dd�� �.��*��f�Sc�s�4\����3mEH�%�P��u���?����C e킣�?˥�@�aP�;L�HxM�g�� ��7�Z�5ş ������:�##���X�n��FG�h8�����u\�Z���	�Sر`$V�.WUx׷#h��̧l�)���܍9�x�C�m��w��C��`w��]p;��KAɍ���0�p��.��,ew0�ا�П��HYL%F��ܦ������JAE�N~�.;����(���?DC����ˌib��)��]S�_�)�+S4^��rT��.k,�Y=�ϱ� r���IOn���gi������U`=q�����3���iƠ�֫T.<� d3տ��'�w!���v��$A��v�0RX
-x3��dt��&;r9����K ϡ��m���O�W#��O_3�is#i�'3�j�]����'�m� h���z��?���f�;�;�k;�^��Gg�Pj#�!4���4v��ܧZXF\X��c����K&ְ��fnR�i���j��&�� ��'.�=�.n���R�dd�Ղ��\���=e�U�F�M� ���a����{��ϫ����\�JJ�Y���a�pt	;Ż����`6�'l����x�dNw#�E��_��/#h�����@�1��Ѯ�\�Y(�'���=w��<: ��^G�.fDh2���bX1p�
���]�C%����BK��;$�7C;�*?���?����c�enw�~��
W�vZB���~��c�O�������qo�qNCxJ@�WM��ݾ'�!���6���O-Q�5�׃���Z�OS�ʐЖ�Ze
X��4+�c���X̶X�-R�����Mdv��p��z��F���}�[��ȵ}f�ZK�u��� ���dR�s������U���H w����~�Â�y����"�h{YF�1������7�"�++H_DV �I��Va;U'~[$Ԅ�&�����j��+���:x��y5VM}߈iF�Pq{��sVOC5��ѣ���p�8��
���J��m�mh�-�;���aLG�E��S�bK�tP�:.���:{o�S|�#��1�7"�L$�`ڞ�W��\�K�(��\�-�>��~ﬠ����ssZx�3Q�o�w,�x>�f&�!�)��?~��,'��7�������������w��q�0Q��ֶ�H�yosK?	
�|Vv����䲰aw���h<~��R���lۃC���~��"��oN��$Nt\(3� t�>�9E�0�G�7fjU���b��
������.J��h�L�ק�I���|h�#�o٠g�j�p�&8�1t��q�g߃X�;~׸��BH�L][��� �\[ V���>���`��+'�)"��0\ħ[0��R ��DK��M�yT������� � 
��N�☂	[&�&)n�7�GNG�3��P���
��m�*��t ��o���/�'����^�[}Qܗ9�����u��{�7F��� ����p�M�-a�j�p�Djip��7"Ί����FK�~|�8#QdAE,oW�Cn6S�=�5�/�l��R(-�+Uz��G�k2	��*����:�啂.'{���b.54u��47=��!T�"��^�+����_�זǘ"��p琂ѥx?�w���
,8/kf�K��G��%��P�١�l�qA�7��rPF�A���x�H���G�p�z�)A���~aKkCa�@��0M'6�'BGuǙn�Iv2K�����DG@�\g�E+���R�H�"8l瀘�Ж��UD�#vL�!�n�0��/v�Sb���np�oVga;\�.��Y���%��ܧ�v�c��	�u��l������!~�U��t��j�f�����3��^B�*�{�5���e�V �n�;�WN;&�"ߨ3�����Р�O�:���I�8L�n,�Ñ� ��q>�#iBrn3uD����(����ɬ�c�7��:�~b<���������4'�G@�s�Z϶����>QǺ�<Df��n��)J�)N
��f�����N�qb��$�ЩM	#S�$�]s���Ԥ]i�z���!1���n�{�ٓ/(����)�	J(@�Q4�(�(��Gx�I1��Bm����}�A�|{��z����lq�BQ}ǝ�h�1=D�5��^�-�zY^Jٯi[�ز��`v��M�Z݇������3U��Ԍ.�Ve;%�^Q�����iRD�����G��� BB��0!�upu1N?zS���u�L�G�(�쐒����A" ��8"��b��|��FY�1�(���!U��������4� ��.4�QUi+����C_
���8p�h8��B� ��bz���@�׻܁S���x��a���w���\�$|qR�U���qX}i�D���	�T�ڵP��� ��|��8?0m�?�P:!��8�;����N����㱮Tda��VM7GyjK�9�
��O?K���-��	{�s/����o��S+J2������������.�z<r((��@�vT�0Vlt���R����'b����:+�f\ڷ޻D�U��Y*�[��o�*?�9����Bn���:k��1􆘩S��{<'D4����驟�I�9���
��y��x�ضiSI72m�S���4y�@����q���*�M"�Y����\���&� 5��Q$��Ԭ� �ƭ�uέ7��U�&�20}�0����`��iIB;Y��ßjx�L1���\}ۍ�Ʋ���@�Io�L��)|�Z�8����a��_�6�8��FN&e�'���˹Y�q ��.���^
q�d�)�~y9KaR����z���%��w�w݃}�8�u������ߌ̎SJ��
���g�ɀP�1�TT����B�sq�%�����^E�'ZU�'B��~)��^vw��-0���p\�ϕjapxb_�S��u��m��Ԭ<���A�N���bz=�SE��M��:��ڒ��[�[Y��f=x�}���f!
��z,���'��
��%����[����`q�Z�A-�g�Pi�� :e�3K��Vq�K�c���E3��جP���S<�B(2�A*�~ʄ����䜢���Ը^G�����(eF�90�U�A�1�זz�]���Rzp#؄'��N����NԷl#�r�v��"n)��!��l�ƈ�#�&!���´�	�S���r#!1�u��˽��;�mb�ڨ��p�1SɊ܋�q�%[�#�W�󙗿o�2#��N���X@lHY���Q��i#I�0��?C����ף����SHj��3�׍IΞ��ü_�(�g^�I����9��C�?��A�$\N��4�;S���v�C�]�kNA�8Xs�1�q���t`_߽c��՛K��D�WN�a�2��t�]����'|u\৩o
,�jCí�О�+6񳾰]���{�3�s��U��B���pBX�@Ǜ�x�@4�pޛ "5�˛n$��8��L�ټ[�b8f��IWɦi-71����O�^��[�P�NW+�d�r�5pе���&�Af|Ãnl�BW��.�*�]L27GJǬ��`�����aC��c)�v;M�ʞ�v�R��~�&�?�U���<������M��ʾ~{��礓��3$���C���b�w�z�A�����ͱ�Q�;j�:k)�ï���%/�j�rd7�P	S�Yo�� )M�	b/"x2���M��5U��W�u�8���VwS�s,Ӗ�C��L��ߥ�8�{`���"#&L��z5�
�\*�uȐ�-0�?Ǚ��<,+|r� �i,�1��R�Q�gYLd�m�g�M�Ij�nSk=P����`��擝����|$�[覱K�4����7��pK��<�	�1�%�}$(���͔$Y��n�mg��%�	��f���)t\;$C������J�ۈX:Y��X�2�7��� �j��_�zl��1o:�!��Y��{���i�����/0o��ŕ�]��ii�}@��.	Y<�D*v�m3�҂�}dV癈��^N�_���+�}OX]��a�� F�	��ϏyZ�݋�^$�ȷ_��TBE�~��V��cw��w!Ŧ8zQK
�|~��i��?s���/����� Of3��4�<���͏*��ϱ�I������������4�����|�� 7�,�z7��c8~��'U�M���?��J9����Ԡ�*$r�_�<'2��Q;�����z�m��c����T�S��ai'w�D���i�dR��pxM8.w����� �V��Kf����/�ҝ���#�U����MqW*,��R�J�!ρ&3\�&�a�Ag]�L��"�?!ܽ!�3!ө�%Q:�#�v��n��M�߁[���'0��J�+�>t*�4y�`������#�Y�[�K���Ā����7�t�e������!�&ޛq6��Õ�Ĉ=����S/�:d'u�1�jQ>�
��mM�¶MJ�1�7\��r�/ �؟�	�Y�Η����:K���������g8w)���Rc�0�x���Ü	њ�o:��c;z]�� [\+�h�{uI��{�I�-h׌EV��!s������`��6�mr��:__��ĝL�v���������G\R֘.�e�J�;Y8x�$a��@�Ԝ/%4�����J>0 �3��	z��ݶ����Z�gk
�m��*��WL�ʋ��w��F��d��0��H�����9��� �����.<Q,j��PgF����|��hOH3A�m�B�m\.����q���G*u��P�b���2<��F;��	x��/v����q��ϭ-��s�E��Z_`ak�y�ԑfٱ�t��\�+q*�m�yq�ۅ�ΰo$)�Z_g���0�=�P�O��=�)���k�x�=ww���d&�C2��3�H%�j8Q�0%]�����4����T�����qZ�4;�Tz#z������ڋ��R�+V%٠l�/7�G���	���?����h����B�wG��_����?��|�ڂ�����}c?�5V���/�3/Vy������Y59�g�ns�>0Ta��k�O�H��!~��=�wu��I[�Y��u�=��s��:�I�t�Z����BE0��ě��	�Ű��+�c)�?9g�L' �x�(��,�+:��$��^� %��o:\���f/6M�8��h~��Դ��ւ�&x&���JmEO��{l,�4{y�6e��c�tF)��cƴM,�R�@�rU�zP���U�5��Q߲���Pw2��{���iV�-Fv�$���P����Ł0|h���u�o��r�Q�M&f��&a��d�����8	��w�@h�.��9El��Mѐ��3�(�9�t���߂y��W�2@��� zLSF��-�?[4c�Q@>�Q���}�Y�HQ�HS^���8��2Ը�7W'��ӿǀ�v�r�Ne���M�i�e(������4Ɉ�S�i�� L0�%���W 6�ˆZ%�Vާ�3~E�y>F���^8"�P���(��r�%<� Q��]j�x1idʩj������%R����'�����X=�qhZڐ �F�["Q�����i�|�/V��":sB��콄jX򴨘ǁ<*�K狴u�A/hȝW;@yD�R3h��WP�'�^_��2s�W@8X1�x�䊝vV�H~8���S�p��2�>�ъ��������i!��!,�%6�D�)}�9�ץV@��Է�I�4�K�&$����le̖�5đ�G�����r�a��~�n�$���ƫƠhb�/��5j�y7w)(ú�izň��^�kqU�Y��6���26y�?��֬������{��-�"-���/:��T�*`�;U~_	
/�	T⥀�V��`Ik��{���~����h{JJ`�q��7���֡���uj׹;h����_�)�$�{*��נu�mא�_���PQ�:��ZZ:���+���_p=�1��ܗ^��u<i��0nfx�N2�&��B�1P3�:V�q�#�r�GF���רȯ
Ł[T�� :eB&aӵ�����A��S�с�/��K�>o�u�$}�Y>^o�0��n����DM?�1ZFOI��x1�.ĸ���J*��m�S�����/z �z���3f���T���B��*��C^H�/���+
��'�D:�ލRV-��D�����ub�G�5����e%����ȶ�'r���U^�
-�H���^���a^+|?1��ğj,�.�smL%�M��V��	k�j�z��/Y��'a0j�J�2��ճ��t��>/)������z]T���K�E����s���?Mvr@�TԎ�w2�&��&�D��J�61�H�?��7��݂9խ��^?)��\R����v}����J�n�|�K=�Q�EOPY�1����h�jzG��2�h�F��x�j���*�J��x8�۰\]f^o<M�D�'h�=s4� ����Y��=����|H9�K,[�|`��P����מ�h^�hvߞ?P���.��E�vQZ����[`��]}u;���t�$�>��	��{aL��57��aXᮩa��a��?`Hh����\�����f��gT��<��0L�f���i�U\�
/�Y%�m��.�H�ߕ���O٧�9�~.��]1#�v����'��
���)����	�@��\Og6�Q0��bB�G"a�9rE�&�?��lzMڱ�#<����z�r���Q�>0,���@ӠoK�s��
�᥈��8�P��ED��}�~���H�7$6}8���d�F���
�B�����yC��~�Yڎ!��9_�Fr"�UL�0T�
 ��k?#�h��?Alc��*2')�������é�N�yC���
���6ZġJ�Q�vx ��!��j.a�=��Β@r��V4Tr�%��@
�dv���-+��CS@;&�n�@��~Az�Y2�6�aqd�P&��̴�}K�q�����t��!̭v�3��*���B�|ziPR��Drf x��v
�	��v�N)5�X�\�����C6�U52Yq
x��	3)��ڴv����_����>&	�$e�ٕ�#ܥU#$��nی{x[������ũ�	��_K�����'|�aG�t�Ӝ~�X�6R���9�%�QyC�cjH6��|T�#��2�tl��f[�C�C��W2,����EK�ld�P�]��.n�Z]g*ʏ(�S��.{�l_^)��̠>�Vj�M7�Woߐ�9���b�d��Ju9�g��歬���6{t�Ee�Uf�Ul�~#t`rZt��H���o�9�Q,L��x�fjĤ�Xđ�h2z���q�-ݕKZ�W熓,�XO' 
��>��Gg/�K��iN?y96���<m#�ءq�?�D$dE�"Yr���P�����
��'��<:��pHb��~$^%����C�h�)�����Z�D�i�E���-��RX&�I}ɘ�π���ֆb�<�p*�tn4�(�54����e��M�b����zE��Ȍ@��ݲ�v��?4�%(�Ł9}~��0+���0�8 ��>ߎ��Z��gF��y�s@�D�]����5!�Ě%��Y;hLSz�� g��Vcm��E�t���?�����p��2� 8S7:Sٕ�ހ�	h�os	�ՅOJ���l�� �p�=�l�˜ ��Ti�U�0Mz)��#-F0�GM!x�NԔ�ۃ��J�F�Il���'�L=�5:pUpWה�-�p�adVĝ􇋍V��l���΅��7�m�+�@[�J�9��c�>@\��5ѿ}7m�S�1>?^$����27Xq�/\�R���"��@{��i��	WU���"���c�5�����(�q��PY��_�L����܇�梖ʚ|g�?�K��¾s-Q"���
�3h�*��6������ ֋�\JkS���m�8F��h�pW0!�H����I�T���E�y��Q����:�k�S&t�Ԉڸ"�v�2ɘ)-�B�J�*�����5�VT�.g�֬f����U�����{,��^�0sk�����	�ع��R�A�����5�W�$Ĉ�B�}���p�f��D����}����L���#>��ǻ��ڬ_��`D/�6^"�x'~����@'��c�ћ��	�:r?v�@,��y?��X0=?�^�
Cn qܝ:@��[]�/�墼z� �%*�@�鎦 ���P���b@'l�⽜�c�/ns�b�p�r�e'8�@	ڶ8N�Hb� '-���\<=�g�> �O�,\�ӕ���]�~���Y}�c��˛��	$�4yHs���L����2u�*��r����oY$��u��`��B�r���Io<!��c0����T�o�='��5]�V]�7$�~��t3�z���v�35:��d�����TI�Tb*��߻����[��l\�>�$ȜRp��x8�#��}��%w��0����JJ�y�^��?x���;ٙ�`i`f��eekbB��M��" E�o7�8�=�%0K���3m�*j@�*��
�t^s�Kt�St~��;W���=]g+��E�7Li��T*��9���\��rAyf62�H��>	O�ŷ��o���:Ӡ�"��U�h�K��k�!cK���@��'��|q���icr7r��58fON�%�t>W�Fѝ^^�]Ld��y2{��&��{�CJ���H��ù�;l�����[�R-I+�Q2�q�?��.�����Q� P����f����Q�o��ei���aj��D�S�����.W�p=[�VΡ��>��j
(�Y��&Ե����V���ڔ�!��QRK���#_��:����¨m��{���I;v&�oa/k$���v��m�{d�?��2���襵c��do�O��<���`�Va�����ч�'j�P\�1qL���p�_r��޿�mo�)��X�<@�5�[mXj�ϵ�I�!_[#�s&4%��9Z��N#�Eܹ���p���e�(o����^H>Z��j�{U1�����f�!��MC�yO�^ CDI���Ǐ��ȉBi���mZ�WY�(+#�e
�Ӈ5��ֹե ���>k�2�e9�����*+���*%�U��?�yD��]�Ɍ7qP!\=OP���������6T�oCZ�/y����Ls��������'C�����H���臑/���HY�E�ߩ� \Ln�@�i�AGh$��AHٱ��kM�4aP]Ϧ�=�9ה����jw�,i6����tMRj7���?�)w>YV�;#b��A��r�Δ�!�)��sG(��"Ҿ�I��oy��[��I,]xNoG֥�s�4!iP~���;�f9��'�ڦ^n2F�%�뵺aAkia����
�� �A���q�q~r�����?�Zh�	b�F�Ϟo�t=G���V�N76ꞅE4��?�xӄ�x4�ܬ��Z`a�"�w�n�@�ơo%`dƱ�.~�׮��%/`�PTx|@]������Iс��e�,%#���8�1���-h��x�Cy]S?��5)���6q8P��@������`t¹�/��΁�]�
H
�j�N�%�T��iȵ �^�G�����S��.��!�8�7j���Iu�x�1��/�<��(���gxsw�؎5���h� �Z&Ń3m>?)S��"�
l�ƅ�X"詑�ȭa�CK��w��u& �<tO�^��qw�t�&��O�o�J��4.΀u&���K�7X~�"��}�,X�9��&���y�Ȥq����T
b��R�)��\�Z���%�V�E�U3nt矱.�� �%�m(� [�c��Wl�����E'��ٙ���Z��,�L#``r��ǣx�ü]|�r�3v:��]��_Y�y�0L��f���O3��昚ޠT1,Z��)�8<�y�r�Mw��9�?r��[EY�>�qN3�[��z3��q6M,6�%/5����k�S�lp���mk.Nj��aT�1��HyxE�H��N���I��ʷ2��d��;���w����z�Ś!*O>S�nfk�Ё�"v,Sg�ea�\�G{��)ǝ3t�����v��/X��s�(@�BG��q��B�z�2�s�Ӫ6���IXQ�S�NE�_,�^$�!�*-NJ��0�xn��_�d2X��A���ʄ����ڤe��2jyh)�E�L\:�w�� ��!�۱�(h	�C7/��4�����ObM���o��˞A�.��V%��9�d"���:
�Y������	���ApJ�-��I�G����Q��t�+�ߤ�OqQ�r82��';�bA���9�G9A& �@?��r �b��'y
[{���C:$H�0�]�aq��s�|a]h,P�E��\Bֽ���&5[Cm[��K���b���8�R�
�/��K���[>�p@����H������<d�K帖��+xn�߁�K�t��{�'{/H�����&¦(��>�j����"Rc���c�4�yů�!Bn\0�)Xw6ƅO��?U�2���*��5��J�
$A�W}{sa���h��E���_Ҩ�ф����H�l�q�&F��৕��9�=&�c� �G�� �Ͽ��J,$ƾ��N2@	���Ok ���ò�e���sՋ�x
�^@ZY�Ѯv<ǩM��,:�2��Y�L�]��c{�w�@Z2��xR����m�ޣ�K��ݐ�F������IB�]�qN�`��o�^5R�����x}�@�{Jd��D��&ڃ��n��M��?|5�U9�a��A����yT�x	��b=s��
�}*Oi#
k5��_�8\4�!6Ǳ{\���At~m�T�����3��!��G���M;���]��'�ÒЩ`��>��:�N�\L����C�{������$m��`J�R�[�c ��c!#b*�%"�lט|%6���}t��O�f��B�Dv_^68޾�]��[e��B0�֪T�h�Ů{B��i�Ta`^N�刎��z}~_�����r�W�h������τ��Iٙ7�Ɗb��c"xL��ϡ����:n���+��FJ����#�N����2.G��3��>h�F�����^wCD�Ɲ���+�E%�:C���I�ͳg���e�C�1N
���	���x��Y�f�9
ν���2X����KV�	�/c�\Xb��Ղ5��Sf���"��U��:RL!��Qfx�)F�1�Ռ���u �Ъ��9�?!�J��M�(�Ig�o��xl�x������N�m�M2_�Ht��韣\��`|�`%��,΄�gr��e &|���ܺ]�\�I9�BT�`!)��B�u8�UJ}�Fn���a�ӱSgAG��'�ީߕyV�W�&T����׍�������-53I6��M+_���#�*�>)G�s���Q޺���䨂L`�Mw��ua~L�M8����E�\�����[�Yo�	��g�ׯԺ�!!��I(L��`%>y��\�z�l�a�ޑ�da��`�L��X�����9p�90\�ZZ���6��(����Thka$�+����l�2盢G͂D�O37C/�poE�f,� �G}G��i �Fv�G�u����c���w�M�
=�Tt4r�q��j��e}z�����7�I'�1���ϧ��F�"n��E��vh���j���`����b7���k��h���ĉ��|#{m{�7�s���E���m�oPF��}C�=9�&-r��2(�wO�ӓw,�[�7.'����B�_m3�}�h5�����#�5R�g��+�� G�+CL���=�8&�x�Q)�)A�y�ʫ9����b�)�>�kŪ?0%ԥ̝�"�W3�q�O���.f���=.E�H���Z`�{N�J��+�2�T�QA��<i�G`���y�p����a�~@y�FS�ꔼ\9-�4���1��f���~)3�϶?������U�M�T���\cG+�>iW3>G�8�����E
�,�FL�GJ� �'�2�VY	cҏxz�U�i�y�U��2�B�䆅�Ye��h''^�����!�p�3��C���vR�:�rB�~�/U��MC�� P��%�Z;�b�[4��FJR���B��b�pN >�u�UDi�z�r��4+�S&��z�į���lvF�`@Q�=�R����3����g�A��-�����ԫ	�w���+�ׄ梂���hY���Ff\^'�����NG�+��53$#P���@i��v{B�8]��Xy�vl�K^�h=� �E�k%uҙ{<����R����$�v�5�"���/�O�!�𽾾�I�*~�k��1'�����Q3.�RVpp�v�t�C�#\O}���1DF�7#oˊ���V>�-	�����>�NN ˠ5n�S$R@�ھ�.}�ؑ�1緯7T��F�yn�A�������%B��úN6R��@ݾ�%an��R�l��� ���`�$��o���*qQ�^X�a��}���OǨC͇������v�R�������_s����Y�������Y�z�,4�wyH�e�Fӎ������ޘr- A;��=�TU��I�%;h�(���#�Q�|�d˧��ŕ�O'�_�!%k����9��0{^gaK�y�"�3
���K7���.��c�Ǝ����5�����I�'32K�F�e�ߊ���!K����	�J7��޲�m�c�K�4:A��UB1,�.���&��s�c�o�+���}��D��O��M�-
b�9�u���F<0��V�Xڭ�Ë���Ѥ��L�]�Q�7��x� ��j0)B��V'���k�(D�?��DP&� �G7�KH؎�����_'�':BlL����r��u��i�g�E��;��z�2$���e�r��L���g<� o5�}Dƥ���Z<3�I��&(�G��%2�R=E&��atuD��n�D�y� P�2�����dKY��_D�⇪� ms�邲+1�G��̣lJ�T���3�|Mu�ni�[U����j����o� a���˗=�i������k��CԊ��\nJ)+6�T�b���Fg�U�L���3��)Z+���U13�r��ZE��8zt�@�?	���B����	3\g��zU�d)�ٿ�Nfd����=���P8o�F.���_9v+�tL�˙���6�Ӫ|#)U��~bRI�K�_�"*Z���A��[fxH�B��^��<*GM#�B%c9);�wN�΃�D*��R��e�O�.��4�@��
ʐ������H�@ ]%c[ӻ+�e�q��V�\#��^��������3���q�Ϛz>���R���0n���R�-�O�k��X�_4�{�\��l���y3�� ����i�l�:�rz��y�:?��U:���fm�fJ�<Ґ��̥�)~=�Q�r�R,~t^P(��<�QDπ�����S�V~g��^17%�b0[1���S�5��F�����:�5��;f����.���y�Ɩ����?���/ ��t5OkQ�ø�$�{�D��}G�"�V[�<ȥkH���o�T��Fa@���Og�����J·Y���_l)J��9te�:�A}~ږ�-£������<�	�S!S�6����LC�k�"6�����!��g@�/��|x�:@Tb���1��8���S�ng�L�W.rN�Y�>��e��rhr�fܭ�9�i��BrRq{��K���Ier�%53/���+�6�F���+�CX'�8����_=��W�*��L���W0�Ҡ{�
�����0d�S����[�������(ƶG2���ny��~Rz�@��ﻼUXsj�%t���xk��@+�C?�2�N�ύTGEI�<�\�B�	��d��6ݜi���!?�6]X�^Ԙc�}n#{/����7N1U7~6�Ebi�k�@1G��Ʌ��CL�P��4�V�������2�6�D���O-��U8((�Ō7.Q�{����)Qz��ט�J)*=]���Tޥ�?�Q��"rnH�Fi�R_�zR�"�,�)c����'��o�v��dV�ْf8[H`�����"H��bG�����ܡ�ֽ��]̸{���?l7��iM�( �R�Qҵ��~A��7�
e���Ֆ��Yԛڃ�-m��,���S)�ߢ���lÒ�8�_;`����OqZx��f2��L
�l�ϴz�"��ɦ;@%�1ifAQX^���"C- �c��H:��� ~D�~�� b�A���4�ˇ/-��M���Zz���% ��ѻ
(�ڹ����a�p�1aa�c�XU�-��b�?M���	Wzj!)�32ƿl���P~�����K\�+7�[d��%�ըg��*3�d������/A��ZD�L(,.�L�� �����k�GmR�'�l�A`�iĊٺX��_��a<�����Z�>�ԥ��8v�<�3Еã�H��=g�;���.f��]-`��-��%����.��Y@�g��$|kO7_V�E���Ü�(�k����3)m����ʆ��fs�U��Ğ�����4L�<����_!o��9��"=����ȇ�rw�H�9xpt:O����ȇ���Űy��db���9�R��Vޅ�ڴ�q��Cފd���>,�|Ϙ�Q�i�q?o�v�����$�`6ڒ��P������RYK�q���;�&�+�5U����8к�t��mt?$P��=��>bw�fZ�(�:؍t�?e�T�	^6�^���� �kMʯic���!��r�yv:�1�{KJ��z������لf~�K¦$�6��_��F)���J~6E���p���>��� �J5d��/�>�]��i$:�Ҝw��4���s�si��0c����68J[���[�����>=�w��Κ-�H�vJT�]C��ė��S�6z���4��X:�!o.�ݧ׽Iy�m�2�Ui!Q����A×�����Mi\acS�P������/qmLž�ԟ���@	$̋ճ<)��@3K��.$��#�\ҋ�)���3�>��e�qc�Ϩ_�|�Nn]�дG4-��%����C�b׷Cb�UP��Vم*2q[��1v��1~M�=b�˞����8�zc�_+�H��IF lu]wH�a��FC�u���g���"�W%DH�Ȅ�͖���f�3-�N�����7$��B�d�s�mf�N���R���8�B/J	�����x�%��S{�@K����_���s��0L��mdHR�&碕�IVط���k�j��/u�&r��+b�EAl"�g�0�IM��qM�5�]L�l���|ԓy�_ʕ?0��~��e���̾<�G����N?iT�m3N���J1�#�|���+�����⦪��ʖA'�o%�Ob�m�X镺w��I��%���X�i�v=l9]~Vf9�S��b�xu�/f�HQ�*p1aP��f#O6��-g!~3�=x�+�9���3~�0}��di�N��[���\p��G[-�&�x�Ma�<���c1w�GX?>�v%xDwcJt�ckk6}�9����C�����P�ǃd�p�Eq�-�"֘)�WM������*D�M�.�^ff���|�b�(Z1Ӻ���+_ �Q9�\���i�G�����‪nȓ�瀘O��yYe���A�0�ɖ�i會n����]:���������O3L�!�/ �'Z�6���o�T�e��)����kb����L�u�Ɛ ��)�!�|�?1�H�/Q)���-V!yx�ZI��Ҵ�#�� �4���6��`Ru� �u�2�$qʷV{+ղ���/�"K��Bd�X�7B�uW'�=g%����Cᧁ������/���n>/��d��pt�KB��ě�����ꮗ �X�,3���Mi��7�I�=]�V���e*�7�X����,?�6�a(X;���7fN6j� 5#A��%�������O<̰�nMф�T��\���|$N��Яb��|�q�B;4reBg6q�{=�4z궫�'$��H�"R������(�F��ZJ/��4_��+�cP#s�Z,���3�;.�Q�W���N�+v���H���|��: 4P�Ylx���c��W��u�v�I��(��ʼ3���Ջm���8��Q3+�ې"*�A��*��b�H�3aYN�3 |B;��ԈO�~�	��Õ�:������vXV���ml�=�¦���ʌ������a볣���AXx/��C��T���4�S�-����+͛�f���Gu��f�yÞ��:ݨް3У��w<Osj����$U�^�4�!����E��l�U���p��?��_�N'��Ț����A��ז�ʷR|~��W���Rd/��������x��4����:���ܤ"����g�$�M�Mw݋����-�z������)�����e�twrb!�&����}���,9n������x��,��r$����M(�M:�~�	��,��I�������w�c'�ws�-�� ����ů
�ƹ�W�ą��/o�7�]F�I3�hO�Ʋ����9ϯbBʻK���=v�U���\i�gN�^��Ņ)|�lY3�B]�_^��k��<�K�%�o^N^�� Q�e�o>w}_���E�&�VK?S>�V+ES�O\���������h:�����гw�������|����m<���}~�࿬��<�v��{O��F����'`>��Dz��� x��D�GPy�5�U�=}�y�̙� ��+;�f��p1P�\�1ؒ$����S�P���Oj�[�j��ڹ:�Tn2�+�`({uр}��7q���'�;�5N�Q{*��w���R��i���P�(4z����">�6����ߚXB��v]�0l1��w>8 ��e���h��/�H=q[�<��'�!J�^��0��h��������+֙�?&��b�����*��k��Z�O�U�G�V���$%ވЛ@kW�^'��t��y�`�U'@6;"��l����<3*�Pz�ܮGR�{�A�Aud6�겈+6t,CP�������_�9��;o���p~����;�u��V�^�Zʤ�r"�0�ӽ/h�4�σ��ƓE�G���0�c�+��𑘀���0}�m0���55�'P;RWrkJ��3���g'*,���_�)��.�1�'����vF+�&��)}:�]�S�������~uE�x����a+E���X���|�E���N�5�-�cV��mWMle��2��Dg�Bc�Y��\��}H��Gϰ�H�Yo�O1%t�k:y0���#���x�#y��!Щ��.���P�����p4O���;����E��_1�g2T�3�77U�g��7.�7�����"�s�>�59n��zv��Z�a*�,n�j��!����	�D��i��M�	�GWյۈRd���j��c �e��(������|إ��5E�A]S�E�BC�1�{�>��w���i"�͘&+B��j�(�0+~�zF���KE�y	�t(���@^-�"k�bh�e���V�L��C>�8��8.�o�x�Z����)�������ڭ�Ng���;A�P�K�i�)��ZA�׀�;�zf�U�����K+6�l)�,�JKg��6���@/�tmuhS/-o����ݓ#t��Ѡx�?[����X��Jb}�|:"�Wd�x�;@f��ɬ�zE빍�K���9LL뱟�Cǥ#HŬ��T��BBR}������&(g�o�6�v�Ґ�ʶ��[cR�;o-��W�-v_��\cp�4���fb��A��׍��#*T��iiwK��3�G�(Óe"�h����Y���XE�.������YF�z|���h��dp���r��?����[2zU}Sr\����
�Md?S�q�B��	�XZp��1�}�|��/�/�Шd~j��j����"���9o^�� ;�_�jKYP(G �������iX4A
��\�	��M�~E�3=����puk�s�%__D%��u}2=��g�0Bl(�=٪����� M/�z��V��[C�Eq� !�d�x����+�F�f���=(��ҍ�G�� �� �I7i�������uw6d�8.����>8�;��_�:��2�@�i�}�E�R�bg_����3q��p��m.M6<�Mv%R�������U&��&�(�����Hyj�8j�.80c�kh,��|���k�o�����e�_�ZK�K�:��/����&ۅ'�\@i���L>��4����!lN
�N>����u�o��˳Y�L�,3n�<k�+-u-�Lu��;TF��@N���l���.Ô_h�H������*|}�!����HF3S���[ك�=�M�K �=;�ڀڭ(�`��$���Ϸ8��ЪU��SR �]h���.�2.3�z	w�J�@�N�;����)���-�n���n��d�O,C�p������Ǹ͌���F�š���f�ˏ'��7^�f�ފ� �p*%!����߮^����j�O��&�����ě�f���u���gҫ�������#}�/u�`a�ʥ"2�]Za���%��U�r���hTxԱ
[̠EP��������7Kͪ�����aھq��S�|���\rkW@[5:_�n��&p`�:�3��t���I���P��{߮d��f�7jC1����>� {+��l:w��-�dg�bL����Z�kI���Oӆ�[��=�0,�����}��
5�9�%��I��"�lg"��uzу��o!�8,��xy�@�ӌN�#n$[��*(��K@��y	��d791U1B�"�Xh��`t���k�@�u��*`�=:�0���5�N�*e��3V��܁π*�J���[Z6�2�
��x�~ۦ�����}.f!o�h����I�L��R�*������� �K&��I��~��AV]��}��B4LK��U�� zS�c=�d���%�1%[8lk��^�T��� ʜ����3���o�!y�:^���L�_1Y���X����B�DԆ\��[�kߝ�~�#3������%V�=r/h����������ř��;$�om{l� ���Os�#��K��pl��#�S�G�E�޵��{���`s�f;"%��>t��SR��z}�f�P6jL)��%N�����w5hOs )��QZC��bIN}$p�ô�:�"=%�/�h�_�"����\C�T��l�$���8�ۀ�1���,��!�t ����f�л�UVr��t����A�5PS�6��>m���I+G���F��������W�X����^C��ھ�̓=�����L��%���� 
~�D���]w�+�A�B�X�o�Y��jᭁ)0܂�PS�ؘ��ўM��Pcb!Ь׷[֣��t|��aM��bٸ�C��� ~Ϣ��y�s<���
�U�u'2Z�{����?F�M�5ن�t����� +��]������T�j�����(���ņ%�����}c7��O2�3�l8��a+ӖsP ���0���́z��2�$֤����³ 8�u�(l���:��{C�� i����Phl�Y|g;���ބ�C��(���i\�	��d�����z�,���1@��Q%��&�����0BUL�G��́|�QB�����:���sM��{CRv���	?T��_m��v��in����f�n���J��Å�:k�df�Q����m�%b�>��G��G�,�0�!��[��a{�ȟ%��nP�M��\���Nz2���;�n:K4�E��wT\�E+iC�b/�b������S���x���F[�t"à��C{��.�B��m_��{��B�VSu�"ieiܐۡ����b��ˤ�m{���݌��b~� щ�4k�)O]K���-�lAY��M|n�[����e����Mxn!ɐ	�ps��������5e�~�Α�V��!_*��e�+"f;R����pd�I�� v���_p�ʹgP,LqZ���n|�%4���$�j5쿒���S��V��{jEr�KIg��@j�Pd���4��D����u��������X�����\l�ZPr�\�zR���d-k�1a��������� >huJ���U�o�:b��X5��:'":�`�EK� �߸�e4S(�q"#t1&c����'T�s@En<Fm��g�F��{2j?�V�j�x�!�E~���Lם� ��4����c�rj� =�O���:��eIqU �*��HGZ#�X�Cw��'��=fM-3S�3�����mj���#Xy������� ����A���A3s�jE��h��$�
v,����>ڝe�r^|:�v헩(B�(��I�̨9E���e�=T�w�1����>�ͻ�Y	�J�7��,�6����u&q���`!�-�Ы_���|���S��+1C�+��,N��2�QP�i���ك�aª��(I�����?�r������z�2�Ÿ�w����qW�ط���%���C�֒R���f����&�OI�{���dn��5�\Cܝ���kk9�h��%q�pj��hC���u�B-=a�YG$f/᭿Z(�9���7��}$��=�<L�<2t?���������Ogy��@��T��=��vL
z[� �(dq+�IZS��)ИR*}T�ɠd�͛X�o�vE9���Ve, {n	J~��3�KQ}+��0[�jZ�����ޙ�wTH�3�;_���_�Z�Ƌ{i�!�����Vm�z?'���h�~��d����E8�d��t�/�Q���Q4�%��>Й��v��.�#�"(^�=	�����
����|fM�E�z\����sU�+�qRȚ�iYH#��v���Xm�ã �As��l7/��6l[E��Z�\���=q��٠s�����4�߶���kT���P�fC�2MT�-��N�mgw�Ҥ�B.4y���7<,N��MO��
���W�4�����uG>����AH���Ml�O�0��VЈE+�G�2�~����S<X�۾�ym��#R��M7iC��(�̐�;-�ފL�(��Wm��>c�E}�B��^S&7������Q=��`DO�)��4,�Q�c�rE���q��bV��/�v8��V�~.u�7j@hK�)�W���:��79Ĭ��@����k�9'[yF����!���W�iU��q��<^��Cx>��F��#����l����K��pR�9��d� �=�񰷹��L���eܣ	h��<U)����V�z-��>�3ۚ��̧K����8,�6b�ſ�Z&��u!��	���`���//���8>���nO���/D)i���;��y0`g_�	���ȶ�s`�fH��z$�	.�d�O��Dc��l%�h����)�C%�w���Q�`��jE|�u�y�}X}c�@�
�����8���B��M◿�1go΃��s86J: �E�=y�ZEk��P�׻n��u&�Y��8)�ܰ�d��*"�,�<o�>	�(�M�d�${w��n��WB7������S�kóxW?�(���G�V1���G(�:��#|Ӫ��d*_;��!�d���m�қ,�,
�'�Q%�b7hc�K�X�wM[C��a��R4Ѿc�N9TrVW��*"��֗���r�1���F���<�k���%!\�Y�"�1�6�<���@�Ԣv��H[��l����c�����lИNY�$�Ǟi*�2�x�Y�z ������c�J�dr�6�އ���S����O��g��]��	�g	d l�q�e��>�W��.|L2U<>|B���nr���_�qu�C�Uȍ��k�"��^L�S�wو�m������yv�w��X2�O�,
h�P]���Oj�H����#*vs�w� .[���/��qA�j7��{���Մ�q��0�����Eӝ�d��c�!�OJ�L��e���U�7�׽� ���{=�=����ް���_ed��P���r�����O1.dQ]�G�;�{Q��
1,Y�Vps�E������6�	�t&S�ρl�x(4�����ڰu��eC�1���~��3�����N���7�Z������LG2�Q�D��2:KL���Q����E�TWȡ�Y���ьl�㙅3%�FwD�g��$�I$�rW�*ĥ��#vz���|���'�{����(a7��Slǈ��-��*���'�]�+ }O���/l܂��s��#bN��kbϳz���N<�<�~�iA6E�:�F�>?9�~_�M�0J����T�b�C��N���V�j:ko���T��U��1J��4�%RO�M¹�X���M��*��Hl���I!J��Q<36��2�\ںD�ӕl99�!��q Ltq��HU��YO���[��b��X�ܨ�x��+~g�Vhʑ�W��
H6����ƿRq�̟�c+w���[�;�o��dm���k�xt�~N�.x�EVC�9�F�D���-�H�=�m(ȌDf�ا� ?�D��EDE�a��,S�7�'�Ih-����5�����Zl["}\��-��.�5�L�8���۔x�E&B._������owʼ�����	��:6�A
`'��F� ��:Ha��1��9��l��Z3]�0Zs+� ����������S]�7����:�~{�M췬��=qŸph�δ#���:<�"F�d�D��x�x��q�������\7� 87�:�}����W?S��ܳ�����m�i�
������ፓ��^C���Ͽ�!��Q93-%{�RZ^�%�z���#���}T���L�y� �Vq�u�d`�|9���8x�~ox�p&�˩u��SНeR��B�G*�'��f�ҕt���:��'�;P9L��or��x-Tm�
�)P�[ջ�E�U�0<P�;��*���c�����#�:�eW�"=�铸�SO鑥ŇS������q�H>�A��R� 4���N��\n��K��c%I-4z�?�M_&��f'�b�Z�>C�bشGu�ki��h�U��KT"����;[^��ɏZ�5j�?�Ҋ��5����RoD����m�[Z�o�be`��8�Dz����k&'�e�H6�\�@�G�L��{�Ye���R��։�f88eo�b�K�5f}��I��j]�>b�؛B6P�)�=Zt2�Q-?z�.�Y	�a�w��(w�]R���w�>y5m=H� ɤ>Ҷ58����Ƈ+��ݞN�"UJ,��`z����DG����2�L�S����㷢�� <J�%�3fJ�Ya�0~������_ 7���<��Fi�>�J�
(���SM¹wtiN�M�Zϸ�d��GffF�7z��!w���r�}�ݨ믊�e��εOC��ѳ�xd7�Mv�|�5|Dd�<`���	]L9�(�F�c�͕-ޒlL�<��DOZ
���'��_��Z 4}*ȉ�Hr�p��f�D��Zl�x�m�ւ���}�EJɽ��S3a�����`*B��p�:Ҷ� ^�}j��Ub�;>�z��4u!�~�[Hq=^ߘ	����9̇���d��RM���Vh�X@�(0s��1���S���.�A���&#�֯g�汝Lv��V��:��E򅓀��>����S%��(�L����XJ�駎.Ym�'�z����w8O�q��L`��޲��1c|�D�����"�\��ؗ�	�7���yߎ�M�ŵ�C!|�3�ba��:܍R�.�2�D*G��R7�TeC?�G$s����c��@xC[a�C{I��;�A�� ���U"�/���_I��a���ϦI��ʜ��po��<-}d