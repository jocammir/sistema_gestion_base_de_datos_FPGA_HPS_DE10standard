��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0����_���3e���ӌ,ne�	S�<\�i����B��wצl ���ŵ^qÍ��/�������c.�)��$�бl�k�*�TE�O�|�e*��#"!�X��Y?�D�T�<�����V�������\ ���𞴣
3E\Ӧ����[����j��/G�q��
�b��G]��=��/���/L���X��7����I��I)�:q?%$[<�����n?�-��:���r���w8���j�	E5�v����O�?�[�3a�#��?��2!�h��K*) �#�0З@�|��ɸ�F�J%O��m�	A) 3lp�ӀMB�X�`׋�]� ������@�0MB�$���:�p����L3�3&�|*)����pq���\�:{���c�x��;1��-XI�W����I!e�&�-9]���𭪙Z�d�����E��r�kL�$��#x��MU�[٧��ӑ�\s~m��3���x�.�v�aV�<X��  -d���L��$�%`A�c�:��7��4��He�w��E��a�&|TĶ��.��<�N�k�I�[qW'�^�L�̕���'d��7���yB`���F�bI47XQn�;Z2H>ڒE�ֳ��K�k�_��>;����M��k�PH�3�w���6n�3�\V=W#�^� ���'Q����W�82G3��s!sPa݊}^��`V���k�wM$�(J�a����9����� ,�@=^�w��Db�
6JJ�]��2�Ƴ��
���_��0g^��gH�#}1Nѐ,Ya=)��H$A��?�]g�C�����Rr9;�e_:s��a\^��@��ɯ����1@e�lg#�E&u#5�C*�ˢN�ՁЙC�l�J+��/Ϫ��8S��`�9=�Tc)b[��	��V�R���Ҿ�����s3!���q�i�bq>��F^�俾	}�霛D���iw�S�� a�,�}mP�K6���׬�����rX����[( ck�ǯa�0����;I���m�jkJ$N�I����M�z�׌I�$�7<~s7��w���ڰ�r�#O�Gh���]�dk}ަ�)�������w6_��<(L(Z��əa�eqNU䤡 ���r��ěA��Ʋ�.�蓛^$�@x���;V��j�$k5��p����m�I��sT�e�|�����'D5&�	���B�e͌�h����0-J���*Zc�i�ŞWro-hrBO��=Y���$�P�빩�>:-���׀��9^;�pz6�F'�����}z��ي�H�K�A�I�k�cD�a7!:{R5�� �4���v|]"�+u ��<|�_����!�ߜ�O���0L����6�?� K���^Tb�զ���}�U�$���E��/-�-@��ș܅_�G"�b��A�
r&Z����M�C��rF�qI������t#�����}�kC�J[]RK���Rm���: ��S7U��NfjP/�c�����Es�T�ҽ��-����,����1�p}|�i�Ez��-�m�N���?� �(R{{�y��t��u��T�k�}����+�7:h?������>��ڕr�WK�LD�2��9�^n�	�J���qAT�|<[�wO��9� f����dW�X�T�%�P<)$y�l��Jk�����(榧}�+��0����>>�G<O�}��@e�DZ%��I�8�V���0C4����w=�' D�t��pw%bY�!�3Me2B��c7�9ߔ^�J0T��$W��\���������v��|,U��#":�l�vC�ȟ�#�<�n�=~dHD��'4�q�Y�Dv_��U��I��������6�H��%5��4^ V�"x�K� ���Ш����@�0��N�I��脺UI��a�FMZjL�����'��ߕ&ȱ�(8��'݀�#��܂���&s�lț��9=̂�CM��$
��V�^6��o+�T��X�ɼ���z�z��6�.�9;�uY������˥�W۲��m�ir���a���{����~vN���-��Jg5�}v�������t���]6�d��
��� C�F�JD��޸Y<����f��?�*2���ι�2k7{����E~�Q,������:����ڶ3��o�IA���JD��ۀ����.�)�'H�������v�G�������������|XPk>�:K�	����v�9� ��j���${��_�a��ծn�C��-�b��t��=K t������Z�:�i4ݮ��q��j,�M5ǎ��&�)��hi!��Rp�H%B4h���C%�B���m^�u�������G�6�F�Aeޘ}�yztVު�x��W�� 3������ �T4XF4�S�q��t�"��a�2�/�U���ul��6���v �$S<3��}:y���xm;������S)L��&�B5K�r��ӧT�E�*}+�7�'�+�4<RQ���gk��ټL!�����o��zh�(»�3� yG��gr�"W�:d�Z���cg�yH�	�I8[_3�U! g3��};�*桩B���9T���lګ�ۣ0��[c��oK���q\k	;®����I&���:A�t?;#��#���`I_�1�T鐙ǯf�����^���펛8.�7����v�-��h�SlP͓�eD&�bZ�#�"x� ɔ*6	(%�~B1���X3��s�6[��cy���p4�(e5���M¥T�M9��LVr�t(�����X;�]<�ވi?�N�O3��ւx�7D �᷄�5�|Fl������/|��:o���)�_=M�K�G�Ce����x��X��t�bu~%���p2��{��!@
	����5�Ѣ�N� ���!p��,��)h֎�~��YZ�ߖ��-5	�5���������>z����b%-+'Q��3M�O�/�R��U�L01���֕�|5a�#j�Æ
{?�)&}��ܭ�EY7qK���q�g����2�/᳄�B[�����>H'����ڱ������Z�u�El֋�����8�}`i��y���q&HH+r�,� ~��59��"T���Dv{M�i>�,�rv�)I�Z��%�a���BCO=�o(���9�ʉN�Q�?\S�@���^NE�J�B�(���{
2� ���SϏ�Q�𲧿�l��emy4�I��ǀ R�|��(���t���+,	
I���z�=#a5`����Xn?���$��2oLO}��Yf+P�XL�L�]׼��@�CA�Y{I�z4�e;f�b�ֆ\5�8����D�bKc�Mv��kS��W6�8�x>�YAW
*��N���On5�mW���+{R$�4��%��W���pn�E�F�v�p���TJkj�֟��)�@�&I�O���qo����TFx/�D峺�j�_-yJ��� ��R�A-;K�G���gc�( ps����*���5��nh���d~;�>��/mw��cT����z�d26�ޕ�����9c3ʿU,4�`!ޛ��S\��+@)w��2z��g�(��f��A$A�X���q��M[<*(xz���]�Q�f�d�hŔHy��D�K#A%}|%�)p�i��0|v�	�чay�G��W��
��;��]D�(�_��"����?�����en;ך�����$�w�*I$��-��2�[�{��Bf���F5&gO�ђ1(Y��M?/�c���d���&pn-��T>,�����"��R#G?!��J�)��RRǄ��iJ7(pS�CmW�/�~;n�	�Q��O�q��"��U�.zq-��2�{���=��^ ��g�ۿt��W9�ܔ�Fa��>��F@�~;�0cٜq����n� �Q�b�;�(Os�9�[gf��fr]��rFn�� ��Dtt�L�o��s���������V˝<茱0R�y�D	z�k���@��0JN�˽=������xN�I]�����eC%�D	�p�ܾ�r���m��G;�Z���b�Y����ЃH�W!�7��,���%;��?����I�~_9����h�����j�e�@-O�r�����1�A�Q�E���
ܹ_�s�"�wFQ#'�\T��\��,�p��9�T�}[��+���r_�M,�h�Z����x5�*�v���1%n���E�U�
IֲF�8s� �(ݻ �m��p���ѡ�zO&b��(�W)�Jp��UE޺l�����ǲ���f�t��y�w�0�a��n2X�<1�ɗ����5^g�h3��&II�0�*���dɌ����W��a���̧7�p��n�#��޹ +f����g[IO�mvu�`ԃ2����ڻ�;���a̙ʾ�����|s' Gjrq�s�� �i:c�A��j�N�$�$Z�b�AW6�h�u
����&�հ�~���a7�@C^�D�3@)�J�V)a�fqu��tI�� E.�9!.Eq7c�~�&`.�:*"1U{�h�4[�.�55
�A��hW�q���<b�o��ߖ��J�@��7]�h��n4�B��\�r��B�3�JL6�׿�9���.SY�"�w�\��e��[�.L��Y�V2����Q±��!����)��]7�%��ӯ1-t��0	��J~ Čj��VE������ŷg;�{2 ����>���uB<	8��������a�>8�Pȵ�r�~3���:���,�2�-�����trQ�徂Q�Ii _�ud�ucr������b��E��L�Tl|OAh%�
+'�&D�vyB&����.K�mQ�<���whfZ����2aq-YFb$�\:�@H��#�(ʁ�n�_e���aqL{L?���˂�Q�[ﴉ���63��;�3Վ/?��Rv�1�����ɭ�����$v痯�D���+\�gseB	~V�	�K�ԹMH��x�+1����0�͟��R��7�#|5Y�����ed `?
���D���P�C�� ��<nV;�:�?��d�V�Z���g���}蚂#UYٝ��_�����6�Ed���=�Ą�{c)\E�Wi����p?�I���$�b�r_{��r"�p9P� ���95F�5EC��ϐ�t��RX������dՉ[2L���3�u�~����lY�-F�Ia�>���/�W�kK�hOy̡��L�(�Yމw�*;��'A��!;�Q����d�|�Յ�]bN,P4R�\�[�@���~7����cp���er}K���י)	�H���8T�3s����ô�z+7�-��Aq�O(C90�Ul4I��4���y>� �6��Dlڗ�BC���q�'�apq�7�UA���`��O#7�	�Ïd���Jm)v9⑘�n}Y��{F��Ӊ�g�wt�ݓ���y����nB|��ƍ��Q0�_�cj"�=�qg�2!�tM��Y=VY�l�(�a�U���s,\�J��e���UaϺ��ϷJU)��ܭ��A�^�U*��p��k��C{�� �㉣c(�
TG�p)��^���u�(Yh�NT4э����I<շs�b�+�&v%~s2���6�$��dgc��� �v<y�&X����}�n�t֮5t.��@�M�OT
92����;�+�#U�Jz��zP�k�+@͕1ö�@6�9k��ٵpԯ�ZP���M�-�Z;�2G�ͺ��c�V�����$z���oNT�.(y
X2���LQag�����:�E��&���� ��w���"(bZ����`6�*;�y:ʏ������V�`L�47t�����9�c�^.�A)�tPI�tR�Th��\uG�����-c{i6u�L�{r��j�.�%��HD��3`]n�j[*�p�:A�;�FΨY���B+��,�5�p������D�vs�)cad0�Q`��%��
܀O'�h%2����oԽ���*��Ϫ�g�:�V���<�Nr�s����cD��u���{��[�T��@����c�
��\DvY��ϳ���o��-r.��\#�q��q�+�2�l��w�j��w�D�4H�7*�Tw�z����IH[�h��t���T('߉������c����*O+�˧n�/rI)�-��+Y�&�Ȍ(%��1�/���X�˃�]�������8�rq��bGM�Y/|��ޜ����!��N'ӌa� i�v�g���C��5{�s63��y�sK9�
EP�&v�����9�N�o��	K��La�^�m	n�*� �^N*��e�b5��s���E/2�7�c�&��Q��Q���jڑ���Cl������	�T��
�6,��U$({/ӷw��
��8z�*w�%$�������g�T�1�ϱ�U�u}Q
����o � 59J�7�M�m}Ov���Y�z5�C��`���h�sA�`Xd��v�
!���L0˭�9�	!r���l��(\LP�F��:I�1+Ul�"xAz'C��إ߭�B.R�4�Үk;����߰�$�:�`�|�7��r�(�P��g�1���t#}�/05Գ(�G�|� �p���j�Y��הs	5��� ��FU5i��0O���JN����5�<�$#?|x!�_-�,-TE��#�c(�azPO��ʢ�$h��ӣԱF�x̙Ac6�˃�,-�����X��a Ń��.����٩�� ����fQ^��D8)f�����S3�p�G|��4!�^�5�Z�<��p�*FPp�s��l�H�P���Y�&2�!=!Qٱt����܈�Kq�}S��d����[������ �:��E��\v��ش�J��P���]m6q�����=}�`�Gv4�h�EDje�A_�b�֢�];N�~�}a�@���U~!�g�}ӦS��=N����X֍��;)!3QCI��&>�����f82ݎ�^��cH�M�oA�E���Et��Zuޝ���5�����#���iVӚ4}���� �>&���)�_k��l��<�3�A1~����{J��F:�\� �"���1�4��wA-׉+�όn�� !(�����q
}�$B�nNhf�1�sI�y�W���)&~x�z���?x���`5 �����Dn�R�
�4�r�{V�2�t��\8��H{�?�D����nE��b��M��/�����*�s�G	�yHS�fI��E�H�x�^�5�B�s�|���2t[��H�It4�+A��Q�[K��,�=:д4��uiC}�^��#��SL�s�?{�sJ�I7�jM9�4�	��(��ھa�,T��Q����݊�������m���rMVXB���fwA�����꭪���"�uAb=��r��A�!t_u�3�C5���(/Ǫ��j�<p�N)�� )q)U���c�ޠ5� ���G�:�1��ӠP���r
�J-�O_���[A��6tJ漘�%�c�����Hy�K��_������;N�S	���P�$����:% u�����	=�j+?	殺P=�r��'���~��_i��q�&�8���l�0L|�1��w�yQ��^>��Ys`ٓ��z��3�EP��Ku����GHn�ȱ��y����?��l�A�H���g��^�j�o�Z�/�^=�� Ў��CH�`Tuv�k��+�A7.KȪ������Y�r�c����h��9�� �����Эa�_��/ͱ�R=<���쀩�4�䁜���h*F�-�.���3��V[{���<�r�)^8 D>�piE��.28�Q��&T��x�f^��F��E�_���CO��dh�Q^�!1�-�����[/�>ip� ]BǤe2|������S���rE��y`3<�K��=Xŷ;볿,���YD�H�/��/�q�&ZmKT�BDQJ2K���~�?�UZؽ�rz`o�ųC�r]����������v���F�/�P�ǉCO�8bH�N�+
@�d̐�=XЬ:��=ml2�Z���(��B�<����$�-BS�P�## ���Y����m���u�[j�I��i�]t!E�^:��g��?c�㸱��7�P��>,����ϻ`nj���3$�
��W�9�N���~�H�O}�A�H�`�@�E2:!�)�[���;�_	�l�at+Zq�s�
|F��h	�L�;�Y��TA��;%7}��	 ��G�ý�;�Z��34�E5=���2熀r�3<����5��4<��'�m�|��~I�t1�ƿ8���_�T�6Ee`qO��w%��r~�`
�[.�R2���ƍ��Hğ���A�2+h��j�A@���_";H@��o�ut�8>��H*%y��@����U-81��x�l����O�-d����>��3�˻:
ZF�
↮�~�C|Ka<�҇V#�7Z�/EFeѩN��C>.Jr�$�R']p濓����b׆�H�e��f�10��i��|���xH/��6����1��	e�<?~��.{	�oEP6��4�0R��������wם�f+9����"E�L�=� cX}���O��%�L����A�jJ<�#0�V5���k�'s`��ä�u�m�e�q�}+��P&|V�	��5^0�B�N�ͻ:�-��ĊEV����V�:F߾���Cv��2���?�_z!W�M��E���l8\��a(y���w���&Cl��'9���gܢ�������v
�����E�4�g���w�?	�˰�7����A{���t��rH�Ѵ
��2l����ߢ?���p�"�>ps�]U�&9�� s B�� Th���m�3��)�9zI�nQ�{�+���:���(󜥉�E��
�S�!�_�祊�>}��j]���җ.��ZF��Ob��2�qtƸ3�p�MJ��'Eۮ�yo�I��e�#Y+�0�k���r���z�7�O� AOcWq^Rr8sj��#s#F91t�Tگ	�}���p�FǚPud��Ţ��z~�p��>]�8�3Pj���dx �U��?�v��iQ��)���`#)^���FTl6�1	����A��t��,wL�&����3y��u�2Z��<��]Cu�:1�d�b�w� ����rU��w���Is,�6�΂/����_�KlfB�WB����P]#),בi��8$)'�q6�i={���p�K���/��i���C��O~�`�ѵ����wR��W��4���4��\%��|�n��~##h���@L�Mq1��6�TP��w�M� ӷ��D��Ǹ�����6ޭ&Е�_X~� ھG7&�w�ݾ4\�+�cU��R'd�qaK6�h��fqo�hLTwh4y�'\��m�+H���LhN���פ�0����I;'��O���	q@��KO���Z
�L��A)�����0Q��Ȝ�w�#�q#P�)����� ��Q58��-�������
��~z2�;��F����$�Gb�eݙEN��̼8ABٜB���lJj�!EE.f�1������qěہЩ�����K`;���6<ܣ/"��Rh�=�>L�p��A�K'AP �V�J��AUW��-S��~Ak���T=�)�ai��E���ߓ.�������_��IP9�%���LW3{�^�����V/�A��/��J�u�oirkC�'���΢�y�#�^~g�w�t�f��/wP�o�pl�FC���
H�uNT�N�%]0���wm��iĢ#f�"?�y�di����}̻��A�Bn;��J��.�a	8����rr�d����������g�2�74K�)p�a���\��G�����Cm,x�mk����-����YS�/�����A+��Q�݉6����\dA�x\�m�?����n��߮��c��_�C����X�!X��u]]^��~µ�v%A"��n�_1��Hh��c�������V�rI�e,��b���m�z�PME��E���&�Z.�b��~�^��(�����y?�_����~��W;��X����ˤA�������G��f����5H��O�~���Q��≜�n��Rrho��R@��M��Q�+Xf����)Z�]���ʹ�����a'�Y��A����y�F��d�=�����9�d����s�0&��?��)���ϝ�~�t�����2�߳�T�n������r���0|�����Tƚi��$���20�k�Ò�U.l�rv� l9� ya&� �'{�J�� ��|<wn_����͵�u�#Yd$�|�*�N��#��yx��`�:�h����(�Һ{���	�4Ɓ'U�d��(�Y�C@��46bY$%��DIt���{&���D�F�g'���<e�u4$YXK",j�.L���Q!��8�������dĜt9���Uzf7i�R����>���*���7
�/�\��s�argͯ�s��?���Z�"<�����鄖KW����\�N7�