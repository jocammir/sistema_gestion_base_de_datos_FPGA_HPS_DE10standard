��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�s^W���0A	�.�P��z�w���U���\��لx�9����og��O	\$�Y�A�v~�5) �M���4Z�2�^�g� Ӧ�"~`�즨��i��N+��	��5�PQ,#�M�b�/�j(2Y�dg���a�=�J�l��M�e.�'�BZ�v�b���.�Zu^��'���
Du@�FJ0*}�F�;��ű��H�U�tܖ��^濜l��Cm��(��<ԏ	���늾ZvF٩rȇ-�f�o�MZ��ւ{yc<V�b�Ș�6+t��OMli�(hKox�P�ߺ�vB��D[mPB-8</ي[�ҽ����.�N�i�O�,��0�$��T^�>C#l[�.ɓ��^�N�-k���C����%Z%�Ӈ���`����v?��J�Ĥ�A���17���l���7����@x��ؐ�^��f�놖�
[k^��%=���A;�eǵ�S�#�9�����϶'n�&Ң����ڠ�����A��h����<F׵j��4<;���=��{���2î&=N�Ru����a�|��^�&גo�,dN�ș�(�1�X�u�o�����O��s3�f��,oV��lׄ?q��f�.�#��m ��N@ϑ	VcȔ�25�����>UJ�l���ݽ�LWI�'��4+���Y�y_I��G:��]Ƨ��b����~m��OJN��:�a��i"��
u�yu� ��7�����R�,(����=���j[%��N�VF*���Ԁ�Z��nWq�LwK,x�R��
!'�T��fC�"�Wc�뼳��O��y�
��pʗI���%7F6�N״�9���D��������z*ӏ+f�G|�����4�>�q��l��0e�V|`���]��k}�W4�>ÒEWU�l��Z�hR� o�)6�22��&��u� ��ɰr�Оꄵ��5��=��f-�d*�����yJ�6wꗦi$�~�&C�(p�@
W�G��_���]���DE��0�I>#v9�y��T"�~y���yRn��
�$��jdl�6�<����7��-�C/��]n���p'|��Ρ���!�*X�6}���9$t'�6�,A��\{�iRJ�t2F�U�d洊I�,Ǒ@�/�_}��,�.0n��@��8���%�l��Hc�7=�)�~�K!��dG<��e>�]Z�3��%뤮���FS��Q� �������	y1;�p���o�ČI�M�t(pf&���ǐ�e2Bz��c��FV�l��هF���N�.��m��6Bj�/�ٺ�*���A|��nb�U������7_���v`�Y�&
(�ՁE�fm��*U��9�(=��e���܍1!j��m�1'� �� uYE��S)���ɱ�����@���͖?���盇ݖ}-&�#�8r���=����H二��BMCI�S?=�J^��:����/ڶR��1[*5��#w,=�3�m��wA�M�/q�gi�W�#)�*�뷕1��*/���K*@��*]�����[y��⟘:�}fD���W\d�Uj�ñ��ӁE�k�G8V��{{&�)q�H�><�Ɗ���o���6t'�5.�~�x��!�ŨcK��(�p���T{1Ț��������ʹ�]���Q��dp,�U��=��uD�n婮<��ݑ���&[����y��'�<%��dZ�e첯�}�X��4��{=�0���4�lN�ho� ��'IWx���P�|�+�F�֚�ћ^ӡ�!�|ע���J"�Jԝťyzq7�����d�j�<i�������2j��%�1�ΰ*����`���� ���l鷈\j�p䧔���)��vn-��&Shy��Y{�-1��!R�����`\������$y]�0*nt��%˕)w�;M�L`Qk��-]f���h��D�A����p��v��&͆:I'�}F,Ba��Z槌2HZ��\4�cUyۺ�N� ��J���'i���RC��AUV�� ]�u��w��^�Ҥ���=?�a���U.�o.���S�-pX<�`��]տ����$t`�I1Z��?�wP9��QN���P�0fZ?d�ǉ�a�U�D�S���k+;�Ͻ�/����׮]��K: _�Y8O�6߃hBR%S9&'ژ/�ɛ{/-2>�s������{��'<���񤕄�q�|���b��	H_M;��<fVy!H�E�s��EI��f{�8	Z-܋�V���m2��N�qт~9�]�\}�c,�$���ޣBy./�F�r�6wb�����meJ@�z��r�ϯ�Y�x��D%ΚE�i��}΂{Kp=��2b����o�������׷�؎32pcj؂s���@�����iY�<�q�#2�g��A�.4�3���b�R��k� �S����ֵi*}C��[��{������gc�HR�% 2��4�L��Ӎ7�T���M�0��yr��c ��߈��J����L�8&	�$Ŕ��ֺ�#e���Xη��FӋ
9�@.�i�dI ��9ڞ-%�
>"��[�z�e��[w��Z.���y�zS "�q&@��AT?�ߎ5���Q|�P���D��W����c�Ӂ�d�n�'�;�r�5)-/�}�'�x�]ADD�;��S1*�����s�@"JO�� u` `���f��"���/2Ot�Var�� `�Ѧ΢�~�N��)D2�'�p�~����@b��>��8�y���6���S^���.�[3�Z�c鬂�i�4i�t��]�����^o � h�LI+�m��0Z��_)�����U?����Ek}�Ǽ�2�v ��*�:�7j��L�Rhf,�k�˘�xg86�ر{�7}�/�.h{�f@4�2-#�_^}AD���h�]b�Si�dnR��,ŷ^3ޱ�S�{Krhq����&w֬��
�N�֤r���<��p��.b��g�i��p�>@ϭ��W7t��Yv>L��TS��G8힥���6� �43�VQQ%sY�ۦ�O�����Jj	8i�ب���)��֌-�<����@{�J�<4��Bj�`�ϜR����G�u���탷{J� ۴=���Ҩ�ֈ�8`g�5�W�l��C�Djv��p7>���e��z�5q1KS���Cw�����|��*] X�:x��J6jP�ns�NLkj=O�$-`�f�À�5$��h�/]u�"�`��L����ӡ��q4��ՙ��B���W���lQ_dnO�ߤo�LO ����$�C��h���{���UF..����A+udB��|��y�Whh�t$�����v��<��1#1����5Z�-,���!Wᷞ���a�rP�����ĵ�z��.��^���^�S�۶�(�X��3��$(���q~�7��}�N\�H�m���9� ��x^�8���Y�_���Թ��"N�Z�<]��Rk���7�#G.Kp��2��kː�Z_~�]F����C���K��	����"�b��<�͂�u?�����+���0V���4���?v+ũp�q����$��Rq��P�J(˪Vs�@�F6��F��^Vv%V�ȹe챡`��?�MB�����U�c|��;F@����~���v�"M���Dg4Q<?�5�P��K�lDIn](U���2�,�
�罈�����$	H�OHT݅�v:�_��[^�xֺ�1M����x��*)v�5�<'�cTaKΐIa8�-�C�v���M�x�ڭ����u)�!K�t�S�P�n��"�-�&�ņOn^yP��~T��`��/��!j=u�l4Z��+��-Ь���A/��^THk˧<V$����C]��̘bQ����I��w�� �%�T��g��:��5˪,9f^�����vƾ/��)$�}���%(������g��X����y2��B�G�X��w�j�e�a��Q�W�Il��e%����B�\���X;��,L�H(W�J�5Nt��Di.��n����v�[�#	���%b���gmEbe�P�Г�:���57手�S2��0_tɫu#��7���A�A! p_p�����()-�j �VUA�'!�/�D���}�Q����w�|��I���癿���I�6�V��N� �ϐS�iɥa���*�&l��^=�s,1'�R``[T�:N��2�jC�H�o�4thHno�+�v�տʍk>� 9uj���p��y��2�"׹�8�.~O��k��Ia�I����pR���5�o�~f1b�f B����v
��E�*Q�;\���x*.�*�|�$����k�{]@;������>#)Pc!6_�U�ԥd�Ó�.׏��K��+2i��.�H/K}\rǍ�h�>��_2Y]�5lH�ܼ:hY.zXk�4����a�}��è-h���(iLH�{n$�!�)�Op�o��Y*}F�ʊ�R0��7	��nYy�yI��Zb��U���1��IiUΰ�|��ư��a�������>x]?�d\PL����ˇ����=���*�����(]��r_몭����^�l�XQGM�ر�6�r���oV�c�>=&d~�����	-�b&Td�67K%[�Yaj#�N1Z�a��Y�P9��]�1��X��eJm}R��۵S�E�����y�sp" �ł�H-�Ķ|.3�p$���:��x�`�
kLc����%Q�@��=b���g�J jI8_Sס����U��_�K����[��K�̱�[�B�� U��k�"�L"�5g0�̶ F�wP�QΫ�r�36�_��^�af�����9�#���|��S5�^�y,wm��J����x�P��A��?��,0ѓ+�6Q�3��Ȣˇ���.gzV\,]���]���lF�����k���26��xcL��٧.�RY��O��1!����>�F����A�%����qV����iC��;@�蘧�!�����%�V��9��_lf�i���T_���yXP���s��& ���E3�N�2����?���d1ߐ\��A*"m�T�����G]����29�jK���Y!q�ij�������G�Q��S��i�BR��pnЯ�
��$�����Uf]8'	�R�R=2j=���P�@��^H������"oWXu#��?��ČWi���,��kvha՛���B��t�q����*.�PXO}��&L����!��+_&�Nz2�`��O��v��h��NO9�����7�\��ׄ�����cW+�Dvg@������6X����T:���y�3H�1�x�M�X��w1~L��:�D ?I��7ׄ�y��[g��K�\��(�a���L��U�'�p������\��J�k���w����#�X�<��<z�qa��1��N2G{�{����1a�������]K�C<�;�A��/���R�?ь|q��ҩlE�G"q�N_�tg9)"�����#ߴ"�:U�	%�Z+���1b��B�ɼS�\�k��m�.�Q�xܔ8�1|W���$F����FDT������_z!C��~��H�՜@�5]r.�9tT'kg�f��"=�v9�0�G�Ȍ5��4�]+�Q���G'o�O/����	jm?'OPD�t��aG4Ĉ4U˩���:�S�Aw u�m���"u�{<aU��J�](7H�_nآ!�g�{�e��Q"pe�i���U��,���U�����W0�0�b��͆l�A6*f�K@N�o6$Cn�l<�\b� �, ��Z�#�}��Q�w��Y�
E�����}��#�¶��tX�?���?�2]�����a����X�EM�707Ƞ7�&{y;�Q��)ɶͨ��&�⠀EAk���v�	]gRAg�02`ʉ7�/�^t�+e���ކ��&�/��#�ٰ��
E�ܥ:��9V�����p�J�I�f�ښ��.(|
"�/z�"�SH`�S�,ۤ䔞�_��� �.�Ld��ԏ:��ġc.�)"����A�g?�7m�{�B��Im ��{)���@Q�/��".=ތ�`���!�#r�fc.�j�uoc�N�>�B������lqЃx4r��7������^�I�γ�xV�⏕
~�3�;;zE*&�������J����J������2��A�� ��U|��G#�v�\�lpf	��췤0mC�iWͭ�DC,*��#}.9�?'4@k��P��?�R���+�sJ���$$�d�]��UG���b�1��Vc	�b0U=VIU����:r�ZD���{���
�a��aY��ԡC�gз9I�%X��/�lC�!�٦�ALN�X�8��=f�vVO2��h��{Ϣ����,�#�Y�[.kj���Ēi�/7��.��.�ɸ=��		4Dt+��	��=�d�ck�#Q+pλ��S�[�ʿ�}R`&L��۟�8�3|M,ۡ��K�6��F�Ҍ6��9��C?�.�di�&���1�PS<[TO�'N����B~�\*�e �q�^p&z9�D�A:�X������J�y��'�rfKC��x��tqa�O��ݺ\�^��gxF�\���(DV����ܮ]�u��gf�A��.����+ft��wN�8	h�|FϨsjbnD&E(!w]Ȋ������>Ж�������4�Pt��\��2����S�������t��A�]��`�J�p���!�QaC�Lc��\t�VAe��Z	��av��lJFY��Z�ؤ�5�����ߪ�=D�X�vE���l�7GI�2;a��]��h j�Io�-����>��(�㐪���
����'��o�(�ؙ�=:��q<\����ъ��/�����[�O0�X�M��5�
�pMC	���
�$T��0�B���˭|⇡;p6|��c��Y��P���"��c+v���<܅}��3�j0���I��5X�� S���/)9˅SJ<�oz]Y��8,W0��8gz�tj̜�;"�_3�$j&�}i5�L�̔纸�Pҥ2D�;NL�Ge�C9��7�༦�#[`b^���/�� ����e���t%C]}i��t�-E7Ug�X��6���Ak�
�z ���"q�)Agꮪ-f� g3��TU%�����z�A�jV�{\��Ԡ����L�]��[���<�M�9����,�cb?-U0�݌}�ݣ/�Еa��~���K�0�S��˖�
���r��Mi�=�˅���y9�Mi���?����y+s�,�9Z	j��!�#�%o��;���=\��uEx��x4+留�4��NPoΗħdwo��섒y�{}[�Aq��4�(l�:���g;�>K���e��m7�<��a'�A3�ي�U�kI67�r�.Qό�Xq%�fa);��tƺz���s�uڴ�:b��v���z��՝�o�y2�XS����P3��cF�W���ۭt˝M|b'%��O�qh��mc�A�5�A)�V%���֜:��� �H?�B-A �0��wSa?�h71��+�|,��VO`X-aB��T�8/��5���Y�PL�k5��Z3���=)�BrQԬ:~��.�^�q�����`J��j[ur
����[�c.i��OQ��!��
�ۊ��XG�#�W�T���P��6������jn����/����M��H��@����R=�PB?�r0�Q4و�U'�hٜ{A�i�pf��+�Úox�=��"S��p�k�>=Z�HC��
崗M�������ꩈ%�L��3����_�潴=hzz	��D��*�W��Y��XZ�o}v6���@Ne҉z�����D(��プ~M�����cM�e�d$� �#����q��?�jtJ4i~���jn�luz����g�A_�����"��/=s��!~�)���p��������I��Y�ST��;�u��������O^���4���Í;�8��r�e��9DðQ.��X�T��cU����H"����D(������)c�r�0�TsSs9i7F���g��&%7dh
�́�^!��߹���~����*#�K����e��Xƾv?/�}�<�0䢇���-��f��fV�S�s��e��C{NV�<Cքu���n�Ȩ5.}�Uk2�jK7d��%R��08M�S�gM0N���brߎ<��aV�$]��BE��w[�L�6�w\�w��"Q�u�/2�U�6��:��-��kB-���B�J��!;�KV��
M��ꏡ,�hi���a]A�z�mؕ��Vq�"����mbZz7��̈�j�9��滽9%%]�2��ZK0�e����3q��ݓ���~o3988����^2�k~)h�2/:-è�����(.��&z+�#���N�S��5:���+H;�7�ͯ^.5(�'\Dʬq��i�h�]��i��:%��N~6�'�i�����AE#�5��rw�lᜄ9�V[:�a#ф��җx�XlϏ��zI�P�N��EE_2�D���ùp�Z_ym������I2F�*�?�H��x9��)�4�Y�[� ����K��[L�`��$�����߸R�V>T�P�	�C�w�y�Xh�Z�ޡ7+�����-;+��F�1q6�"ƨ7n&��̥�\���1�몬��E�EK�;��v^�pĸ�3�%C�g(�Y��,�o�`���Ƽ�]�a;e6M(�����s'�O�dA���P���U�	gz��B�\��m\���T��� �\��N2ٝ���tG�����@B{h�6���w$K�|�����@uE��f%��f)����|��i���f���?G"���5L�G`)��B,B���`�m�9i�vH߰0�F�x]e�[h������T�=�=����s[�F�ޞ'��/����e�H �x6o���4�r�52�I?7%��-xc�p�	B���toqpYo9G-Sp��`'U�c���;���@���W�g��b�V�iS���Y-F��~S���A�����"mY��}����<Jܒ�B���. %��me����zZf>��������W��_֗�X���{�r�k.]b�f�����^�N��$���\���d����'���.��F��q{��v Ufx�;F��ɲڧ[��� �"'��E��1�,.�9��(�E����[��:C7��m��,
���g���E�=�����?h��G�q�Ϊ��cw�v����?��k&�\I�cۙ.ԗ��b@A���IF�Rѹ�.�H��aȨC-S["��_r_�;*nQ�j~��%�<l��Bȭ�'���L	St}8�i����o�	�@S��G��R��V\�f1�q�ċ�lԞջ��ߦ\�����������Q6}���D��jħ���L�-��/}��l!iT,!�eYf�~#���6�Y�Z��SO�b���(.�����S��Xw8=e� �Mȱ���֜X��Q�'�!
#K�=[c�h�&U���!���( u8q
ew>��?��ryԦ����[�ң��$-'���Z��3T9p�'E"���#@�����K�@a��R`}�P���ejJ06־AO�];��l�Q<���e�p{�+� �?�64.rl��5�Xȃ6������D�6�d^��s�&�db�K�Ç��t��%@#���@ڛo�E�QY�f��'a��'�7��֮����K������HFk Pjcek�8х��:�aX��r��Ga��Ð=��j��C��ʤdF@�t��V��o;�y�*C��!N�{&(����Ӵ�£��SH<7.��@[/��h��4�:�`"��T��3|y^C���g��s&{��~��X�G�Y���Nߏ�u��F* ��#�7��ݽ�K��8Ǎ�1�;|�{��u�Ч~���q�[`�=SD8<מ��A�,����c�D!P�gf�5ڥ�3\���P�tK��~�:Pq���C69%��U��	9S �-|�	pi��]��*yQr~�y�׼9͆�x�dK��n�l�&$�Y"��,1��"µ�GJ6��z��L4[�֗b��|x��@��F!��d9ԽF�� ��3�%oLmF�����Ѭ�,:ϽDY�����ƚ�;��RX1{�5u��=v՟w!Xa���o�/)-v.3k1��Όo�7��M��&9��\�����t�H�V�M0��W��f3u*�d���������,8I���Pr%�Jk�)Q:�g-���l���-��ˁ)sM_b��GD�b�2�tz��@������Ư)v����ى�׺�r!MJ�әv�ɂl,@<��^�쐇��j�\������H��<2��O� ��2�� d�D��5��!���ʸ7��i?�8uL{�!���N����Eb�	Z;�ۄ��f/M����Q[��<4�4	��Ȋ�����&�~I��U�z��_!GM�)qMAߠ3̄��!s_e��A�z��A�Jݓ^��O�G����[.r�;����hV=N�M�U�#��L�߰~K���t%ې�����6qB���W��Ye��sh���1�4eKbBIX�����V��:�IY�b�G�d��	��Ēc�uw`_5B"�)�q��_�����ZxR�ߵ��`��C��Bj�?�^{Z�h3�����Pq�)���I�2WP}O��-Z�HQ����D��s���WD2���|N-��<�V�p=~���f�.�B׭ݫ
QQD���^�T<^	i��ϛ\��V~�)T�Q�� H��4����y�}�����P1۸at���˔�=��;BPM���#���E�]?�����)�ѳ�����!��[�B�O!2[3�v/����qt���&��
O�Kt��_���$m4é;���ه�e�U�y�،�������O�[�s@�>x�*$ׯ����Mx��O]��b2�YwkOs�)����k��>�d�#�J��Do��f������l�l�����*K��� (��j�\��Y_gCX�t� ���t�<R�QJ�GMXu��f�JH�e�K��t@p���D�����w�Z�z��FA�	�_�=���(H5RR�6֧+w�+'���T���s�����_e�)��NF�+x�����@e��"�H�7���MAB�jQ�C�8��� ���.㹟sO�XqpV�kS��Qn
='�S�m�v˦�!q���M@Y�鸹���{r0d�5�=  �w�PTF����P�+�}w9�:F����  �#q`�i��CP�C3��Q�&\��s���6����o�/��%k_�����u3X�r��(�}����\xR �L�^\��"����;�ԩ�[G��t�@;�����P!f_,�����_�x1׾\����� ��?S7k�2��f)��ZC�"�����6�HYS@�����
��o��e�[&�dJ�:���F��͓�ؾ�Ɔ���<aڣ�Z`���e�^=��������\\��o�+�.:���/�6��dI9��I�o("P�aEp�H��[\��Е뭀e�������Ѽ*l~oֲJ���
ij��P�P��O���Q��А��</"�Y�\|���;��R�,�ρ�	��L�<ցuV�d�	I�v4�Z�Qd���&� �G}����%�W�����$%�6�o��)�Yo��?Cq��|����	��م���$�x�|��7�j���X� #>���ހ=�Y ��G���{�E%��|����pea	c�b�ɒ%E����u���c#/�ՐO�a���;1R��!r&�%c��x��`l)����k���K5�f�)[��R�'�:�ɿ��p����tܬV������刺qB�������{s�X�N��K����;����^Ov>�3S�
���(Bvk�j���mJ�a�G��w:�!A��"榳x�-AGw2���+���J��y�Y7X)�]���G�rn��zgl��_Y\��1��a^7h��m��)���P%���車���(b��"s)���U�P�XɳvQ����@���?�*> �[f�CGM��P�~��ԋ�R?�8Y��|˖<ofi��5�+��S���u���JOo������i�>�x`����N+��֯ט��)�^y��ث�$nձ+`�F��˷X�F$[�A�p>&[|�		�D;)g��V� ��"v�fel]��\)�U\�χ;[R��; ��L������QQ�lx_�[�
���-�E|?�/�I�s�N��Pm���7�}=NZE�:f"Au0-+?a��^�?щ�7���G����K(�������X��1�Q0�1;�E�=��8l�y��n^�� �4�1�?��.�1��D��9P[h�������2+���E��mS
��h��d��8oY�� yԒW��^��A����NS[uN;��6��PQ~�%��s`�g>rt��&���L�λ^h�B�����\�Cw�n����.�Bj�R��mk������o&̓;^L�>�Q����!Ɇ��ϙ�~�$�>|�W$W�����9o�
�Y(:�#���S�r�!�k4u�H�
�a�8z��Cnk7�>e��A�/2L�p�}�x�$L����#&���J�§��^)oS,�O����������2��:�*�⬊�i�����+�N{�݅J0���#��X?���j�4�V���{�!ze��N(c����x`̢�,��t�/s�u�bW�z�+��.��F1�"�Q^ٿ�}H+z�N�2�y����xdu�ַ��ߟ�]7 IjŴYj+�C2s�n����Ԡ��A���v`$����}�(jD�
���p�����uX�3/���YY(.Kw�n%��W����K7�!�U*^5��L����g֙���I�Q���&�����G����B]b/껮Q��ԫ�mz�S�)5B��?ēy��&��(�����%M�2�J���74Mt�%������ [��G�Hڑ�C�ii��RR���`R2�7K��B\�$�F��j�mM$��q��W���{�"��<���9���:��F��������U~��*�+c*�`GR.1��OV�v��5����I�˳�J>�~�7m����Az�c����6��ݲ�� ��*SLp�[ҍ-}E�V���	���Ħ�#[�,EE��ϛ���x�sx&K�҅����<�~{����2�<��/g�}�ͦ��}Twm��x-w��o\>���$#E�|�o4��G �W�*MR
�yu'�~r���`J�'�e��꘏�<�M�+e� �o��X�x5&Р�vR��������.�ϣτ���V�����U����Ale�q�}Z�7�t���  r��[����-3����ĩ�2B�kʡX�D6�K���	?M��ݗf�U��%�r�~����Ð���x�k�:۫�7��kL�6�a>2���I����®}>�P8�۔���`���/S�������:σ��&'���-R*���k�O'GC���� �,8a���!R$߬���Ř�;�ң4t����X�uh]1�q`(��a�<�Y�+��\X^�Yi���R#��g,�/��aǌ7@*�<ؼc�iv���~�K�V \��62^?�l�f���Ć��p0܇�kgS�0Z����Cww't@gU.K�ʈ��d'���E���C�/�-bbhU�vl"�˕fO��^ϖ6 �?�g�n�3f6+���-���H���(���Df��)Α����nFKԞ9���Q�k}���Ҕ�]��^P�������B����[ua� ��ãE7�����k��2�h����D�[V�^�ˤr�f�SxP��"��]��3uR��Ec�,լ���*T�4G�h�
j��Њ��p6DH?�[q��5�L������7������$� $����ٖ���a�{�eR�ٳ���(κjFv�;\J��˸�N	��c�aG�ޝg�7�q�`]�Vy�u����sW��H7Y���V_Ѯ���IVQ3����O��/��ZI���t��\�D�LS�d���(~h�̻i����x#�����Z��l�'k��k��4����N��fN�rS�(��,Ŧ�Ac��7j�2�������$P��	�$�v���NE�]�-:��w,#�ƞi�2З��`�h�w.eeA�GB�����2!Q6��<�c�CE�%ԩ�k��1� ���oD�{g�wg~1�:"x�M��iX"Z7c�k��GQz`<@�0�i�m�?�
��w���O؞7x�
��3��k�e�A��.>�K�=�;sV�vRW��:��� ����5�#��E��8�p�#��Ƅ�\Pa�a�4}������2�z�k�����f��V��1#�6;��=���@�17+���թ��^��:��9:�Ĩo$���CV��7�qh�#�=\��V��,0g�u��ƼTP
�iĭ�P�u �q���|�����=�~��k3�Aﯙ[(�*EDc�i��L�]��O��^��-wI�vl Z��d�ϋ���2R¯֕/�����O���Y/iX-�i���&�8��mQ��ShN\ o�-=��A���s��ʐ5�c�EBk}a�l�4�e*���e!^xF����#UQ��D�I�h�Yq1�e�x��U�h�V�d,�7(?��1� ϔ�,�
W)��T�%�]ݺyw� E���{X��N�g@J�=�4�^��-��โ���A���� �T��E)��:��0�$0[�=�]/׏r��󼱿������6�V���Ϊ&���O�����O��аh��61!�<�&�'��M��ȓs�G	�ulӭ c.cc��Psɱ�f/Y- zL.�F��όd��;<r�eVp�H:À���Q_�i�2��w�딆*{����B�V˗�W#t\��]o7HT����re~��L�KK\}ho�or�F��Cѓ��~B��a�o�"?K]Vr�����(��:�aym��J����Q���AJ<EK�[O�Ȃ���2��[��ա�9����� ��L��ů�S8/'���~��㼛�4�����Z�}���S8���^�d�TP/fȷ�QP����r�h<�7�2{B�$���s◿n�����>뱺�|�_� E��w��QbIɛ����ؐ=
"���Ѭ�y��yE݀���A��4�Fx����{Ij�P���\���2�%j��z�0�P�d^WW� 䕎fo
�C�pҮț�Ͽ��w3,"�@��P�]tO蛫�Aq�V8�sŎf�m���6�N�C�1���Q?�c�`�g��?�������FKYS�^�'����?��������Wi�kGAnB �񳁌���tз��Q}�/���$�b.Z�p1���N\@����p}��/�	������؉��3Xk�E��->{a�������N "�W{0!{|��)���+��ef#�F���Yfy.b$S��=��[� ��zyq���s�X� ��y��k&��N$Q�����`���?�w�X�dq�O���)��&(�BTȑ�]6y��&�9�K��o��6ܻ7�M��9�>�όԹQ�*������ny���Q��O�*�NiY��A�^�d���D��jWW���y��$6�[�"�ò׺m����np���^n�4��*R��2p�&8$���сN�kw�Z�t�}�x4�!�H
;^�H�Z�d{jL��K��v�q|��k����{A���u�߷@���(���ۑ0�@��V:����{f��(��Ҍ�-���:0j���kq}ww�'E��mrઉͶ�g[��K���IT���Fa��.c�~�=q;��bk�jA�����y9�6qU��+��7��ξ��I7�����h��5U�5�+[J>�����J�����1� &�y=���W�¯�`9���rj�m�v�_97�c-�	>2I��t��f�|�!m����AV��)��A�/�ox���X9�x�ȻķV��#�R�ϸc#�tUHQ�P��`�Q��p7�9�Cf���f�^T�q�6W�x7t D����<��/'we���X�)�7÷������,�}�����?�9��R�{FwKV�*D�$�
acA#\9�g��4Edvj�7뀫����ݪb�H����/.�P��1��Ŏ���&jr�g �i{$�0;,Y�$��.��a~�T�ذ�\��UB�b�ʶ'��^:���G�Jn�=���W�Z��qn�2]|�#���~
�ll���N6 �4*?Θ�����{���܆�n�J5zr��)�>�o2��N��  ��f1{��_��o�)Xk��]�;x� ��P��5$�Ox(�4�̡���'<8Nj7:�bX4����0o��pц�'0��.cBu��(z���=�1��V��Y~���ѨT�\����1g����0�
��HlUTk�\��P�Ծ�Ǥ7�s&���e��^�0Ww,
[�7����Þ[�>��=x�ڏ��m�����%	�l�hk��k�����F
d�t�طs\y�9*���.�w7`}O��Y�tð��>zK@b\�Rt�֩)�Kf�׳	��e$<��R��GK=K ��o���a�����xy�)̻��bs�\"n��C���c�آ'ҽ�VT�=���{� C��]�Ŝc\��"NTj]��V@��<�-`>\8��D"�쉼�_!��{b���z��1���k>�}�]��|�⽂3>hh�%xq1Qz#�<Ni��Q"�5��u�Ը���G�Z?����	d�s��,7�hvD�KׁI�C�ȕO��;&�uOYtM 䐋d�^[]oT�x!$��-����m���'�q<�҂Λ�)iH�_N��U����TH���jm& �i��}zx]ܭզ��+q{D��&�r��=��<�\>��Wt��j�ʭ���Ƅg�6�<�X�
��c��#�/_�^�#�$^��x����_���?������N#P(�Σ{��j�1_�ܳ���{�Ө���'cVeXL��'$�w�~݀�_��@a,T'G�[V��&���d\�j@��t�U����¬��S������E=������d�U�s��b�7ΤU��i�}J� _F�ɇ���<�&��E�d��*'1!���碙t�,�ah��#5M��H'�Jwx(6��G�rZ�xY��4�1e�%�r!���ɲ���ij�\�&C���u(²t�c�DMr.�P"��'0�G����������N��iu�>L��-�B.����r7Y�MG�x�A�U���ށ��)y��EW	��IM���{S�:�կ������?"B����4=Wgj{�^d�9�!D�����.��軲�dY���D�{�A��2���ƶ0d �'�X��<��&����Öϯ/���1'O�E�oY�����@oլ`��v�3�����۵^Ĥ�l�*����L��'���<o�˱��m.4 ��ύ���=�5���$�z�=M�^џ�Y��O.���Y����sÄ~_^s��RDd��v�������Z��
�����+qUڨ7�نp5�xz�'������女%t5ͯo�6�
3+�	�T*�Z��twY���in������0tN��O�1��w(!�p�v�'Ǚ��G�*��1��0c�.4��U74���寤�Ӿ��F������� ౔z�,�1�M�+o%���d��,YŢ|��,�OQPXp�����1DVRr��b�H7iy=NAm���u�y|(4�������d�ʾPo�=��Y&�'��K�@V�i��97�lm�=�f2hK2�5��5,{uW�FH^g`�>	�[,	�G��M�G�� l�޳\Y~o9�W�u���]W܍��ƹ�FCn�f�lJ���;L$���;(n�G�B�XW|����t]�r�$&��Z�M��?���/��)�����?S�{q/E�����bQj&��-�:����~w�A; �G�� 7��"?���&֒`�)�{���^�p��S��R|����Ug�ո~*(��[�X� �c��	��7�Iag�g7�	�"�ٝ��� $�M��� �4bd)j��Y��4�8w�����Б��ų���Oq�D����Z_�+x��6��A����\?zV ����0�ѓfl���E	>i���jۚ��#��uB��9k�
yxj"�;�,	� �X�b�A>�o{��g} Z���l������c�C �X�e��� 4>3��7����U$��Z�,BӪv�I��-���E��&F���|��o��7w0��<G��t1�i���v��b:a�`f���=3��f�pn�7k<Ս���C�1c�Ȕ.�A��ɇ7��#.�7������O�8޹S����MS�*ɕƱJd��4x��)��m�r ���������y4A2^� S��|<� ��
P�����?��HB�E'6l�`)���w��h��г�k/TVq�t�KO���rv��*�[ȯ��xP���>nH�E���FV_�������������M�Fp��X�J�R��*�u��]�����N"r-t(%�gc�j �#�25J��^���(~ӗs�G��W˕U��E͢Pm��:y��j�I:�ʮrv�j�rE�9;Re�N�,Ί*P��ua8-k��(c�17�듏��їk�i�=�S�ђ���U��/����,��3����4�/)I���c}�8�}x�%�NA��ƒL��*�7�]9��b^��%��i$|����>�~�Ėa�����N�$���b���r7Q.M�������P��k �P}��:�.��rF*3 ����A�LF��B��:�P~ϗU* 7��M���Vs�}�ȓ��S��1gl�
g�#���C��1�5�c>�S 0�l�Y�=l�����	su*9�.3�E���E�_����ي\�����*5R�bi-�Qwnv��6#y��yh@�.�9�ʭ2g�`��o��7?c8���;=�ǿf7m�-w-������(j�u��X�Y	fڰ��P�:��� HL��+&��r��_2x�D���4�G��D��H��=؆�hq�t�1ާ�{=
�:��v�c��&\ �[D�Af�8A����,���p��` �Y2F��q`��h�������]�t�����Q�	;$��ȍ�kE���,
D���������˽xhDK�e��:/?h�2a<ms���f�� 9�p4����HT��˕��=�+w�u=�ܞ�	��rCkzq41��\zS��q�@Hѝ��
�����Ao��6�MQ��`V
<h��>�5x~�*2ʊ�=���c����-�Ѹ g<ŏ@��A�K��/���{�y�w�A+؃J�<��;���
 �r����|瞜���Љ<|,[1��6z��}t��>C5��y/{�ɫ�>WQ��'�n�s���K��҉cYS�x�&�a�(�&���:JT˅hw�w����6D�_��:/�~.����]?)�B��n!�s.�eD��y>0�z�0g4O��Ö=Zti�[��d�iPP����c�{�=�/[뺯Kjw�$���/J�ixa���0Q�{�E4�_B�3�!�_�WK0��5҂��CL�I�M���I(i�+�
�ܜ���}��D4���_���T��1ٟk)��D��O�d�pR뭩#*Q��cd����,H�'�w���l>f���7��J�[�(A�F��V|}'��J( �Pv�6�?t܇i1$��W�|������: ��wH"���N_ȊeB�����M4/l�T�]���nĴ:�*l�!��0�%���7��&�j$�|��>XN�;Ɨ�m5B�6��~z���[5��q���'��Gݎ]-�I'��ӭ�������f�3���׻c�^�����j9�Km����v�-1�5I�YCE-�}i#����Лpspws��'�f��*r8�A����CEҿ�(QQ0��*��)��
����IxL�Y�%�+k�~aK�4z����p�����|㑎��}Á�W�dnN:���A�u��Gµ��i�Yj�s�f�s��By�Σ���ٽ�%s� ����ѫ�n�|��$ξ��ߧ6ͅ���^C��E�|�>eG	[b�"��*Tb�qn�֥�c��O糮yB������x]���0:�,�H�᪔O���i����/ĭ�6����c��z����pʀ5��5$�}��5��"u��N˖�5��r��o�����1],�~��fO�U8˛��X�al��󥖾�'!��(�"�x9�f��,�Ӄ/ �;׉ĵ
l��EZ�Nפ��)�U^b>�̒CTլ�8�6#�SP�&�v�� �u5on���q'��3��Vf{��H�M�]'��__���@������9��Ƴ��43L�D��9Oy�I�S4��Y���0�[���u!�8�e��߁�tE��n���nf)c�y��?���T�0&ϟi��:��`c(� g� �*�B�+!5�u�_���u0��p�[�����o1��ݨc�}{7a˩�\�1{��X�k�@O6��QR;/v=EhVTt�M�U�=�&�iObV����
���V��S�(3�0����&e	mR�+�|x������I�e�Xr���S��(Q2w/䤻�n�tɬ�yq]-ha&)��(S�6,-��"������p�Mʅlu�2��dx�L$f/�jz�w&��P��nAbĜ4U~�f�Y��Z�x��S������ϝ=��J�u���$���Q��]ϐ?#�&�\����qK[h�/�m-�7Ƭ�4n��)5���*�PF�/_��t��_v��ܒ[h��ݧ��e@��^��i~���ڕ�\.׺%~�GiWH����/��0��K���,3zHc�O-Ca�&}���;�ע��J�Lb�]��G=IO�8F�}e�_��wTə��s\�`���Q������̮4���ngQjQq���I�� ���ț��'V��f�J�(�r,,�=H+��)T�(U	�>�yc������8�"Z*K�_^.�*s@�?v���)#�C��h����~�\��v:ߪg�B<��d�vK �1�ƪڬ�T4
�M���9�o)т`�T7ԕA�hxt��~g�}0��޵ׄ�0y� �M#6o
;���t��&�\%�5�Kٳ��˟1��4����8�+���g1繩Mn��.��E��720�J2�'i��d���%�m3�Fd¾��=2��|���i�P#��ϧ�
�}���T%�Jg��W�9��?bASv#��m&��l秴�o4�x/j��άgٞZ_o�!T�h�d2+���3����N����cncO� dd�;�5h9�q�j������\b����e�NhQ�}��v��7.��l�6R�O��ן�w����YA��:�3�=װ��=EF9�_/ (>��^�oM[�^st�Z������jYᬜz���|���OuA��$bG�Rf�D�	*E�n��N'rK��@]Z����R�￿�)ArN��@���R}���(L�!�v��zޒ���A2RO�l+��_4T����Ι4{�޸�郳����B�2`��5�Υk����4�F��C�6v���t�#}��^ ]nI��o�w+ơ���ts�Ah8�=9��pD�n"yp��y�����ָ��ʚq9s�I������S��j<Ϫ|��m!�W����P'2�j�I�!s!sΔ���ϙ��-U��S#�-d����%҆dm��P�#�A_���:掳T�дL�'9����ʹ�$����+ك���n���Z���Ο��?iK����oP"y�B��{�w䀡�Ըm�֍���n�U�'�$�~'+���0�Ꭴ��3��;Ld���̸E�s{/O�9ퟷ�Mu�!�$#�iVߠa���-�ൢ��3!=��rѭK��הYCI��B�KEb�W飘#�RJ�l3+U6����p�:.��e$��T�>���Q��=C�
YS2����Y9r�G*U�X3�0�gr�5��D����^����Q8�4*��^uo�ZL����S&��i�7��1AD�B����#����E��c[bކ;�3f<�ԇ3�I��^ �����,����N�2�ݑa��ݒ�φ�J·��u,\4�%A1ۭa��ܓ�4F���c})�O�3����Ⓧ{�0F��w��q���"�AB*��O:�h��Z�b��6�JK ��Wt����o�����2_�����(tN��G�b*��3�G?łρ�/MJ�a��\'o�M��ԗ�?����{���3
���3w�t��E,7�'����S�b���?�vD��b��Pu�u�,s��ݛo��evB�G����II���6e�LCS�x@#����L���bB�Ks��uw(Bo���eȽ���k(�Eo�%�M��άb��v8�PfXy<��rOc�2����F ���؏�=����缵��U9�~���֚�� ��i���JP7^tXB#N/�^��������jQNu�pW��7�l�)9�<u��g��-p��ɒԇ�v��C�'���k��AՆ�k��2���,waMf��(�m$�����2l�S�z�p�,�ժ�sr^HG%�,�_��p��%\=h2n��z������:Du�w�g�3i�%��!pԐG�mC+x��JW���1M����^��͏y⧩�P&�lH���61�o5������"�䐽��I�;\u���Y%@�}�L^x�Cٍ�����P�D�}���A�����K���vݯg���u������zғ9+0�A"�M�p�Yՠ
�\9�xUBzT?��	h��{k)�-��o�m�o��Θ�Zŭ�<	��[�7��U�iN��Gb�w���p�3�x�j=��vB��G�bY�4n���}#�2�G��w�L�
�ry]�nw�Aq`if(��� K�T��>����c5��C%�ymόg��z�郩`��¶6Qt)��f?3[J��kq�Gc6���A�)#���q��6��XJ�� 7�IN䶗�),��AÛ�U��#�P�[�"X܇B"m���4]a	X	�t\�g�m*g�/�#���B����9KcJ�#�B8���t7ʛ��G��>�)�(x�����R�Gxz��F�4��Ϩ[K�x���w�Z�����`����3��;�G�� U�^+<�.rzȸ݂;$oWS�pԹ��m̃�1���B@�il�F�ߚv{#Wť�}E�B0�v��!ք7;m��z���;�"Iș18ҟ�P�=O_�}e:W쿄Jxk㲊U���H���n�N�{��Xm���Ļ]�T��,
�`7Ǌ���:U��H��%FFm瑖���#u��_~V (����3!n
ÈK֒}��9&р�����N�sy��N��a�ڧxw!��VL�/�<����(���=���a���#נ�`� �'XA��w���.Q������5m ���-�a�B2 ���zS����e}�B���
�dEm� "�����#�usr���A{��Y(����kO�
��{��]�X1�.���~7;���w���]ɖ�ZU?��ýe��)u�l�c����ԯ�p�~O;�HX��9&��=��zf0�{�@���Ύs�~�(���x��Dz}ߙ�捉�M�ASڪ2h��h(mv�w[\�S*���-=r۲sRp�'x��ؗ�S�E��qJU�"ۆ�P�����ļ�=���''������Ekp.�6[�&eI��7T��֋�\)�@_%<�F}�Kʺt�}[&�v�n3e�x���M��)̱��u:����J[���c�2�Վ`�_�ļ(z=�{��RH�|�u_��2U5�A B36A�}�蘶��g����T��W�WUX�C�v�/�=y�D%�#�%��xà���0�*xu?Ǘʈ,�M�f����hEh��eD����$�зu	�k�!Y�0G��s��&10�zg���LqAr7���*�^�;Z��
��!��F��x�=dQ���)~���>#r�|j��r�bY�`f(�z`�f��\UZ�b�K"����}_��xw����o��%�Q
sA~K�&��`�6#k�,�����M��.7�y�ϸYM'������!���ĮH��@�M��1� �@�5�_�:k[p_�@!��Jt�-���O��J�s=�6g�[�[��g( �~��B㞯ߝ�p��d����'�<�4���EdQ
d�u�����T���a+�υ�煌���?��$U�`$k�6�c�@\� �ـ���Р�.������"�tX�)g��' �cU
�ª��Fy\u����.[�h�<����!=6��%`qlK�9O�h�pJ&V�j� `j#P=ϜЉBb_F�8�w��zǢ�_X�}x$�]�cz��R�,zn�����kla2��_`}&Q�&���+�ˎ�?amU�;��L���ÿ,#�D�$̞/�s�/��ʛ���'��HX��2�T��g��Ő���ו��l�(�!� �����;�c�]ϖ�Y+�V5N��w4@y.�Jn����;����\��8xHX���b\;���d4��n1�)�����=	��gyNN)acM�N��Xô|�D����8{�O��e���A��D,x���*G�L:�|��&\��
�#�}Z����ṷ�fl�j�oK#á9Wm��
��s��k*�?��15�� ��Bs85�����"��lԱ�zȨ�E���kMh3��ݟ�Օϳ��Km��{ڕ~�J^ev�������q��2��r��|(�1���Y�gF_�e��Z��pYɔi<9���ő(�~������x�ܯ�
 kD3Ȋ+^7A#u�]�M#��8�N�@�;8�]�������TK,=�}9JMڔg�p�(��-5��D��ʊ��w��d�ӭ����_�Q$�V�؀���\h@x��f\�z[e�Ю���J ^��۪�3�Q1�� ��\7a˵���I^+��H��"� ;tq2�H�q,!�6���*AT0�	�j	�j3�^E�u�;���q5�z�A�',|�>�Gl��8���D��ev�ރ8$$m�Iz�MCz>�����P��>h�hik���ƏkKS����.׃1�\�>%n��>"�,�#Z�Niw��1{IQVv:]!��p�n���`
P�����U��U�u����H*>�,\Zx<�X[���*C
��=0t����BB ��	�I[OԲ��{74��/�#Y��5�[t�ƌxe=\���,�y!�Z\��VB���\��pt=�b�I7��敩s�u���t����-	Z�`�|A�Z���P�������uU:����p�@5@�\C���<!P���T��0��-��D�HY�F2	�Z�Z��D%�.\7׸}j�?2��3X���}���0Pfdw���t+M�w􈺵6X�O؜_��.
<il�;ʽ@��O�i�׋�ז��
"vDu�ݶ��o��S�
�6�,�{w[�g&2RI�%��$���{���Y=���U��.J�-+O��@*�N|���������vG��ֵ���4���f̔�>�W��"��)�8p �<+��Y�c�>�o/*d�v��;��r�k�}Ev��l�<!�?��Hf� �_�y|�%��M��s�0\����6��}9��M��攍�Y�@#W�:�kSAi�|"*#�Np�+i+����WǶp.�F�:w�\��z��i]�Q��}�	��p�em_$�i��P�=W
ң�i�}\�������@���w�k��e�R_�����!��U����u�ى$	<�Fw�"�l�Y���"X��R�q����#�L)�ڟ)�@j�9��-��gcV�Nz%8@Da�9���, o�o�n������3��-�V_G$u�QV�v��2���c��o�b
.(���o��/��ٳ��Y5�mrOSb�v��U��;�hލ�a��zF������ڈk@~��X���V<5D��^Oi���p����9�N�B��Y@l�+*��]2�R�3z�{�Ѡ�ɷ�K]��PK��w,�4(�J#Y3o��Kk;�[���VP��uGS�6~���+.#�f/A���!�@lZ���~ �"4��s�mn���1��KЙY�e:�̻�g�o�!)�$��ve�.�n%����������p����n�g�\���,�I��+�x}[QyP���^ao3[@�����Д��o<p�t�W�tr�����6>��oU�vP���;�P�ei�	��^4z�n�"![����$�	J��)d�`��EeN�~���`h�@�u?DZ������Q镋�Nd��i>D}����i�w����%��~�
�|HA�J1�uR$'�,0��f�M������u,��x�I�����D�;.Q�_��굌p�X�$j�\�|]r��x���M�8Y���$ǔ	�P��J�1>��Ů�%
})�긌Q�v��F�E��?�3��C����6��!o1 �M�e8;>� �}Y}Z�Y�C����|C��e����&�`����D�`�$�?�(m�c��$2ݫ"J���d��
��㲊���C��~����%R�I)�~��|Q㈛R���.Bw*������M��f��T�s�Z���V����v+Aǣ�E��F��!����*�=nK4�������9c�Z���+#��և�<)G
g��H\*#�I�ZJ@W#�����f���^���/���I�M��i|j�^��&�
�>r��t���-�5��o�XNs�)�ި7MG\cd�ƿ/�G��E3�g���?���G�0��S�V<T�����4��zȢ(���q��A?�l	9
�Z�g��`�6o�C���\�2<$EC#��w�X�*��Yt�$,<�����;��>&!�M��t�e=|��L�,߉�UD)������-��|�bK�/����ط�y�ϼWX��ظt�ث��w0� �7Ob���R���:_6�k'D4Aҍ�-u��R�����TVl��`����a�3�c�f'�؎�g&$�\mۥ(K��(���:NR�v�j�q�3��!��<"7N�"��	e�n�K:ӱ��2�- ����a#�N���h��l��kh�{�a� xi=7��f����
:r5���]h3�~Nr���"�ٍt��*�2�k$DY�D�K,�`���{�y������(5����r�����l��|�6uwfǉ��뚌[�zL��Sy�$�d:M��g�ӊ��V��}}���˽�����U ��RDϐ���M���U�Ҡ��RY)�?�
x�0�MH*��s��t9o��yO�,]��B���i=�������H���5���3�g�,*�/�L�A�#`�����8���8DR�^J5��>������V����܏`��Zm�3�::z(�?\��o��F���jYu��ƐS�c������,�[�#�x�'������k�3�^�='8�yi4@��5ZZ�X{�ꙍ�={%_�����ݚN�2�AW߼�B�Pa�ӿ���X�c@�!��`u�Q	��j�Ъ�4�}�f��4 �/OFvs�L�P��C��W�E��й,&�i/��=Ѹw��5��f*�A��ڦ�#V�M/�@ƯA��;'����F��J 9��<(����J�/T���$��M]�ٝ�=��i�=c�Ё&u�j�����Ť>��9꼺n�co���"˙2MB���p �5`Ę���?��jC�~e��T��p5#J�s��Y���17�F�7�ɻa��yۨa~���,_%ߠ"�2�`�cZx7%�8���F�~%W����$���s3�ܠb�QsO�����7
����%G�c�3�Ӵ<8J�E�C�/c��1\P{Y{~�rP��l~P�����Ӕ��U��lC�ܭ7�E���ڵ0���N.��UI�d��]ՠt����Hmu I2���ك4��Q��3�����W!�KF��r�݂��E���a���P��/�G�8S��uU���������S�Hgw2U9�6A�G/��&Og�5�[o����
�g�4~tc!�{�ۄI�����w���S�z���Ҍt��M�,kmͶ��R�N�uF��B�^n��[<}mj����5d�41u���-l�#�!h�©��I)�� �d����W2�9����tU�#�>2�8 ��DF��ȕ�fj
 ��h#��^�p�\;�b�S<�2E�k�K\���#�]�F�߃S�!)|�ZJ^�/�;����c !jk5�����DBѠ�*3���c�3�
�_��`��n�����=R�km�֑�����09�j�����Iu'�N.��C��?>��1��I������ ��&t�<��"3a�~������o���k.y�B�o6��ri�M��l��w���i��ɄXk69����[�!�z@�Y	|�
P��KZ�э�3�x[���OΗ���-��Fs\N�=��<�� ;2��A�`�)
�ar!k����`az��y;^���}���0�U���/	��B���ө�\\sy=N�	��O���0��,Z4�U=7�Z��K��E!��wz�{���ǰ�픞䂅cl��c� �$G^G+����7��Ԫe�;n�����02�y���Vh�Z�	���b��/<���س<���_ܝʟ�Mq�j�? �iQS:U�Q���W9�x:�{<)��@��9�a^��'��s��H#�
�w)^��:���'�] ������_����pλXZ^�'�d�}�������iu��f�vu%���G��-��5Бjx����
Z�a~CM�:�`h�>�}�NԿvYh]5}q�p ���_
ݬ�8��c0��'�y+��l���P\&�H�T&��z@�/5�/�T8�fP�8�݉�V�������|�:���Ǜjܚ}f}s���Z�$��%�'�U���B�u��E�?eM�z�!!�+��來�!@ٝ491���#� p$����dN>2]��A?�P��~Xڇ���NN�cf�n�7�t�眾#� ���c�ɦ^�����JQ�@%)��ڶ���T� ar��ȫI}�j�E�	�%�f;�ȅ�X�w��{��>6ے�2=g�W�n�@;Tk��1���*~[�+$LTG�� $��F�qMj6N+Z5;×�rGi�Td=�w\���bX.��#D^Y^��,��3M2G��doM�:��%=���)��׫e��g����R���c�nȒ��F�u@F���LmP����?��QV�jF��a,,���/�(�f��V��Z��- �P�Y�t�P^5�VS'�-�4_�����߼ m�i#�~n+EDd���W(���a9(s�$	?��!��w�B���Ĝ��Rd�e�j�~{�}��ӚX�C�X1F�3釆�;�{�ȩ�R��'R	���'�����u���/֚�R��eX:����d�6ܐ@�r0�R�����M3�[������"i`(Æ*1bCzB"C=൯��(b/yv�f�x6����u�9G�QX�� "�o���M:��J?K��6�~���Q���1�e3:�*�L4�DF��Y��@7����!���W��95�d)�M�jL���;]�ߊO�(���MV�H=��-�y���j����4{"3�������u+���e�|��s�)4�5ꋱ[W�a�{l���=�#�7E={8��+��a',��J�'�r���il��E:�v���l4�K���F\�W.֘b�-p��*e�+F_��{�b���Xʝ�)� �I�jǺ0�x7���u�1��*��bd9Ǭ*b��X�ڒ��NKc0�5����>��R��a,؀6p&���_'(��_���=�a�a+�x�pb�-(��	�NQy�ޓkT�Һ3�@���4\\�K�K=x+]4H����yEϜ��%�����z�,*�4�H����Ź�;�y2��"]���Jf�9%���J�ɓ��է�w���+u�-��;�0�?ߤ8��^m����-!+F�W���)�}=)䲯0��ȋE�\A��ő������z蛔��Pʓ��	��c����<N9��6�ݷ�g�� i�@'�<f��k烟� ؾ3;����Lٽf=Z��z�zKtckj8���6�$
����ʄx���^�z�p�����IZ(W^�6w#�So���N��rƒ���ς*���!G�y'h�`˰F�9;W��nŲ�Vp����r�q&�����g�D#v�g�݁���a�ź���"��Ҫ%>��m
�\��\�����e ^��yk|.MJ�Y��x��w�rn}Xu��m'M_`�uo̍�B�tX���{����
E��? �}��U��h���y�ŉ��C�2�u�Ӛ���7[�9�1%E�	c� P�[E��x�����X�l��TDߦ��P̐L�OSr�C�8�9a��ڠ	*=[B4�̌z?��A�:0ٯ��D\^<�[�ޢ=d�B�` ����R��P��.$�F��l��������(C ��iG��ʅ��/��J���O�>T�@xh`j�L?���؏�L�財H~���C�e�fI�:]��5����'N��BX�&��b|�w-��$rYh_m�������I���wթ��Ĵ:�3��y����zcC�/�y3���� �z�$%���|���m����&�5#�F��d�ck��NJ3۰���\�Q�9������!Bn�b�)�z���D����GB3y�ľ�$�o_L�nĐ����ʹ/wn�5�EJVGxI^���ū�3	̮
&'���s���Q0Y�1�4F]:Q�R�fT��]L����P�Z֙%L�j�j/�'��{X�Dk�����h�jX�
8�D=2�	���x���qpqa!9�xT$]MHy� Gt�??B�O�J���D���k9�@�DM�G�h�����"��u-�O�4���ߥoi�^9W�贋$������m-#�.�8���SJq���<�l���S�2^�in$��!���0^Xh}���Nl�_*���,cA:�d$2�Z�H���_�T����%��y�7xH�	)NMćޭ���!��d߁�=��\��R�	3*���'/�dV�j.>�:�e�tg��[�=*�"��"�r #��,^a+�y ��X��4S��e�|i�`Ͻ�:�^����a��FRA@J?S���Q��  k �c���/�9 ���߀jĤ�E܈�b��9�!��F�{�0zk$�l�Y[�\��l-@
s���ʵ�h�ܝ#}�2ds0�|�2ת���u����l����:�ӅU�f>^)m��k3#
X�;*Յ��j��%�UE~ �8C��k�(��/�]јx���U�ĬL,+�rL_?��-�l���D�Kp�DZ�rְ�=�{S�i��7���n3!Uw�r|���Y�HK]�h�@����+T0T�%d .Iᶗjx��:XWEG~�7=�G�uc�2�X��.1h�`f{j�/��k��
�6��v�m䄌NO�Iؿ���`A��7��oG_����aN1�.-��s4�=�mMx�T��pU!�=�f�D��Ka:�?���y�YjM�$�5��=��?Q�����p�2�9zx��ע;�sqSY;��CK'��z�M�|��
bؚ��y��I06��R�^�7���i�l-#2������ɨ�4�� �L�D�$���h����a^��y�{\� :V��c�8�R�"糹(�����#-t�E�9.��C 5�cj���ڤ��z��p���%�o������Z�J���3��t�� F���hGC�v[�|�ʅ�����@��z
�숭U)�m�L̽@��UdՕ��a̓!¼�ϟ��	�%A�=�*�hgb���������VO0�xJY��t5%���L��,�+u'�)%Sn�#��Z������1�T�;��߽����<�e�|����͗��w%�t��G��&7��ۄq�η�4�c��H���=�;�}z"�K̚�F�p�3z�
��%b=c�պJ�z��]�>�����J*�A�� �Ft��)��d
G˂�t! ��Rm��t;��	�Lx�m�	ƍ8%�˝n�
*9�Ae���j���t�J��aM��,ց�r�Ӆ՞���=Vc9/��4hk���3�,������S�}��j��m���X��:�)8}t�n7���+�0��ܿ��bϹ�r�,�t�i�>�C��O}d)���2��T���(������Oqp�7�D�@�U�o=�����Xm{ϝ���A�ې�jS&t}K-P%78M�aA��{z�y7�O:��}��e&��Â�*�Q��t�6�!!+֏9ǻ�& כ��b��s';�e�.v6|����l�F�J�L4Iv��oz0�����?�3�����J��D"���Í>
OW	�԰�X�o��-��V���қ<,\=��� c���<r���KO-���Y�8E��.��h��b*(���9�-�I>D;P�����Eke�ѝ�y(���}7b�g��j]1K�l=y���H�/y,��My�HK�Ň?��yOu}��FTǭ�E���05���F�S$ܒt��	%#D�[�#���4|��F�z8%��Y��<��O#�W��LD���(Ia`U��ǚ��eOx�b!�`���v�a^�3m��a���Aag^6~���"�x�� �ɛ�Q$�����S����0?2�:z��:�j�_48�]̕.RIn��O$��oŹ�������W�hxA�V<�������]�G١l���J���r���b�d1��[�h��&{�����s��TZ&�_{���iP,H^3᪹��g(N2D� Na�J.,ɡΚb&Fߝ�����W(�>W4�i�f�������!�W���;��>��2`��~.;������n40�%�Md�??��9G��iOm�cu�~D+��e���*��hx'v a�W>�k�B6��i\���`�S�ؐk	1�0���Ɔ��c��.h7PS���-���o��!����T�{X�wkQ��>�����b��A�T��M�D��.mb��%O�<~R�nPC<=~�S��)7&��G����}n
� �Ŕ��.�F��ɒ�i��UTG��k�a����IXIw"]�Al�������|���l��KcinQ�A�~l�p�)��K�
����ƌ
��@/�����������a����<�E;0%�b�pt!�ώґ��m%��p�袶z�\�8�Ђ�)����Ĭ��},��73l��ZG�����V#�B���Tr ����ٽv�.��%�߬x��yV��&e���6�<��P����TX]�Zx�q2�2h�颽i��).GLX�J�SlUt���zy��h~�<�l�4��
�
I�Y�����v�f�����^� H������1Z�4p��SI�JA�9h�]�݁}����1V��\ؾ=�NY�v�}~pT8�v�7w�M���F��k���H�5�'Og���ŏ��6����z$%�,�wDv����t4��>9-\�q��8���S�k�;"D)��������桧v�z�->H��>"�4��|U�&�c����W�:N�4�Q�`� �HPΠ�xpW}��>�PT~�E�Ρ�/jN�H��Y'vL<dJX  c�c���7ny�V		��J�Iڀ֡�g���'7cV��h�U���8��򲂁�I'B�`-2� gq\�(�?���"Ԅ�cu\��Ӛ�QT��N8�j����In����&S��;BmK�{"#����gU��R��2}��o����i�{�[R�-Ҡ��Pli�ED����k&�v+�1�ߪ�ų�5��s�Eݰ�boy�	����GhǮd<��1�	��M�_	#��PX���+g�=����#�y��1��|e J�/x+�!�-�i"$�T�ǜu?�Z%(0.�[#ݟ4��Ǹ���?/>;e�B�1�/^�O���z��ʙ���c�aK�֘�8"�����pPh��%WD7t��)5*a����g�~1�J&����_?C�8�r�����.�����U*q?���v���\u�8������8�Ҝ&�>z�#�̀�b	??�zn��������8&i�V� �34�/Q��S�_ea�u/b+�W���Ѧ���,_�.A\�3�Ш��'I�ھ�SW������3`� ��MY�F���/2+�]�e�[~Bxp��5����h�Ow����׫6������9/P4�<�r�dݚ2�9��r�_c��%�gb�p��`ߖ_�_u�'����&9'35���	��<YL��ݘԧrw�x����ob��ƈ	a�4N��y��^3O��2chz(�~.a���-P:ě�6�?k���m���ގ`ϩ��u������>��*�]$��z�T�i^�-~I.�JO.�G�Q&yW�,���R03��E�2���E�z��F�#sX�s��R����vU�I6�����9���Ф�nO��ʸ��:m�|�>��o�}HwR��6�����"��&�_��Q&�eN�}��_]�	��+xs�Ǵ�S�1Z#�(��S�7;��	1��!�b� U^����ƴ�b?,�&K�m��Gd>Cw5!U-�k�6Ï�TO��*��v�Ȳg~�7�.�;��٧Not�������:�Od����l
ґF���pN?kk��������|/L������&.$/0���7��^�{������V<T!����q���xgt!׎x��*]��-jpX\:5����Mp�����_�M{��Br��1���RF
u��.����tM5�%��5�x�̺��UbY���#��
��EE�J���f���t ��A�pi-���UX�u��e ͌o�$/�3�=>H�T��3#��88o������-Z�!�<�.�<����݋��
o5x��I�3�y�>o�q8-.�_>��� ��ȃY麵�)`����U��<�~~h�����a�)}C�F�*ՙ. �l���ܮ[/�j�N�s���mw�-UdL;؇���z���<���{��_bg���:�[e�S����ހ�47�7g�7�YF�3����T4��߃y-J�m���š����>���p��>�	8֌\��=^s�
�O�č\��U��Q}���5���O�2�1D��JLP�.��J]����;����/B�l�S	f���X� '\l!�H������o_��it8�+,�A�z-P�ix�v�Ŕ`�a̰���
g$8o}������8�ts�.@��SB�O�i�klE<�`H���~�$)�������H���D!�5>�'����^����^��p���^���D-�Wa����2�E�K6���K���q%�BȰnP��˒��˺�9cD�#rt�.�}!�Aa��������!�#��~[}g��#o�_0$̀�Av�ij�ۇ��>��j\A�h5�X��:?�i�Cg��ʴ�Yz^����X���&z�Dߵ�u��sP61H�3ϫ�s�0'�O�t�,b��ft���#3��C��`�ntX%����h���Du����0v�(�;p�bw�i�d�$�w��^�	�c+IWc��\�k(�	��SăB��
���]�LO�-鹵W�-������f����h���-p@�ؘ�� �:b��s��0?�v0�� iP��-�қ��r��Q���*��\��Ly�LдY"��xzj?3[(�0T9�����Ri� ��E!y�QI?��I.	t�Y���M����GJ���$����T*�ގ�=���w���cu�!����ɎOlKg���~|�z� �ĂΐY�2Ъ���u��%�d^�v
N��N0Ŏ��������p='��=��U��5�!vJ90y��T˅�49�.s�ۇ��=N��4XZ*'$c})6�s� ���fꎰS�ds�mc�S�s-),?�J
5��ܗc�	�ϔ<T������0�s3�"g��9ൃ�����Q�^az��<�<\;�%�����{wRy�+(@Xa��|����=剺���vO�E�5B2�iW-����@Xw*��3�O�6g�ݎ��æLww�xQK��?�W�#�@5AU�����F�0��b�4��&f��5�7���Z�#�+��p&��+�yy�����?"��}4Z.�Ŀ	��-��տ�#���a�pxN�%>�=|���G"�Gd�b�$	(7d��S4d���/��݅�}����9L&�������#�%�e����=	� ��E(�,����*�g=/�:�wJ�97��叩�U�
T��Sv�!�#��S��@}����j����n��2Vn_(�ʽ8�&��2ԐN	��"�H'#GxC�J���J3����l������:>��fP�Id�`�ױ 9�oS�j��_�>*��COn�0ظ�._'�f�*�$�l;��!�}��j�����bM>Τ�[I0O��IW����ZT,��*-�JL*g������?D�@�=��_����\�%�A�-C��{�E;�Ɠ��b��3>�w�YWĶ�9�7"�zf����ۉ�!5�֌cK�o�A��a���>gr�%���4>��hqP-�;�`�C�d,o����*-�^����	w]�)��p���:t�\�.��Oq>���;J�^�4�N�������J����jKaIq��	��Y}%n򽧷n���æ؋
^������E�c�l��s��=3��������Jhǥ���.�i�.҃�q��RUmd1(���*K⒠�?U`��1'R�!�O'#�/W�jc!��S˝��,N:���5��j�"�K��n�L]@���W�K"�5����t_�f5`���30�\�Ĳ1��䔻#fn`�dF�$.�y���x���`Ɵ.e�x,+��|��[���D�k�����}̎S`�)"���y��%P�(Ĳ�|{�_�9�G"�D�x��xW�(�Y�2P�l��\v������k�����j'�U�ѻ��ͧ���roT'�.vc�-��{¬7�,*:�Yӌ&�V���duZ�W�$kEF�ԌP�e]^C����p.�Q��4�~��OW�̜gki����Sl���M?\�}��2 o_�Z�v!��`��uL��	�[�ˠ�}�^��5�M?�T��w�0@�M#��O��f��z\ �j��2\(�g�k�>��`�x��l4/��3I �\��p�Mlee�
#ks�^��s?�T�����,��2`������o��:�҄��X�R����1I�T(>���6wE��"BpST�k��Ny�ʘ[�`�~��gH�f���eΔ�\m��/����=��`�����J�j5���V~�(�F� _焎�ϔU�Zf�U���&L�}��q*���&���0T�L� N��	�W}#[���&rY�2�Vo��BZ�:,X�B0�pV������S~��B���p��Y�alU@������pD�wά-�5��k�R�F��a��F�H]`ʯ���)pSEW�Y�-�F�#d6 y~�?R6�K 9FF�G����!.�O�m-�ɠ�ތҴ�v�u�����K/�d�Y�4uZ]����Yt�];��ד6�?��k�w0��d���m��^�C)��m����ؓ�f�� fc�y��"
�̈́����m���_fnvm�uޔ��~�*�L����8��	�r#"&#�,Lo>�g�gM�@��-|��b�W9�-�����{�s��?6���`v����#l��g���S~1��U��a�l&�P0�td�%���K7q]�i�r\�/�S�L9�>E��Bt7lP�n����B^��7�\�����2�P�QQ\���ቹC���.c=Gp��3�`c�QX�	��u�	�4Kk���Ey�7���2�%I�4~ �F�S�pT��19���z�W2/�_W:��z�e�"�Ȥ �d�Jr��<�j&�53^�^�����qΙ��S�>x�z�Sd]M���X~T�J�G?��#J$ �"IF�c<���'!ps��D�P���z��؝�⚑D	�C�F�����eY,�sn��9�f�-�@_<��% � �dLAjB��������-I?�w�(#pD����yp
DF0�޴�l�l����.��c7�2��}Y�J�-��՜�:��9�N�+�K*92�^O��$��ݍ����=�&��Qf�v^�mU;P\�J���MGD�8�.j�=hT�]"�F��
d��d��<�*4�&G0�W!�AQ�ɽs�mr��h�5�d�$��l�M��m�˝r�
�s�L��P��E����� ��h_>O����%��:��I�m�A=�і�GH�EzB
��#h"��o���pU�Ho���>=��u��.Q�����ݳ=���a(&����uɮ����0[4��������;V�F�0稄aHI'c�G��ϙ݈+G;1����5�E��}#�Ső|��10��L,"�b4$��zTv����YB5>��a���( ?2�U���yQmx�ߢy|�-{��;�Au��9Ul��w��u����f���z"���J�, �����tݪ��M>Һ/�p��c���U�����r�ĉ皴�腨HO;����ba
�bf³T��Qu"��4�J�f�N�qn�(���@�5y�7P��I�����
���X��IH}��10�b���3�� �Ӽ���k�G����?��
�yLw��R�5[^�:�YC0U����ć�HI�h�l&�S`��j	�&V2"L�#bx;�����W�fy�o<L�`<��i�]���"j�b#mdAl^���P�O�u����� ��å�W@ݩ4��D��	���R�L��a
�1ݶ��<��=.�$wESh�$3�#�et}��A��b�@qª�^������`!�"]%������EY7����w�3�QcE�O�:q�I*�� s�����_�2%HCy�]h����1u����[/�XD�B B7���fr[u�DQX��0Nw�\B@�l�-�hN2i1"�)�`�m�Eb*�գ���~�,*�����M�$5l����jvO�ћU���=��!��R���� [��:��\�;��5y\�,r꧊_(��F�Ѯ,֬Aؠ}0�]
��&j]:��{�豶��K���Ir�>��l��$ ��j���·�V�3��%,�m����t&����E��^�AJ�+������"*n��!�%�Y�{��I+�ig?hs�s,+�y�gypV��y��|���t�ᡆ�Br_�Zo����|`4l�r~e�V����{�6-u�\��E�X�{��z��u�$���#�ק'b@Q�Fh!��~��z�cE��>�W[+�>��i`���N`�QHT| �O��:r=�y�M�Ǧ���s(��xcI�7(��<�v���pdr+Cf���[����B��7l:Ei'e-Wm�a��t�7�����z�RLB�:p��j`E�6i
���O��$�+3�I[*!�*�I����>�bH�w��I���'^��eFEn��#(�lp�5a��Sw�G�L�4_��U�d@-`��уi���j��R8L��	رl �?�咽�a�u����v�z�`��I�~��d��� �JlQ����f/U`��R+MktK�;�������b�3}��4h�����C$�T�����9�nIئ��HJ��o}�� e�D� �9V�\�@X��Dn��Һ>��$�mjx�_^��`t
�����c��q_�.��j�Aa����,��o=d_ds��aKF�L�ٟj���<����ു��Lț��~�8遶��������Oa<y>Y���M�q����9����k���X� �~���F���*�aW�]��D�}Ew��<4r녮��L&���4h��ȍS��,$��� �!D7�y�6��6S�cH|�3O!I�6=Bt&�]�TR&T�"Z��7��\E�����_i�߰x�"m�f�G��p�|�km`]YiUn	ZW�]ބ�����%7l�x99ҬɈ2�d0��T�>Jh�/��w��_��H7�_ΖCB���i�b(�j,~2��.����ul���}%���=���+�9X�e�sn�M����L��>�����*���,��c�5T�L٬�7��B}(�u���xZQO|��I&I[L�'
��ѳ9�+N^B�=�
}�h�\�V� ��	���vd���:eg�����q�Wx��q+�`��%f�X�vFZO��!���?g�E,r-4�w�c�$[j֝�H�/^W�OP����w�V��ssa0�`���ג�/���h�֮!>ݓS�>/�'8�����L�I�1'�C��T����2��Į.�F���g���Z��?���eȅ;��Gx�=�)j>_��`�R�d��څWI���@�E�
�GT]6�jY4���P�.梢<Ǩ�?y[=Cp�>�x@F'��zTg=�#�py������J0i�٩��O���\�5�
�J����:��ˣϞ�.,v�q'�i�R(���,�������p�4-���"6���mL��"��	_B/b��ͭ'��p-;��<��^)y	6��ga�97�Rh�1��&�L�Gt�O�����E�{��H+eW]��y����sМ��\Ǩ�X	��A��3��t���~J���������J��1�o���;�*��i�GٿS+�m�J'3�XY������_��*�t����U o����>'�����4��|�;��:.@�9~��^��h�����`���Fߋ��
�w<K*P���]�.��r��j�1�1��+�W`�ǃ��C0��E&��-�O藣�ڠ@�{;CĂ��#3r��&���*�@af��#����l��l%�Aw/Ġ`'���U�}9���
��͏�OUP��.��G�m��w���{E��	_����_�UȎey���d��Ns�c�'m˛ɼ�m��B��F���d6�����0.˔�����A��\K���^���b)N܂�Ht	$%u61�ս[ä �SG
"W}�Tp�P#��w1G_��K"��{�`*	����kSq2"y��R`�z6xd2���ޯ�b�sB�)�����N8P@*@�7",Ptm���rC>��ZS�C�m�8y���z���i������F�H�j��W*��yr���-�q�Y�`A	���{[G��3�����D�@�SҒ�o��E�5d��[��$y��q�E6!ݹ��� .�����]����3�г�!�4w�����8�!���{]L��6wѪ�HxQ���I���Fӱ@��}��mR_a&uH��l�Z~[�i��/de��'�>�SX��@����_�����h�	y��y�8)�(�MGR��qe^yT�{Eī����Pȶ�'B��u�8z�C]�{m����W/��� MT:K<��@��|a�*i�� A~!z�y�h�-�^��p8�#"'�k�vnyy�1'3]�N���n�}0���ҧ�}�^�=T&Y8>玬���g7�(D�Ha�G5���I{(9���xܭ�ӍM�;�b;�廪��U�����f3��N�+g�'o�ӈ��:�
�V�6LM����2k�$�S�8���Bk�`/�Tb���1�F|9ג�ZЌW[��)��VZ��&�vhz��bEȼ:C��SL;�75h�՝��dFQ�5`���򋵵��[Wͥn͕���/��9��P�0��L�a��5A�����~���KE}�Y�����`���9����u��|u�qd�X�%�Vs���5r&�w�}��[3�螆�6#��(a��zj2��4 $��|��>\��c��}C��$�5F�K'�3�]��h��:��պ��F�PU�/�$�˩��=cB\���{M`���I�gw�4٦�d6� �Fz�CW��O�����.KT���5st���*�qJ��<�Ax��d������7�1��̙�"�.�КD� ?\�HB�4�Bo�jG��@<xn�͜ŵ�:��v�܉���E���rgبN��{�!��C�k�$5�B9T+�p6+�ױ#[�	�l�v��!����2z�?I�l�y��Jf�c$�.�����`!���S��|{)����P����o���;��z���N̊�8��;rwcV^�
�l��Ȟ���y��|���4��\vv��:�����"���mj�`%�s�rOSV�~��������o�h(��:"�]��3l��f�+�f��&��̙ٓw�udJ�`o2*����r�=%�n�m����d�T/�U����6	�����o#j1� ]�e�R�<���݁`n�ʍ]�G'l�H�AE����S�N�M`���Ҡ��'���t���xA�>�G1E����3��l�N�2O��X41 �E'����a�3�a���X̎6Yu��ٞ�f�����]�r���:`A{hͤ-�9\�@����H��0�����J�YҰ���+�d�3�k<|�8*� �yJ�2�&v�Jlio��	�(8�&$�0~��Q�5��驺�&��N@,��ޟ�cB�e�{j�׏��"�hX�9!���Gb�O�0�wߪ��XK�DHYS�@��Gx�%�F�r�]��wRx�{"����U���<R�d���%�Xי"�H-�o1ω���{��]F�嘠���>�'�;�]3�u�.v � ӕ!S]�%-��W�ؿ�u�:>Q�a�����x��b����!�$�4�a��5 ��c�VK��!�]�|���B�{��]8�p-�2`�
�08�jD�mܱK�A�A�G�� ��k���c%2���-6
LC�Z+{{1�D��M>RoLE�������A;k��_G��	f�����B2��1�3�a���4/7s�OR^sG~Hɥcg&�	��� A�b!GF���c]B��jO��z����h����#O!|/�d1���L��#,0��tm`m��Ng�g����a��繱vD�>�Q�.S�gϒi������U�����U�J# �[�	tЮ���:vv�=����[*!��qO~��T@����cĆ��{*.	Rk�`Ba<���D@��#����*A#��m�d樣�۾�'O���4�N�����	0�8�#�-kS[�#Nk~�(l�8��J��u�_~��\@r�k��x�Ũ�c}�/����ؚ�5�.�������d�r�@,�䨃�3��Q)\x��v k%}�������q�%�������*�]"fB��/���=U��)�i�B$g�93���l���0#��1c�aѼ����v���"�b)D.3�od_G�y��L_�]�;j���	���v����ׅX3N�����G� ��G-t�.o���]a_���`�9��J\'`L�{���i˺�������#rL�}��S/�p9Q�@�JI� ��2�<�@g�!�:n 
^j�WW���:v9�g�@�x�2��ܾ���x��B�����=_H�k,�~3�I�ߠ�#��xS+�+k�8�a�����Y�^	�!D�r3IC�	]�U�Ll��ffJp-�ٷ!�\\�鑵$��p$��c ���vaa>�=�A�xxݻ޲�oq�C��?q����)Cx%w�1h�X����p 2E����w=����
�1�M;�c���q޲Ti�������ǃ���}���ZS��%ۖL	/)�[X�D�'ARC��d3b\ԉC��v˩��k\a�,�T�s���M�$ �c��\I,9��2��aOd�C���:*i�r*^�F�V����`7��tօ3�S��̼K7Tj9��;�b�-"����?�)��UeD�"ۮĀܭ� �6m��ӊM��˫c���{ Z����2�KS��dk���X>>����n��
�W���IpK�$�E;׍
~ί����c'�
��J�����\F3n�J�B}T��+�1��4H��.�`���'�mJ(e���u��T��=l�L+}��!5�A~zS�c^��o�'��A��g들`�ѱ�����؁i�_{�� �x�����7����s?�hm_9�1��\��������G5�H	o_ϊ�W�I�f۴�?�scڔ�����ʺ�b�Ɖ�X^��*h>��lH�d���[+�ڴ�K.�.j�{��_�/� >Xܝ[�ҫL�/��ئ���KtS��g�b{1n1K0�������D���������w{\�s�*�����{y�?5�!=F�)��2X���Q@���7��i�d�G��Į��72������#&9 ���p����$2�=r��~�+��M*$�IG��x-����F�P=l��aR���	�O�7��sC̾QħC@�?,Y,���(3X=�@�A�{�~�[���	>����wp�;\#��$M�S�3w�k	��`Ʊ�w�>���T���)h��y�+��0���2{���e�G]���&�ZI�e4� ��@�,ţ����J$�.mY����)v���W9%@ byez����%�FWE<#��-m��2��Rݮ8��蘋|�����&^�y���{7m~[�)lH�$�zU�~����mJF�}f^є$�����؜��n��3����=��&2K��~��oi5�+���P?e.F��L[ٵ��<��i����b�|��=�@J%������|���;CLw��7�I������QcsW�,f��x�����a�^5�<,Īrd��4���=��<�m�~�W�A�j7��8n?M;1��rfiZ�.�2+��Q��z74��~$�S]�Ŋ�~�``N*��*U�u~���d�
��nn(:�:Xh��w��%��'��u7V���֊�N�3�����}��k_���+Z*����>��
�����R�Fn/'X@v K�i�۪m���Ō1c�t��S�d��6� �Ql�W\7�.�C�j˼(�B�������P��1:�N}հF��{t���R�Zo��.H��_�#��Iw�}�4b���N3�I^������87i�p~f���M�"���Q��]#\j����$�E�(���P� ��{�����{�X�9�������?Iȅ�)�4��+�à�uHOc�+�T�@(�������O7��ArZ����i�Ｃ��vofx/�i�6�X}Q�Ӯ6�S��٧�	Jy*�r$�q^�V0�+�0��ڐox޿\�.6�ɛm+��zU�C J��ZL���+݌��4�+q��U
1��~@���V��)����?��
�=�����L�;��]�����D1��n��(��6ѩdi���Ż%��`��Y�H��xn��%}�=��yh)������,�#�~^__[��ann�A�hl�Ț�X���8�V?�z�D_�WY�u�,ռ)����u�I��w²�=!i7HW�"h���zﴯ�]*�*��̉��}��խ�``f���O�{�H���4K����\3��E݄f
�j�L�C�D�����~�Y�R��<�9����f���,C&��^��x3��B�:L�*��f?}��f�/�%�
�9Wϛxߟ����-\�-dx�;Icʮgy/&ۡV������й{�r��E��T�
�^�޸H���p�If)F*vS�;آ�xF�e����#�����*��̴����J��w����_������G��!�Qx�$ج'[����!u�s۠u�H�!�P z�Y��ݱju�6ҍ�	�\�/0z�N�28<ⅆ筟BG����]���꧖��a�Jz����Zn�i9FU`�䩓�*�y@��|��Np�Į��X}B�u6*b!�Q|�
׭+��Z�s�,o'��aG�����8�0��,d��x�ϥ�	�N|��M��@?���	3	�+�BKV��i���l����ܦ��>�N�b)<<�g��o�x���� ��R�Q�|�#�"���=���o�u�����l��Ti<2�Br�� 8 ��W��o����ݴ���ہ��1{��!����S�@�2���p��'�0o� ��xoEf���8��Q0���<_���F'�o�G�,b]4:��M$��{�^c�U���Ukܕ�\$�W+��]���O�u=/M�!rT��b$�D�:fZ�\8�F�Pc�ɰ�i�k�
��Xb�m<��N�֍Y��y���' 2]�6�$����Q�6�a2�t�7�6�O"nK���?�˭���hX��mwb/�2��s���뺵�*.�}v�)�!J�����#�롈�ZT�������+ŝ�9�^Ũ�jry���m$hɖ�N�����g�J�ǫ��J�_��b��ӡ@�9l4�g��s�#���'e塊�,t�y��Kx�m��i6�	Րe��������O�+d+�c��4Ć㸨�Vo3�+ݰ󮶖�EVd(��>W3ѠFz�h�ׇ� .��g�u��B��8]��+H*'P��7U�a�_�V�!�+��16��^��~$U�]z�h��s�����`�s�8�[���]��_8+Νk[�g�D����W�,�#9GY�[}�����7���"4O��L����M�j��f��B��E2]c|(��0������w�z ��]Tk��	�x�ĺP-F�P��/�sX�J���e�8���GU��%�I�,�}��L|�vW���N`K�R���Z�0� �7J��z��_����9��x����R�J�Tv4V��G��T��6��؀����7�9�<��񔻏Ze�	"�X����� �i���K!ʥ~>{Dt�އ����������ҁw~飱���3%�&�ۚ�����X�m��;���P5�t�0g�	�oz֜]��7�Kt��� F@0U鱬y�+�W���e���(t-x�#���-�D�J�����ի�+(8ߙ/Z�+X�����y,ތ*�������m�g�1�ǚ��/{"2S:�x����D����D�����y����j��A�#�[w�!y=�Z:��T׉�w����_��l��x��e���[r,���&�� }�:��P?�D��NuhB���[��J ph����ͯV��f��9��`��#��손�>�����on /H�A���x���e����>�U�v�b�|LG�h�Es�?�^�8q�׺/��)`ᮚ�>��ʖ��&V�O�Q7PQ��aS��UzR1N�f�� ӊխOȰh�IV��R_bM�8�Z��>ue\Z�zv�ͪ����|"y�=�q����a�Z*�8����������8���A2�"�R9F3�¹ϞC��k-ڼhA~)5�P��0 N
�=ް�v�s�s�*��fy<��ƌ�[�R)��#���ռ\"t�����s�h�̤K�NN�<M<#������;��+⦦{�|=� 5���M�����2�aӂ��vB�v<��Cm�#����Ė��s�-W�!O���8hA�(�7[o��RQ�2��6�JyU��k�D��^g���/�GM	@�<�q@Q�н��b�p��\���p��?�"�B&_�߸�Uy����.K��B��9d ���@�KUNC:_�8�0)`:٠�0h<��L�f�.g��g` IR>��1����<�E��Ǆ����|X?͓g�܏���S̰�C>�+^m�ÍM1�������/��W�b�~����vU����R��{��d��1�j4��UE,�y���5���ӵ���Y3�X�[�'�m%��V8=b�Mz܁�os:��b�K���q���jf�f����c����ܟ�~%Rq/�g���\�&Y~j��Vt�1eg}�>�b�h�Ixe�V���?v[%� :���a�:�5r((��M �N��1�v�
��6�S-.����;�����eR va�+�Ld�12|"J�p����l���wP��Ƅ�L2����J.Q鵻�g����	�.n��`��DO'���5����/�y=z(����$o>�f�^��^F����ݡG5�"�$�q�8�o�<֎����1�Lf�*:�uN�R=5�ԶE��y%@ ̤;����!`��^�C"�P��Ǥ9N#^$�-H&�~}D?�B}����.;�� ����+�s��Yh3ԝ8uu��V7���3~a��Ђ��Zg��El�ŵ=����c@�,�uF��t��J�5�E=�HPJ|��{�9A����:�w]�n�����GZ�SZ�\�$�dt��M�z�g�&/����r�/��q�.m&j���f�Ƭ��>~��A|ά��M"��w͒R���{�`��a����yS:S}�̘+�pr�c��!�Q��,s"���q1
AI�	����R�z'G�����l�*�N똇�X6�'֕���$~m���H�v��ُ��,�V��	!/Q�P@oȭ%��P�:t.�r�� }�&��{˽Bδ�t;vP�vg���"u�>E�P2E�,�L	�?�W��*=X~Z��?qH.�q�G.`���lB*Qy��m�z����,7�fl_�?? ��FtX6k�Ʉ��LI���,����;�#zޏ����$���œ�=��Sd3O�,���&8�(��^��Գ���/��T�Ew.�Ɨ�`�ɵ;r�^٥^ȧ�]�$e����U��݈��!Ы�-�r?F.]�^]F�M�թ׼�J��٨ ���Y��M@�¨v�]��:�E�i��s�s��iݒ\��fKo�AR遚ך���5-�(3W��R��;m�C���#��d��&����D��]Ave�������h�qMd��E��^���F�*�v�����$�@i�D�A6��1u��S��� e��Z��F��iø�Lg�x�/y}��E�*�m<�C����䏍����W�l2�I�oI��oY�T��{�rJ�Q��v�? Z�z�vѰ�ΟAjm��c.��>��ռ�9J:9J�/�k��v	*r6g#2��F㷕�/�ԅ �*y�!fZ��2�r�W-����\�2^�]��+��Q�L�C���Ue=�B��"��Vw/��xӱ�a����8A�}�������)�U~���=�=��iY�d�p�&��["���Y������V�ɲk,ݘ8���TY��J����.$����P"�C����m��^��I����A�k+�́z0\�`�������Q9J:M�7?V��vsC����śYW�@����}հ�\�
�־3���ڔF�US�MѢ¢=�儝#�&Qk�~�W�w+3߶�3S}�:���_���u�&o"��|F�(�^�$�j�n6q��z3��>���(���[�V��5�B�G���bJ���f���z��T�[�` ��1�鞗�e`���������J1&B�D��n�U����{��vt�H�Yi(�`��U���9�O�7Y�MA�
:_�гbJ�{Ź���ͦ����8�0zm���f��f���t��؏l�jfʆ��[��Jb�Dx ��Z�uo�k���S�8C���\�V*���.w�W	��>���Q�������|��f�G�p�ԏ�N���B��~"��4�o�Eb��?,�u�����Xʿ�)�괮6�v���n��ɉ6�l
���cqBÚ=Џ�H�D9���N\uf��c|`�߳EV�e��.UNօ>:(�6�''��4I���:���Po}q}�Yx���h0E
1-�=7!��+{�{���Z.1d�+ �.Ƿ&�H5�)�켍^!��@�R7�Z���~b�a�}b^:��5[�<c�Q��|"���e�NY-�@��@v%[�Y.��!_�0���ɒ�J�9��1�4p�$� '��KG*!1 Cm��������U��o����܍�|Q�ɲ��s�R�ƃ��]^m̌��ѓ4�����_d�L����s��*�I���>�6@�̰􍀲¾�|�R�����D
z���7D���W�H�cPƋm�Ak���� �!�&��0�&�u�}��ӡ�� ���'�@Mo�u9��j�ճŨ�I��c�1WyVz�qG��U�0
�ץ���з����Bo*�	��u2��0Q�7��+��TS���-��;�#T�6)E�ڋ
���	]A^$6������f9���!2y��y_J��~u�P]o��R�ѿ����Ҡ��9���>�*T��kp���g���D�QE}"v�����C�TV@�ͬs�������(4�\��f���G6 ɥ�y�2���ͥ`��}r�r�&J��R�4&t'*1��~Jrq毀ː�s�J�pp��K��%7q3u"����rh�ˡl+S��c�h�M��q��tI���	Л����_dJ�8C�M��jʹj�I��V-�:K�ΌQX@��-��g�k
�6;�j�� ��(��k���gt�14]��/-����g!O��)�]3�7>s��+��a���?cq�ԧ἖+���"�$0�g@�e>�'���2LX���?� YDܤ��N�Cr1�t\f�Br�(���璇�ne��w�(f�H��E����7���i��i�Z��\*�$Л�����(�����3U����ʃ&EEyo1�ޏC�?��j�e�ƚ�,S�6j�W� n^%1�������0����ڠLE��C�'���AZ��O�5�����c$�� �^��\�l�J�Z�*�Mw|�\*)�o�����k_dn�N7��[�����2���]��6ԩB!�mJ�3D%R�V����Ig����N���H�2�P��/k������x��כ�����ۚ�L�2�^ K�s��/�x<sהK��e�����u�|
p�ۥ��ʪl0o������7��r�l�Ғ"Rg�Թ��,P�=�w�9��K��b�/�Ӳ��y͆*��Z��3K-��X_ObYy�S2�����U��Ñ�I]g?>������u��3)G�$�4�?��i�<��(�� iEz@�ȏ�縱α���ݡT�C�#k��N���_8�{�����<C�)�X�aq;J/w
ԝ�8F�^j�^v<W��J���9��G�އ��V���k�2S��l?���Ɂ����e��u?>��<�-�] �{���&��c��S��>48�GwG9&g�I���)��V<��yy�J���� @`̅ڝ5Ń�Sx�i?#qCt��A�+DK~�4-o�55����x"9-��a�� }�M$ϧl�Q�+��3�����{�*�l�.��P��)ft��\ ��
���ŝa�ܳ�w�O�f�Ш�uBe��\�D�!�+��MQ���T
?T�U���N�s(���� �&=Y_�x%�E��A�7��$�s�o?M�d;[���T��F�r
R%��G��|+��V`T+�*�X�S����p����[U���1��K�Sf�:���wJ�w�Η��T&�r1�+!E1�(��e�Ĉ�W�ƚ���L�st�����{�V�N�`��8�.��Ѧ�i�*}*�r��{�:Y��b߽�PN�j�ǫY�z��z		H{���d¤�Ê�o1�3׽u$O�<W�H�Kd[�����S�UOI���q������ 	�H��۾y!��f4O�������f�Ö�G�6��Zw`��ՙ����v�}�ַ�㴏.�k���܈�N��0�ҌP٢��*��E@��3��B�t���Sb�`�f��s�1�e����r�����l����A�*�t�F5߁��e/1C����#��L�;�Gh̒�9��3�O�5��zo5�Ќ�
��}��!��_�U>�h<��}B_�\k�σ�,�6g 7�8��1i��Cvȵ��g�NC��S�:��5���o+b�]�64��V��-?/J����ƭ(���%����̖>l�D���f�n�\��]����#���إ_�*�o��u��l�Y����	� .}�%��Cd'�̴p��1���s��� ���#�p��J2�u��>�4I��n��`LZ#O00A������.�a�^�0����8�\�	�t$����0�-��/�т8���⇟�ӼJ�UJ�w���<�R��4!���.�� �O�`��-4���0dʓh��^�F�W��:�F�v�%h��ª��
�[��a~RN��+)c���E�Ƣ��j`Ĥa�ޯ�|��N��ؚT+Y0%R�H�T����D���\����,��h��NU��ϏFd
ׁ����R�bh&m�O��9��tw��#?����L��^C�WG��n�Q��L�PV؉��!�����\s����L��y�g�>@��0M_`����i���N~07���/!y�BF~��蘙�j�]ʄ���_���Q���>�O�!#�̀�̐��E�b2 �{@���ek�0�V����{ ��8�M��`�I�^%��\�Z��(�n��n����t�.Ƞ��ű6`��ex\�=���	���%w.1�0{�s�
,�X*��i�Ep�C������}3�*�W�`�����V�2�X�8�� �E���dm��;j	�����|�^]|���@>�e�є��\���t�2�����BE�f����d�\�?V�sW!��-�?�,~W�n��n�C��:N��Ś�!^�-�h�mA�>W�R����H�k�%H��74+�/I���d!J&�E����#�ly�u��v�P��!�\�>J(�j$�GH}+n{�< X6.�5~uo��\�����Q���?ۆR^�zP�q!`%�2���M5�F��[l���5`#�<���]�<0�o�up�Oj�q#+�(�Hɒ���"$	eEW�� ��w����~L��:ww�������v��NP{�>ƾ^P=~��R�c%�%�o��Z
.y-�.6O�(�B����%4B@燜UB��yS�V��T2���?�f|�Z��c�%q����ն�������gsz��o��`S*�_�M�,@/�,ye��]P^ւ�=��6�C��m/����`�o�w�t[���ע��_)�> �" ����Є� 2�z��&��+��̓���_�P�K�t�T�������k`}����0qjc۹x�3�n���,"�،��K�!k])�_%����\�Cl��B.�8۩=T�4��UmjE���5��!�a;��^�5p�`F��;2���v�̹c��qv�U�DHE��U]�$��+�=S��p�����%�Z�eBC��jEq(l\Ye�G�V�O=�������r@��_�a4�r��)tm���V�����h^���.�5[��+�6�T7���=0K�{{��y��4U�R+[�@� ;M*���Fy�����R�D�F&s���3
�ld#��=��l���+�J� lc�sd|�&� ͌�n�X��"2U��W��3YA>�@�h��SB2�Y�ϣ?�/�?�0?��7
.<:z��"0]?d�|�}bNs�QH�̭1�j���-O�%���[]C��LG��f>���Z��la	�`�q�ħ{n*�>�� �<2�ˡ� ���=���r	�:2_���9���m�:!?�}����w�I�'v��7����B<q�p���üץE����@��Ĩk�:\t�Sъ{�����q�kF�r����q,����f���?��� Fw��W�R6� -�`[�	_��4n��`�#��/t)�`�5�F(a���7�b�=&���?Gbdd_��������='��s�ֳ�M ������đ�d�~ld)^:���v(��5me5>�F�nO�x�R5��.0}m4c[��$��3az��I��b?�'�Qm;Æ=3���d��h�����y�-������xjR	�VwxZ��0�<��\�(�Z`u��i�E!�L��̷�\椎���&�-�د?�S���f���wOԚ%\օ�I���iM�P�H��ؐ��E�JX)j�n���*ӿ�z?��v���\��"'Zޢ�̊�����mo���m���n���|$*�*������=,���m�u��l�Q*��"����!E�Z'�]�	��m<_�~�����+x��1���iF��B>'�t�=�ii��IW��Tķ�j��/~G��Lc��v�����2�%>�t���w����mq�E�͛��K�w4FG���\1�K�ǙhL��%��˧F;f?�N7ϧ#��O\(�.j:Cv���zT�c&k/�6\�,�,�(k/!�+��G���`D�WK�T~"3��j��U�ۼ�B�4�A��Wf?yZ�+i�)Y�!����=��p�CU�yX��!�������W�z��(�� �.�ƞ1�m�%$�pvuщUZ��)�G++y�i�~�*�?(o�+�8��aaUs1y�Ԕ��w3��m�3(w��T��Ǡ`�G�T��'� &��No��m\�q��[eØ�x#����W�2�ɪ�ϲo�wV�_���2�zl�����#|��&pۧ���Ѕ��ll^c2l|�m?	A�3��/��BUm%)�$�D�뙨�-�R�i�>Y�c�R:遼��f����� \�~[C���i�����-x_-��T�*aG�$R��	�I ����w*ṏ����8K�Ĳ��iS����ڞ�oU�Q��z׾�ɀm�W�%��534�����`�<��:�V���B����V�w�����~���ҙ��яI���g⒃��0�mh~i^�b�\�cQ,�ۂ�B�ƠZ?��.:��t��vYГ������������Ӟ4�3`B��Z�]�m�Y������q��i\�$��ϙ,��b� ���)���:�(PiI!�gzB�Cr����R�ۿ�ߖ����{�c�Z�ۙ�ծo$r+35h��y����l�������!�r�Ȅ��nˤ=Kڠ�dpџ���2�~h�� 'Հ,�si�X�(�l~=��V��J�0	V8�~�����{��ȧ�Py)_��};�¢-���_ X�+�xlUbp�0�dܡ�#��2p�.8$_
˴][(;yY>s�x�&毺����ZTI��9�>u�?��->̣��V�a#��%�nM3�mJh�Oo]�P���V����r,1p��L�r��xX��e�v�C��g�+��@��"�C#�P�fdKU�&(�� O5ŕ8q�SL��F���`F�9xc��1�|v8��/�Cu�I9�o��5B�<�������(�����yq2�|��=|A7��(o,>CQ������ǥ�Gį���uM@����Bn�(B�xN$OKLD�j�a /�.�̠K�v}�R�nx�?�����	9NG����Ԇ�b�n���;JL�{�Y���t'�Ջ��J6}	!�=������Wbx���1jB��
u�]�k�$3�Tc�ր� ��*����g)ӂ�`������K�'�o�f.p#�6���2&��a4} �����*����߮(&��)Zx�R;����1DH[�����h��R��6!a��HN�"��G�\�V�\܉����7��Y�c�8ǒ6����2:x��p�"�D�@E�r�P��'�>\F\��c����l��F��BY
�'��tE�J#��'��O���Y^A�u�c�5P��U�l���՚���6��	`��K����;y�[��)���BT���sin��
!{�<�������P癈(�� �����%7_᪟#fȂ���c]+{����4�|w�t=��BN�۹,
`�~��(�0Y
���^w��������K�����>|B<��FN�L�'r��e��ʜۯ��S��� ����^
�u�PZ���y$!��p�X��`#���%����P}SUҍ�=2�r�ϔ�Q���[S@�|�1�m'�
��Wh;T���K����lR��+��|?��!��(�F���/B�\���,����Z��.+aT��i�;��)����m����i�S�vO>�Y�nl��?�}X���2�!��q-��x3��fc)4��:����J�p��Ǜ�-"��ϼ.�?ElLSp˪.�u��C�Kn�ȊÑ
�5��ϭw�~�Jή���.�[�	�u>#�Y�?1��\�H2��zB����!�� &�����"�W�^E��9�(a�X�'��������(���6�rRzG������#
~V��L��:�b�b���B�K@x���y�cJ���&�$B4��7�n0OAH��3F�i���%���m1�
��z���L�`BW�t�^�b�HX���lק\�w()Y�o�ֈ��߭��x,m��:UZ<掂��\�C�h]�*7X@o��{gg�����in�:�-�T�A��>^�}o��Q0�"���� L��L�$!��F��1�A�g�ﾪy��E񔲀�*"U���X�~V�����+�EK��2z��nV�N��p�D��)HeJ��K�ZC
bq���x�n���݉K������=���23�+�3���e$6�u�ݼ_15�Y7j_�s�7O5l�L�bG*�����{�C���Lؔ��
[1��8Ţ�Od�f���+�z8�*�WLC`5(��#����	�]�%�;�_O�4�}pf�&�b�lxX�g��w<9n��~�rKK��/rA�ʿ��p 5)���GPy��(.���~#U�%;]�S��]<`)#���T'�k�<Х������06�LJ�������a����?�Fک)�p��T6���t!i��s`�-�`�]5��6�� ��h&L��Q�Sn�1�ܞ���N�A���n���=�5��M�-�3v�����3O� Gd�Z��,؟�I-��T^/��`衠�M�J�,��r��i��w�~"j��]fXM��Lc�����q�����\�JzTgtKէI�pW�>8+]$�h=�uK��78|�_���O�<&��-�&��E莓^�u��y(��t(�燍<N�o��ĩ���YX�P38:�#��� Hi�F �d�S"�Phά�b�-�q.�y�+~�=����<:?��%W\$v��}o��w���'�LU�`y!h��o�!o�˔4��T�ƽ���aFX)�% ����x.N�Y�[��LfQ���y�	��w��_J9�ci�H����9s�A���LDv�A�q�y����4�c{��/��8t~Q	������<��l� ��?��*<���8�:�Mna[h�֫
�J�b�wtPrw3o��p�N��^\}h 0�v�n���_���Ä�:eQh<Ѫ�.��c���9�m�v�p1��V ��	�m6	�X�ҕp�CW�+1j^hD�w@Iŭ�D���(��u��ޛ���]�D6���M��<N
`Z�;����6��]I1d�lV���ĝ\�v�3l]Q S�ʲ���#ݸ���2��n/VLH�D	Na2��� �,�s
&[aٿ� �+�WS�E�]ث�%hw�+��p�]�2�1_~�8<Ɂ�"�q4=\�k8Y�W�H�"ob����P�f��(��c�:Pdi��[ށ��836s���\��5������4���iK3R?6@pND��t7���4fKX8)�c7�;�S�r�*p���f��!��{�2͈o�B�b���[2� �f���Mn�fr>G����2��Y�����w.��һVn�k��֘�@ R�a�[t"�����7=�)<�펩��߷_��[1o�����ȁm;�����]�Y�lEo��N��Mw��2�S��ı����0���Z4�����59� �u��8Cg�!Ձ֟�J\�-v���)Z��"���s������CՀ���Y	7S�6{i���N���İ�C���l�<3��B3 ���T��o�on>�dߛ�U���ñ�d�N��	��eUX�GT�&
-E�l7��ތ�� 1O�c����\<Lr�'x婲�P�b٨-��g�ǣɞCXt�7��L���BSW��dB�lʫ�WC�Q즠��[F�l7-�HEsn�2��=����a(�ь�^Rpr���]�����u�1��Tɭ��.g�:+�;�Ȯ�&�o3�4j' ��#I�bS�kVb�O�(C���Z\�
�1�8�m�~/�L�wh�.��Rࢎ�7H?�]���?�0^���3j��`�W@f|��5��m���`�R稶��MMY�B�B��E�BF���(z�G�ݶ�Mk!L}��G�nϜ���X[��a/��7\���z�ڧ����[:��;P%4����6�B�zP�rX�'>�.�E�_.5�o��ː�F3�dx^�L[Ȑ���u����g?\�>1��Gwrx�fU��%�,C�V?�e���O��H���~���SK&��1F�YކN�:R˜��TƬ匌�<��J�]ߚd���'AEPز`��/@KJ:k����3%�y~+�鸞T�7u�9��L�=��2��=��5␃0(�?x��ޏ�v�!�� T{2�>� � �Be�&�vFjW�t�h�C#�"�7�5
5c�� ���4��/�'�����7��2׼SAW��uOg��\��B�L��+Ő����ă�ʡSF�O3B�M�M�|K5���>F���(\ab!�S��ˌ�7�BΑǂ��*n:��;��R��q}��F]�� 
�F��yL�Ur�i����	Sۖ �~�:	�f,�W��O>X��/��.BG�\JI&��� �Zi�]�
t?����TT���K+35l��#j��46�L�Uȶ�J$✬��')"�B�ia��16t}\z$��U�A��0���{�^W���c#z&b�6�7��&�����&,�|��$��r�=�i�E�~w�� wL�eG�[/����W����~�{��l���?C�bƜC�t�0�9d��%7%�8����������[Sěo1Ix18���A�t�G*�z��=�xo��Z����L�Lp�D�X�.
b�L@^�jX��a�Q/�R���ǈ3���{�q%Y|��{un�Z%�7���b��W���D�e�g�E�y�sKM͵��8	��k�=Ss  h������}8�+���;B����r�q{�P�%�y� �sp޵B�� q�e�̟b�]I}."+��CC��CWu��GÌK�;!�����5P��\ъD��K9�Q�		__�Z�b�^)%�!�b2�8��̤��ɒ/\#tV$DyG)5c�4���rhbI;�#�;bc��X$'�p���5��9K�3[������jH[���c��L_\�)� ���3t �%�'�l{�8LUR���Ъ�Ka˰I�i5(�Kܘ�XFR'�fȖF��^kAK����<�7�P�:�!3VY�g�b��o�۬zlI!�ɘjа����4���
i�����L;�ڲ�8��	*Ųa�#�$�_T����3�J�����dTZ��iN���C�;I�fYι�0��S��\A�D��S]�N�T���+����-T�Q��S��Ox��|��#^����	�������Gcu<� ���u)ū �u����?��-��θ�<LCK��Ip��n��]z��K�e������|k�D�O���is@Hv�������l�/�j�����eo�iŬX���"~t�"`��6AY�h��
�x;��7/��D1���{�D��\1@��}��z��_V��[������9	C 3�_�m(Υ�� mFʟ��K�-Yſ�����L���9Qu�ش�P��.�%I�� aٲ�(����9��-�������B񯩘�dC]:HW��֔���?3Y&���O]F����C���O.�-�E�7�w�M+�ǇM�7���"��J��g�Aa��v�����b{�D�Uޞ�;�"?q��%�7{��Rl>�$5~~����̢��h��Z�q3��8��P1y2yn�p0S�a�)g9�S�����5�Ѭe�y��9�{*<<y�B�z^��2��g��&�����ı�$��^��:fp&�A����*I�� ���ؤ}c'3������̌�Â)�Ώ/�]������K�"��u�v�m�ޤΊ$��&�ODN�`` �"t�&/�̰��t!�N��zZ���+��^����#���su�H;����B��D�GeAGWYi��F=�\~0�/�R�]Y�:�kUOM���_����݃�|�3NΪ�r�q�-R�oc���)��+�;VoW��!=H�"�c����]�ؙ��ٌ.�K�Ϸ׽k�v�UiR�G�J��ې�5m�|����GE/bH�˭��ϳ�S;�$B��.]z�&��cl=��T�坈�x��M`rƗ����3��ã���<p�Z2� �/TtC(��^�T��xw�D��,[�#�S!�s[����@[}����H\�@�qkxU3�=t�zk�����z3ܱ/'����b}��]��~rN������̼���zhK$�Ó�,㫥o�����`�?'+�i�q�~���aq݄�m�g�K,׶=TU����1t�1��Q�L�SE�K�C�"g�����G.N�":za	�H�8��M`kL��~6�E'��t�艹uˈ��	A����q�4�{�3@���E�^;�lr?��Ds-�H����-���u�{�e	:���Й���9`�g�1|0���q��!!c�x���Z��Km]�u��sn}���k��^<�,[���G��@*�Ky����G��%Z�ٚs|l�Ҹ�����<�ė{����X�ȑY1�+Ⱦ	0�6�;K,�����%���i�`��[Xh=�����F�ӐLGD���}����ޡfEfZ�iN��l�c�1�vf ���a��C���Qӧ��@�ۋ��
 fW���=��l����Qv��em�Ѐ�P%J���=
xE�����s��6�K(�Y	b�+4]��5���&���M��Y)�3�ܠ��[�6/�#�mZC�h���e�*�l�}�gQ��
�u�g�+z��cSǊMŗ�v�_l̇A�!���?A]��qR:�>��tɝ��NOv�w�����+����2��"�}�����^wiW.�-�HWm�X�b�V�Dw�{��M=�K��82樏jh}��{ ��I<0#1<�ᢢ��UѢk��9�z{:���BF;I���?�(�̚�z�Uӈ̲[9�^ʏC19k�SbT0����,4���d	����ѯ��R��sR�Ut)��^�`C��������1 =�ܥ�ډ8����9�Q�4�Ndџ�a~H>�������!��M�g���'��g��L:/�r���͞^?���	�ϰ���g���O.���_���%��(j����%
z"�^���/�J�L&$�agM[��
N�qN��+b�b���?&@��]�ʫ��.4�m;F����&�7�WŘD����?��^O
(��+��:pSB
�Ac�e���%:��Ev�Y6��h��pu�`�=�����8��!`�L�#���n�6��aZ7�/�y�6#]���i�aԫf6�.Ή!���@�U�M���?�iΒT���)��
�$mn��v2\5���K�W	�l������[!�K_��k�EO,abQ�"sx�yis�P�/�v��˷�T�5n��s��ע��ꇋe�	��f�ђm��۪�q� �x��$���s\x�e*�/X.�a*��H_ǰ��T�"vn&��F.�\���i�eU���y[�g��b��Q��&
X�_@�
�������8�]|z�9ד
[��&�kV_�u��;ez�졪cJ�SL�����i��)b�.Np�����6����*�CB��>ݻ�Sv��Ųg�h��})�V�a�E1j�N�Y����n"��0b�_o+���zjȆ���I6�~M�@Z),D�T&i� R��{2������q-v0c�j��<O��\zk��d7�zD:y�ݛ�L^���,<���_P�<�= ����3�|#����w��I�u�T��ŋIЎ5�8z�)����~��c�o�׏7�mJ��Z�+=K.���|is����hfej�rk:;C諸�ۢ���Q���l�����p�ƴ>��($�����H�
�3�q��gy
&ag�J��Љ�Dzg�ġU��w`�JS�{,S��Xר�J���@V����磅E���ł�.GT@��\*�B�e�ks��	U�_��3�I�c�$���k�d�F�:�X��w_�F5R�Ia[%$q�J�dm�R�%�����0�)сV�Y��7Х=�c�'�@�=���,��W�F�d1�¹L�7�s��f� ��_��rf;� ̹�����@��I/Y(�t;���9-��R�B���o:i2g��'���-O�b*)H�-蟷)�D��2���3~����q(��������K�� %Kţ���K��w�������n�a	)w�*q<�T^C�H"�
̛��ُVv0f�H�B��k�u��z��+-�.U�"ɭ6¹����X�i>��?����;3�lߩz�1P�*@����������}�*B��7[��y�:��\�E�p$b�����U�&
|UF�CW�&����0��)�8�!�n�d:I�0,�7�ցqKC��+��]�H��M�X�-�m��^��mb!y���?th��@�n����_���CL$̻>=��?�G}���w���**Ԝr@�43S)]0��Z�K�yH}�#�/�����bϣk �騦ٷy�׫�05�Ҁ!c���I�U�G�=�:\��cO��up	pʯ9��QR��B�f.V���|.��M��>u�5�O�-v��3|:mK�3+�j�]�ڠ&��2��ӌ�x��HoH�A~*!���*�O��mоuϸN��졊�o�d��l����e�*�������mV�y�b;�O��ɏ��CYS�D��+�0�C�Ns�q��ZZ�̡���ib�@@&��,i�i�+��	'i/��t ����
�b�_>61��z���}�]V|f�}F��NJ��%3]�� �ؓ�5��I�r$ԑ7��XMI��������GH�x6
��õ�x��ΘU~��#
|������=��(W>Vd��T�f�3o���E�ouW��C�n�4�\��FB��-�34�i��G~�`�MDc"�@UC
����@���N�3�~)V 4�lRRS]�m��a�1 e����C��G҂v%�#@66�Z#Bb4�v�[}}~�R)�ѳ���������Wk��璭����@�0�S��sv�~y�J"1�(|�Z�P���ϕK`<(3�jӼ�3Y`�vr�=���HvF�B�B�K� ng���!㮝(j|Sj�u�+�v&vDłn�z֢o�]¿]�/kD=��p��/Î1�J�N݋�:���-��(��Y�a�_�"�U^�Ѭ̰�0�k�z���X�~F׭t��cˎkk�C�ok��ZVF��a��Xhg0ԕ�A���-���qAfK|���P��h49��X-�@�淅���3��K�
˿#wn�����G���}�U�0�iT%��M��l8���X��у�M}��]�+��>�M�l�g��b wm�3)D����0��
+q4�)�$� �0���!�54J���㙙�*1M?����9Nw��X����PٲÌ-�aӉ�x7��������#d�;휧!��P��"��[J����Xxs��h����nL
E�  Y��a���|V�9��&Յ1��ZX�J���<�ٞkz�6|ܔe�����CdJz$|��\ftre���E�l��f<�A�Lc�Uvju�h{�~����U8u�^<�w�q�:"�'ɪ��%cy(D�R69mzX�ѕ�x�y䜀�!`w�F�Q$�5T�Ħ���p@�fK]�3
��7��K�+��������`$�{w� �7N��>���&װ9�p!��%߬���ET�_����Ä({�~,�lM���IdO����u0�l�.�Daa�	Ѣ�+i����t&\/n-�X$%�'��������a�>\��>��SOs�P&�>E�c1X��8m�QR�W�/+��]g�i:a��%��쑥G�Y�<�12n_}|�e��,�Ԥ��L�#�8 ����Mv?���N���*�j�0�4=��1��b�mJ��o��w���M�;�ݢ�p�7�҄��$akUh��C{i� .�N�l��բ,{��>�}��	��L�%�O��e��PɎ6 
2���|�5'Y/�:��ɜ��޷�ro�� �2 �D"� /��}V������{o�� F����ۍ�׷�Wh",q��o����V�-w�I�3"@>��@%� �?����Y]b�qN2���(c��zn���6�߈�&1giR*ū�kn�Se��G#�٩<�.h*�W[�����.���nE����&Cp����/|�Gg�rh�=e�L�#�އf�&�"0gdq������|�Al�H�N�a��CO`L��B�6������t8�H�h�5��_�/Z3����sL� Y���5�"��~���*��6�-��̋`��	Fs�p�i�Y����ʒ�]�A�x��6�G��T�u`�o�+�q�����6!iuH<��J��Z�y�ݻ{��I�%e�_8�KH ���m��Ӱ�kۡodA酌�Nڊl�I��Lmnm��O�ޒ���+F�䡻�^��Ϧ)G�	Z����ƢW�8�!��V�rFms�3���݂�Ij زq�^���9��<,Eڼ���B$.�ذ�[>\Y�?�1���2j^�'BM��=C"R%w�#�����ѓ�k�W�*<�|aU�P��	��2�sJ$�Zs�H/���f)X�۸h��f�IԂ6=n�"P�	�Ț�_?'�i!}���4�22(�8�������/��/+ݑ5��"���O�!���=�λ��[�5��������M��ĵz��嶬5�;�T��y��ð�ѸE�k�Db��t�r�Q��"~/��� �!`Ә�U�ڏ1����oD�/���r�yM(�Wg�v_���%X,�1���?��;��D*��.�s��1���mRk�!a��J��*�#�<��Vj���Q���C���w	|$��ʳ:�1��.��Wzx�Pl"����22���̏���o!�O��K�2�a���\�6��e$�y!�u�5v��O(2���P{��B�*>D�[&Lu�#�IP�Vȍ�K �g��XShn�m�#�X�ԩ��$V�`b��>l���8�3<�L��Ӿ}��}������[FT-��BpL0N���i��T��8�-Hݖz�#������.��� k)_�@�z��`~L+��
������I�{���\V���`b�dk�f>�H#<W�L�K��3X��/�n�gr�ƥ�$�S�|Gn�C��T�U��Y�
<�)�������hI�\��v���+�n��к�y�?�xd-����B��P�f�ѿ�-�0;B;@��Z ��{��� FM�	��Ѧ�Bҟ�Pv�wA<�'W�b��˖:�TK�e��м��L�����,����Ri�H����}+�+8t�:���`5������D�@o���4���S^�~������6��w_o?x���\lhl�)^
g�̇��fL#sRQq��W�q�L'�q��)��=�go�?�`�� ��D�Ap��lkp�\�VMvX="-�O�?H/*!-b����1���[P�O�?�2��ȑ�M���Dyd��U�!�_�-���q(�N��5�w�~�2����� ��0��8fẕ�V����\QP7R?�;2/��M��,�E���*�0(�e�� �)�A;��J�X0z��'db��������{5S�\]�2�Xy�eT�'�K��L�;ݳ�xy=a�2����f���:RlYg��t;����.�(2i�$����<x|^�����GQ�:I���_&`��,i8��q����L2�	MH�*��c�Zⰸ��*v���Е�����j��
*���d%�<�f�9�9��ʓY�_��H�r]����'���'2Nԫ���^[���z�]����f�-��-�_A�B�UI�"��Q�:������3_\�ɀ�X�N����w;p.���S�^vu���8kJ���c�?��\jI��z"%�+�N���*���/���=|��|0� ����1�֓[(�n^���A�dw'Qz}�;�$>��t���@�)E��Ќ)N�b��7���d��K