��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0����_���3e���ӌ,nc(�B��N]&��;_h�'��g��ײ��A�U�)SWn�(���I��jy�i�	�)�j+.F���4h@��2؊���d�rqD(�nJJ�L�%�U�C tD�=��I��E���;o��+`�Y[����|� ���I�\�_R#Z��g���po0�o�tm<&D�TEHgC �9l�=,��;%Q:��p�J��y�ˊnӺ����#���x���<�����`6�E�l.����p��"0�f�����+�QKH�����|������O0��*��^ɸ�tb�l'LM�Gr��UXѐ;���"}ɗP"��j �X������yn-�[��dZg��h\�;�0�j��\!׍��YL�	���#m9/Q���U�',��`��NN&v�bʯ���V�Q��n�RMt����gG~�r.B�sŊJã�QϪ�S����ž#;��T����-򙉥��(���<�?��ղ jp��X,��頀.�}�\g�E����T�'�3J�<�$�\�[F��@��$��������0��EÂ|�{;��p���K��L�j����R�$����6ءT�	c����f� v�p��_t�c@b�-�.Tf,�����ܤ�gi܄���FG�\\^�C�
B�}�ա�F%h��э6̿����n�h� �-R5��'ݏ+Nn|�Y�
��L�i#��B��[�X���#P��4���Y{~0pfYҡp�U��Y���{�TL@���{K�
����8�N�yo���d�!��<51��t��eaُ��?�?��?,�Y�䙕�y}�g���K�bf�:�5�z?"���Ɍ�:b�?���/L�S>�nz��Cg{���VLؿi ŝ�1����ڥ��cq��$y�)e�#γ#^��x�Q�� �X�#׬����(����M�,i���!a��i�L�	��'�'#6��0����ә{��s3�-�v!HJ��,�;)�s) ��iՄJ��m?]�(�^ lI���)^�����P���ۣ��s5�M�m��5�KB�r9	Tczn]��5���Z�q'a�nvZ���j�w��_�]�A���}��Ъ쟟%P_�`�t��a�Z���.���l�L���a.�И^EkR&3q�@5����E1"�,.Іa�Y�G�S�a#����� �0)���{�Y�i��4�f�V��.@z�_v����6�m��A+brE.���l�G�B�IZm���
�	6� _<-�]54! ���T�O�����*�}^}<�m�i&��������c ��V�2��%���L��t���uc�xJT�Ÿ�)�������������aL��?=�"������t���Yq>;U(ʳ���^ZX_�bs�[�r���tNq���7��1G�����o��L$�Sv�o�7jnI��o�s����!z�Mt��Us-��ހ^L�Ⱦ���l�D"'�i�t����ee7��x��8��h���~���j1h��E^��t��c��Ĕ�}
D�l�1�ٔ% v+8�@O�C�|egm'�������0C1���C�?��ka@�����DVq�5*���.�n#fn	mt�KUb���&����&G�Վ�+��%�d����}��%A�Ǣ�{:��D@��Y��lq!�X<8�'�j�*�k����ދ�q��̷7�b}��1�9@lU'�H�n�2b,�g�u��CZo�*�=`+t�5��؍$W�w�����+��t�4q`@���i�HC1-3Њ��C�����m'��&��N�� �����Mpz�ew��(I�g�4[D+$��\�4��ٲn��Z�5S=��7C��)�����]v�gf�O4f�1ص<�4N>��i6�a��O���j����,��2,�;?�z���A��>:����&����-u&��S�5COu�rg+�wp���M�����I�X�Y���D�=�h�}�j1	K��lƳh��/E�K�p j�Zd6��~��o�h���{t���3�-���`�
���f��8��74��x0�iA�����W��wۿ���VƂ,�n2Uٽ���vU=��Z�{~�\�g�R�+���Y%�1��;�z��J��l�?�)� Ġf~]Y@yr�ty�e_4 fP��G�3it����P���*��g�6��-y��Aq6`�I|��g�_X�zm�fy�����0�ga��1URy�q�˼���M{������B�Ã�ིY�Q�!��w_��(�k��ɸD��<�d���� 2����|fיK��-p�K�����(=n~���Up��Hy��]������Em�5��w4�o����008��F�ﲗ�Gǹ(�����
^��N�	;��h��'��~;��=�#w��9�ut�s� �+y�.�کYl�� �:c2m��2�.^�QAVX��Z.W;�j-3�ނyP�C�Y�
��'��X#Z�BkHE�gy,��6RKR�S#�9\�t^�EZ>�A#xxa����41�e�o�ٜ����̫���y^�H����ƺ��i/�u�'�N������o��;��$�:���8���V����Z��z:���_H�,�w�G)