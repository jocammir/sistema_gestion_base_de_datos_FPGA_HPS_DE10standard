��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����{`,u@=.P�.L-|�̯�	�恫f/$�mv�Qf�~�{���,���[� �dwk}Cp�dp��Oz+��x�R�#O�W��	ӓR��SG������k)��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0���]8#�T�����w{[V�VBcĹ���D�
x������j�#��G���t���~б@�W��]����7iW;��&q��� y�+�wlo|�AV�%i��)� ԫ:CW��#`ƚӊ.$���~\�|�
��`�S��hL���Ao HaP�G���/0�7�\C��õ� �w��'*��o[�xaU�C"^^׭x��댱T�J��=F�څ~��+�9�Z�.��Wh�z�C��@��H߲V;
��+��1X���;�8of���5q�z�/$*@��_y}gJ�������I���	�3��R�z���O��\uZG�eD���h�!�[If^3��Ι�)�u"��6Hmc� 㠿J��(򬣣���x���J{�:�u���Ӈ��.�
Ju3��T���ui~���m�1�]y��,N v8��]s ��}����n���<}��C �?-s#G)��%�*z�\�^ �����0CGz��<G*�k[yΣ���P�=�s�d	|t��4W�uﳫ�D`���x��c�B�WZ´�\�Q��Ԍl�ݿzUj����^�8_
���q��%n�����:����mm@=uؤl���8����޲���c�mJ�7Z����=S�w
^��z+A@9u�Ћ4��������ǾZ|<�vӤ�P�\pMp�{۩ܳ;��C�P���s�pI,Y��߭�\�p�+堍�̮[�˲^����"ŉS�И?�F�T�v$=u�sK_�y�갠��Y�8�{#��[�5��F�Д��R��CvE%��7>*%��������oR�C6x��8JUW�;��7gX
�(NZ�fL\�E�"�˕]�\�������N�v��-��C\��C�Ю����dO�N�j���[,�!�O;э����зՠr+}?=���Ͷ7�j��y~^��'�(��=�YZ�ʸ=o˷*�c7�@L��좳�F��-i|��r6����-���o�4� �N���?+�+��L������$�8����4Kp'�Pݯ�C�_|Gk�+�r2�2LO@B�e���N��3��� ����M�J;[l��;���x�H>���T�S����~g�b}yU�(Q ^,a�-f�R�X�0<JG d���Oy�f�v<E35i�=zk���ݭT�u����V:$�ʿ��a�����Y_��4"�2/r�Ե�f+{fج�5dm&����M���f�նT���(�_� ��+�qG�����.FZ��#�i_���v�Im��r�5[����\7Ř"G���:�8�$��&'��0%���*�Hx\S��s���M��Y����*��E?{�|��BHF���� O��|��9��#K�%Xr²�@�M�� Q_T1�c��&�a�/T��U2bU2��0 G�3���VhN?4.�e��7O�	������$�cM����S�t-��vURN5�Ea@�I�Z�+��a������,2���D�_v�G�,}����{^Ύ�����0��I��1`̢1`�|F|��%�ϙ������?"�[J���7Uh�_if�5�v� 1�s��pәb=ty ˀ��)��E.{X��'Z�����T�X����h�� ��r?2�a$2Y�Ό��O+B8�]��r]�	|���<�����d]� j�`���Eo�V��,����6��͋��Aل�J9m������"l����^\Z9�u?2�%�(W�j+��M�[�%��S��^A�����Dj�)�DNP��)�}��+1���BKS�/�ڼ$�?�?� �pU|oX�#�mv��T�96g�vKf�4y���2�t���71�l��1Y�pN�m�O)�F�@����)]��l4��V�@G9��M~0����#1�Ûl��\[�Q:���z��S	,�4FZI��U���� U�����	l�L��_�c��r�x��F+Wfc(����A.9yD�p�����4_<&1��"/�(r��P�n� �ݮ$�\�e6~"��)(�v��<�\��c:�d�K���6����P��)}?@�p��_Id��t�q��a�r?�' �ڈ�a��>�����;�~pqwD����������޲&�#�2z�����W����b��D���ϩ�\?� �a��R@�̲�"{���@Rj���I>#	���"�'�:4P����"N���U�<�s�{;r���u�%lN�V!�5��S����ٷ�S�1$�֑LUC/Nn��U)#|Ӄo����=�������}��>WY`[xd�(ѬʓԚ]��6��t+��'q��F#���
�}��ю�|���I��*�x^_۲M�p�ٺ��VǷS�+#�"��,4��W�ܼ!�|0'����U
2�A�QY����M+�Cx�a�^bXD�}�i ���&�k�c~e���<A������Z<�b��������ɕiψ��n�Pf�0�-1Nd�&��+�&�׳��⅚�4@���x&�l,A��3���>�87��
�M��lc���\`þ�w�/����@�~��N���w@Ny���Lٰ�}|v;�- ��(A�z}��BE��d��S�I߉�Y�Qx�k	R�[�: b�~���R�VI\Fi`���x�O���Vs�N��z�1U��Ʊ25UQ�1'�]��d	�����M�P���2I���/�DU�������f��w�t�Bu�
��+ːz���Tm�N)�*eõBU����?Ǐ�!�Ɋ������Rr6tN�!�7��L渵>�P���3��;�a�X��g��C�"�9tN���y�<X�H����|gm頺��֦R��R=w�W�G�� i�Y�=�nJ����A�&X+�{��1R�OyR�Ж�!"	k��b2�]Cޜ�(�=g�GEo��&���(**�y��X.K�d/��ry/ˊ��-���-;��2���I�	��E�( u;.*�sբ�n���S [�� ����	)aq|=kG�[C��]�� ^�:ٞT��.*�_��n^5K�����
V"���`K�mu*�;o�s��g�-�������5"uB�U-Y��4Dp�]������IO���m��=i��w�"I�����4�ݽ7d�4OP�Vhs���3(���Lø-|�÷��?�)�՘`�ӳ�+`���&��>��$uI�3�/\�In��m�ȿ�����ź�Dzz�~!.%���^�q��T�C�2��A�`����*dȑ�$���"�L@A6prse�'U�h�X��d�BϭU�4�_-��Y��������'�UU�4�nF�ѨY�>AsQn=n$���V�o4�ޅ��m�!�l�mQ�<Xb��q>��ҋP���g>|���0�\�ZM]�Σ�q��8��bI"yP�P�g9�B�حtB�:gx��ŕXݤt���59��|O�s�k2�sh)�~�/Q/Ϫ���w��U|W�i�gfŶ� ��A5r5�]95���8n����ný�� ▯��'[�>�aw��V���
�� k��6��l���m}��.˄�O8 �.4���#��*�G���j}[K|��bV�"����ܷ�'�M��,��<)Y^�j
�Q��"��8��(���o�=]����4'�z�y̦B�^�:5�#O����H����b�|tsNf�9F��6$w�\z��%��@�d�OĜ9�c媼U��y(l��#����(��m�d��)�_@'�4��r�A#�ݛ���v/�D^�#��F�J*x�Nc&#`��B銩���#��z�TR=߬.�2�\��-�㠌��\���zqjӟ 	|�Ջwax��[^�
�<�"�[HP1��y�oG�T(=!�@�g*qP�Uf��$�+G��� �YK��}��������U���D�l,�^ �j;���خ��]��?��U%$��,d���k���Ÿa��^�Оw&�����ඥ��[3[��՞�Olmq�FOk/D?���Z��M�� *zcT�&E�ϱ�ܬxȪ>@�UH@)��S%K�Ϫ�y?1���PN���߫�pk6 |�����C���ػ�.�U�htC��pf�U��!���:�S>0��~Ų�
k� ���\J�$�;m�0�@_�m�G\�`�v3c&B �oD���i?�m7�����_%�$9(i����g[����@+��,�D��#
��Z�t�Q�Q�(I�z�����R�j|��v�D��O5D�[Mޡ5��Π�0��Ű����I�'�g�}͹��![�n���S��

ا�H�b�;4-��dS��֫D���(M�\�{�?t߳�HIx��Q�$XTQ��ifA���hJ��av8��ѷ>!/Ő�9L�)¡YI���Dk1��G�$1F�\�� ��;<�l�d_D᧺�qi�c�=M�9c�PK
�9AhO�&3q����Hq˝��oqC��6o���m͋C+�!���Y;�̈2�ѣ��j�2�H��nl���N4�؁_��t��In�kRDi�\�4;~󸚴�Ԅ8��Y=K�xP�q|
IIV)[�瑲�4�Z��(E�x�A�-ڛ"�����Q��D=h���o��H���u�5nZ��ٟU�S!h��H-&}�[�1�f@��T��#�����I:��襄���fj;��,�L�)��m�^�Ԉ�d�'G�tH�he)�.�5�tb=�3�y��wt�-��9_;-NRO�?{O����	R��I�-CF$(]C��v-49����gxt@��c���'$�D1�R�8-$�u����o�|����$	�6����݁ːQtG�P�(R�R�,��!���/4`uP��⦸�;����^�d�rq��F�<�L�^1� `��6��&�%E�zvq�V98�m���#�5WU�
ˋ��j0�Y�Um��Rc�Ag*i�ӧ��2k�������5���+ϣp�DIR}F9a����;��׭�k�١�G��ڊ\����~6E�6	I�%��Z�q(��"�zp`X��抝�1��n]���#�JN�|[~Р%������}�(�f,���6Xq�A*��O"�| �j+"��l�m�q zӊ�3_G&�Bq��xۢ�y�B6�4Ӝ�� z�{�7�C���0��చG�K`6Ac�����𾭸h �AC��u��` ���-AR(F҄2pv�&��[2����AZa��|us��B8}�d�a!�:�@�V��PX���f��0�p�f�=����Yj �#u��XJdk�&8ȄON�s�;Bɡ�����}�t��#�e'9�����`07��{o/	�["�د��21PFZ�=q���s2�
���u��#��*�R#��Ya/DY��iF�H�eq��S!B�Pȳv� �/�����|�r#���#�0��m�3�E��� ��b�S���H�8�?�U)2�S�
��^H9M���G��f��|FզmoP1�܀l|׽_H���9�S!%�Y:�R���K�owh�B����!79'n�J:���D�*�ur���3�8Wez�@4��T��z�ف��S}-9�p�H�Ȉ��:X(�c�U�X�՚R��N�IiT?����b�쇫���|�����9\���-;��-iN,�=: eǬ[(�N_r��^�Pu�D�Js�������(�doJ��6���
�"y��SP��_>8a*�v��R��=�����2�� tgZ��	��7�a���f33I��KZ���a	�ux�7�G ��o*�y���J"G&F�}~�,��(��oNQU�Mj�.{���7�ӝ<_�T�!�p������X#ǿt�ϐ���ۘ�@W��&f"(��2g9B�+���B��c���f�B��1ngnĘ6~jpjjEקRqc��`73�)�	Z^��:�I��"����g#���	�y��fȮ�;7"ø�	�����ėv!Ϊ�n���h<��ݢ�3�"�x\Ʌ"'�h- IۋaQ���ê�5�Rep��I��қC��
/j0���;0��T�r��*�n��էg)�'Iޒ�|"9C��1�O7�&�p��_NL$]�$�~��{�b�W�H�"��(�*���A� =X���X1�j����\�1�T)J�D{�p����KSC$�Ov���.�|���_Q�NA�<(,}|#O晳k��h@��*�Մ����!�X?P��V�vi�����֕���
aM8?T�\����Hs��αhG�#� �3Y-?L����}��} �
~����N�w�j��v�h�#�D�7Q�{*^�ǑqQ��<�#���Սzl>u�����D�0A\"@)�<�\�\+�6�$�~�r���W����<su�7JRA+Z\���ڎU�	tX�W2�J�T�źVvj|������%j��O��"
 R�q�k�޾/�w��~�;�MU��[�4INO����Q#t�&�"4�V�
����S�z�b  ��5	�jاD�:�9��7�!)�7��w)�?�7vXu|�E 3�,�|$~%"*�_Z��?�YG�|�]�BR�x���t���8_����;(���\j��M�X��M��r	�[��P�ѶnUѹLγ�\��z��b��=/�o����4盚M4%F�'Zu�.��&���{F;�"�vz	�R|6��>r�7 ��5��]�ܔ�v�v��� ��(������P��gHL���`~��bCLˆ4��tQ�*IQ<��%�d��u���1á�E��2�.��p�q
�x)6F1 n�J�U�����М�=����1�	������^�L�*g�(W15���do+#9.`�}?��v���U5���wc��4�]I���e�#ܹ��0ϔMx_X���JΟ.�[+�<�#�$	�t��I�-�ڳ�Mh��*n�#��0>��k���b��M�E��`���E"�E���Ϩ0�rR���?���$����X�9ȱ�P��^a,���%�8k���q�؟���,t�W��R�����I��,la~���}XQ�O�-�m��^w���b�rDD��!�U����:b�v�~�/���Q#���h�j0#�:�˲��+l�,sz93�;�#�h���Q�'%��u
_L00�BiHDBHھ��m��3^��rJ�֋_e���X���7���� .��q�~��v��k�1����WXJp��ï�+�a�<ٕ|n<Dȥ��d���Fw�3�k��9���e�5	D6 >lLq5��Gjy%H�~���0�B�JJ�4��58C�l��N�D�Rܴ"?�{O����t���Ό�N8��˕�b����5P��0Y�{��?��Hd�����;g�Ъ�p�Ą*���=�K���ƴ"��=�F&���.}��vs,^8��MHW�F��%��#�^����8���s���PD�O�Iq�%d,ɡ0c�v��Ϊ�'3ޗ��gfue
��8�žᣱr[�W��"l���rHuo�v�[��S��gu�m{���1�K?0f8��PI��/2-]�-��l^O��ϤcɆ@z�4���Ӿc�K��8�I�<���>�xoo�ѳ;��_�Ǉ�0s@���_>8S�6?jҟ��A��
��qJv3���i&tuZ����X��x��$i*�BL�H�����̐���ۄu���>+���&s��:bu��� dt�Z�%(�y����unk��{t1��n�ьT�R0�uc�F��98���T�j�H��m���}�w޹���ﶧ�'��z�x��'$��l��;:�� {�����G��5_�G@y���h����בſKˎ�cGdu�Ud{�����p\�ȣ�����h�ky`�L�\ ͅ��y�E	"~��u��lr�g�Ο�7emKc���@���a3��&��V�O��� WfY�{p��\�~��44D�}�~pQy@所�CQ])�ȋ��~o���7�>�����_�j4�<yN��_�����1��PMiǙ-5�5�X ��&�9a�
��r"��>���XArY3i���֊��C+�1�WCIl(8��D��n�Jj���a��q�k����v��?��"��Ƚ���<bG�Ź�)G'_�'���aq{�Mܔ�fvq�1A�􎇒�H&Aw��:��X�q�L�x�B�3���֛W�e~�v1lKo��5�H��l_y�����Oꀛ���
�Idw����+'��e�Y
�ġ���q��	�R���c �����Cz*h��M�ƒ�s����p�S�����%s^I��\3�^84�덧,Ͽ)+XX��-�k�;�-?A�5��z���_�
���I?�!�޿�.g[h|��tC�{\)*2��`q�Q�S�ô��f7�Pj$2o��oS��s%�u���h�n#䓘>�PQ�Й˙�Q��V�P��)���˖�X�Pq���4�6����ht�g`C1e2
��X�/�Usq_�]$�Qŕr"���7�+జ����1����ߐ�!�	=��6b>km9��S�R����5�x��O���z�:�f����P8;�¬_�5?!u��YB���AD���L.#�󎓇��UH}ѫ�.�3Ik�[��X47��-p�K�*�/(�ZZ>,�+�J�^�� ��/�9Ƕ���L5�}��qK�}�0�C��E��/����2K����aW������iq�_')
	�T�q��Jݦ_+18Y����/�ߵ�|�O�����B$Q�C�K�)e9�v�a�5�B�gD6�vU�m�C�]����E��Q��S�Ri��Eu7����c�_�"���7�_��_0OE���D2�C+?�8��p�����a/���&��d��*<��q�B���ί����	��y[�5�wDL��^I.����(el��:F����˦�bf�C�?�R��������U�2���}g�"��ρ��!c�A?9�c@Īb��h/���2W�����P�p^8�u�?M}�e��z�L��8;V{ X�\*�/�h������hޅL��fz���ޫ���9�D�
 ��wE��Q�����r�k��� [#c�+��j�5t<�J��g���+ʫ�ܣg�v�)ͣp�^�m��T�k/Y!c��x��Ia���>��I��wkq�/Y����Yte���"j�9%콲�!mt�^k5�#��h"�8��vnX03dz�j���7���\DX�j:03S��:���&ª��Iي.�Y;���]K��Ÿ!��FL��7�BƷ,� s���v�/IHX�#�{7�,�Sf�M���j���a�gj��_�s��Kf�o������������'ԅA�Z�X�j+����r%��������2r��U�������u��hw[�.B
"�
 y�\'*�G�@3�t�DR��ڠ�s����N:��u�T�cryo�F`ε�)��$]��&��yn�gAX�N�/��KZ����Ҍ�Qޏ�4�ؒ:�� ��w���%�!��z��@�sba1���������3�?�yh�M��w�]W��g��ѝI���xވם�i�x���
�W/�P�t �p-����[ƛ�#��6t:����d(M�+��G�����,6���C���mJv8�U��l�c� ��vS>7��^ڼ��S�2��ݣ w��"D��,�W�V9�E�P��O���Y����0�퍺��~|:t�}_[t�N���
�y�1n�|�p>?Z��4=�3�'��̍狧�ɑ(��U��y$�pS�0�ꐾ�1�U�rE9^>�S�
�֐�g���Fi5����(���a�Ec�/�EO$N�V�o��4�2��%l$D
���7�̲cG�^��DH��j���
�謷�Z�)�i�ʅ�����u"�4��7���3�yhA��Z��S�����l�*�d O�O�ZYݝ~����Zi�QE�r=�W��ǲI���1w	�[���3���x4$�л�������_}L���yZ]����b4W���Z��f����:��VC�������ϐNofo���nh/�������O�x%��6^c�- �`jNg���W�1��7�<j���5�e����O�m��ս�ۙ�5,�$�x��P�A;�\��	��_nP�K�p�'g���R���$�hV��c3�����#�w��ZJPIDnm��.��⌃�%�����4��d�&����mp���^�%�'o�a]�~� ҳ>s3W��!?��e��.X�}�p�ķ�
S�g�"��&��j��B��]��?�q�kF��1��UA������ak�h`B����1j9>�R�[{�����V��h�Q<��$-$$�s/��M�J�&_H�~�HZ�#�z��'�'͙S�SuZ]�⥞kKߎc����߽��.���]D���m'�� ��k�)�z����~4����SQ�Ը+�_"��\S�9�b���,n�H�W����6"��n�Ir[G~�B�ʟ$y��N�L5f����Wni�y�g��W��R�� ʿi���8lPQ8�Բ����Ih����Ѫא�����O��S[���w5�t_�c��?lj��jh@!���	o&d����fp�Ʌ�I' ���)�
�Yk9��U
*���'x;����6_�X}�;^?�&L����$��d#g@���7х�(�3��;���bǭ��"�;ŵr��ʄ�ka):�f��,��R_y�F�Zf�G@�����V�����>_`�0`k#�������L����HIfP�`�� �OnG	��"����	Қ%!�换�������gF�d+,Hs};_�*�t�ѩ_4���餆��,�-��K�P�zѬ��������C�HaҤJ��l�o,�މ됻5~�%��Q��oD�ٜ�����w��������᯸�@smͦ�����S�ܯn�:�+2��6��+6 �%UA��^ծ�ߍ�h��A�e`_;I�FƞƷ��(���H�GO��8�U�g�dK�nM54d�|z1�!�B�L1y�����)��?�����]~��Q�2�q��TY���<�U6�g)��Rj<��@���OK��gV�ll��ӥPԗ��b 2y�1��Iֻ�s�!��`��19��c*φ�2�.�?g��ة�9� ��"�y]��<���b�~�%b|p�R	_��N~G_��sfMc�r�b}����A��c����",��ܳi!�<Ë��3��yF�M��Z�A��.!79Q-���}������'S��~d�a��"��}��U�9�r�M���ΓRoι�"[�8�:���ỏ��֣aw8u8�Q;	D�8a��u�a��$��ǆBeߐW=Mz+9�Ӑ�m�DRB�N�ܿ�	VY)������U��~�����֮^
�'���?dw���gI��������R
�'�}C>?�钓,���­��_}9a�ԉ�.���~�Ζ͞�z� R
�o�k2�����
���؍$$Y(�?��71�Zԥ;|��\AM���� k*���Bh���;��F(�m�sa���:q&?��tԂrrDJkg���%PX�q��m�7�=�s�8e{mmKNk���d}�v���y�-�$��z���O�<؅J�~��|j�n�k��_�SvW�V�=kQ�m�`&jʵj��V�/{�J�]��u��cY]����u�l��G��S-��~IK�,��l�l����4-���U�ſ1������i���x��Ŀ逋d�J����d2q,�HgX�����x��\���㽇{���3)M��veLB��;6��n�L�&��F���0m��V'����t��"b�[=�o�>��;'�?���y2g�`���n�T��=E���
[�|�)���B���/�E��3��' 挫�r��a�+�{wt/O�N�����U�"ڌ���ץ���h��][EpL(��S������(!(�֏��Y6�� �[��%�1�ݾ ;i?]�uf�`v �\�fGnSQ��7@�8�[�O~���3{nW|��P<Z�u'H�4.]�:��H��\�}��fQ�|7&'��6�w"G\j������"PF�&��K��s'�>�AeL��ђ֚xlw �㨙�s�&��M�aYt�>�-f �%0�Q�eA#P�uؒ�$WI�I�
�ǟ�)M��ĂM���;�V2���}*����rՌ�@�
��Ud��#ƿ_��Ӥ�T0�!�q������6�k�.�D�6�D:��ep;4��W�>Gރ3���<������m���' �#[��I�Q�&U'���&�2�W�o�_B#x �|= �Td7�њ��%��|Ղ��R������ ��-C����УMq&R���0����W��λ
| -w)�g�����q8�<6�3d��W6�]4I�&^��4��9rVtĳd� �bu��~x-��ᰵ+��(y�i��N�����>��'ऒ��]�O�r�;�Ў�9�xH#`C�?N���ǫH�\��j�0�֟Ё���2d�
�1v�J�$i�c� �W �����i�������4ˉ�Q�r�y���૭Z��%�I�l@(e�I5��J�*�k��ᆍ}�d�3������p���� xQS�?���֕����x�O�[gxc��K�G��]����-J��CY��v�R"	p�0�{����E�SW�����z����m`�Lֽ6a��T@���8�⍖�����fk���iJ���N��J�C�۴xs�����e��� ��X����,�q���aC��� L�7�5���P zq@C�S�Wϣ9z�В	*	�Y��Dc9�p�t��P'+��t}�N證��J�!	Բ��̣U(�sZ�dgwJ��n��~�Gl��K�����>s?��q��%��[���|�|f�/�ؾ�,��Jly���:�ȧM�#esr�&w;���+�N��^��Ɏ���,�oc��*f��j�O^Ǵ�ώ�|�gb�})^@(ǟRQm���W/0e�c;��'�ڐ�߾�`& 9��"��,[�3\&ӡQ�<�B+��4�ӶN�⋀x���I�,�69� A1-�#	���EX.���-ª	�=I��髺��ԩܬ���P)��dO5��3x�ԑ��w��*j������O1�FV��9�o���6����V���j����M�;�2_�
W�*4��A+o�3�eƋ9����m�-�<ן��[������qҪM_]ovS�)�yc�{����>�RZω�ָɃ%�檣?5n�.a�*7y՞�83,�e���K��j�n ��z�î�g$�q�������3~��McQ�lƇm*�7���*�5��%���Hڟ'_��D�@�J�PFQ+����d�T"3���8I7I�.����o�[����1f��	��f�d����������Nc C��?!�z�r���O;��9`�Xs�[8������J��ѸE�7�~�a��r~-���j0���#np�P�hBL0�}��T���S�96kW�/�Ǎ����E}�x̩����T{�� � Ы�ẘ`S�b�����*�� e
�T�REW�&8����b�$�aȸhT@��+?��=b�e��?AҟO��I�,m����u�V�E��I̩��n
>%]��	��`�m��H�r
�F�һ(�;W�rE8uƣc���a�M�����-j��%6{q{��r�Ǌ��'�[4O�|ciI�O��u-,$~>���"p���r��`������z�ZdB	�ԟ��6e���w������A�-�� MH���Bh�0�Ĕg��_�b��.�$K�9��4��!0I�S�����d�����b�G�!,W֓F�mO�9Z��4&=P�V�-�D�b��0
RDc�g�(�f�q�)�%�Q������9�~Jƴ.G����'nnƲ�#��`;�c����GG�MHtW�{-��=u]H�R����C ;�<bsjh���/ɊF9��!��!nvv9��
&��
^�@�Ҟ����T�d�d� 	�X��v�w��;x`]�BiM�b�!N�9�]9�neN7]m�� �Hl�D�_��������+��
.�[]���T�ۅI�o���e�gkm(#w2�F�akv* &�"
��yM��>�ŵ�4�c�����vI�j�����zUM�G�+	����-�v-�R��f�S�F�
P�L�?F~}���U����/��y��]�'�� $ٗ�F��6�ݒ�K>���v|G��J��.d��vj4�Ֆ�w��f햇1��\BQ�N���c��YI���>9[��p?C
��y�oa\-�tu`W�d��:�'T�.Q���rMn��t;��h��	=��)��p
�}s�$~j��d��#��H>��{)!���̏�M�5m���8���f�ZoZ���*n��	bD*Q!�(��j.'
�g���#����¬�dξ���!�z���m#�j�.<*��]���J�$6L�4���$�����._E�6P�jb$��r��|?Q
l�u/;>щ��)C��������2mf�v��Q�0���@C�/-��\rihx�Z���s���jBɥ֥Z���&ܘ6~-
9@�`�)�#H+�9�ӑA��t�J�z�i��-��1=�<�x��	W�*�[�Nlj�ibэٞGhHt\��!����H1H~����M��z���u�,��d-X�݉G
~;���g���K[�#?��>V ���x@ߕ�H.�Pj�&��i�*���ߒ�x/w�7lgp���Ԓz�̤z����>r��z�/,���t�M�ĬZ e���[WT��R��_%z��m���+��aCe³oO���=�/L���9�qH�����r���9O��<Ɣ�������̀�mw0x�F�r7���*t�(�p;?��b|�S�vC����I�J�&-�^���z3$�̛02�1����q�p��N�n��E��q摨/�r}�����)�pqB@�Pk�K���F�u�����P�������w����1�e���w�X?�9e!�1�CY�rn{ֽl���3����n�m��2��B!�2ܤ�)9y
1��~ay� ��ZWVO�9���q�#������,�惰��m1�������Sm�j�(��ʬ�T�����h=�����8dE�Y_v���,\��4rZ
n<��A���_E�_�>�;����c�6�`��_r�᭱����V�[�J��Jt�M�T�T�/8�==܉�?X�1'8���_J��X!:Ddǘ���~�2��B�3��]�m�F �2��<���O�\=b�h����P���x��Gz��b���{9�&�N�Ͳ{"�>v+�g�>���i �g¥W����L��QR�8�����_*�h�I��u���*��R�� ����Tz�BY@�ڪ���o$�~Jv}\�8��%`S{�]y.��������8�f��C��.��XS���3xW�H�>@��	�� "�]��:&B1h�Rx+-#��Ż.Ɍ��zƓrk6,UT.�/�r3<��%R1L�K'�MmH:��D�����h���%x�oL�a�gt�V�7P� '����/y�w��n1����F�[G�S�b�c�y�eU1����<���ࢉP�ww�KQ��>���l0�y�*̤|�B
[�or1��3���n�k�(։�!�ݳ�[4�tw�.�@�,��:�S���q)O	�	�xx�zV�)�������Iɴ��6���ΦOqa��R��Ds����c�����UO4T���ӛ����y����<�~����
1�ҧ<<#o��Ͻ��r��iGU7��!���`��x�S�4���Χҝ���fz-�V����; ���(�S��D�~�ع=]:��)&��KVS��{���Sa��?<��pw�2�Yzkw�r9���S�{a��_ LІNi}���9�.��b��nR ��[����6|�g%�ͱm��$��p4T_��Ly�[a@�<�n�_�?�¯����Yˊ&�:%�'ڍ��cLW[��NF�L��63Q����(���Ԅp���,hE<~�y�+7��gj��V��F+	�W�m�_1�5��܋�uyS����mXΉ�=M�x�H�����cϬ����!v���N�g:���v���*� (��H�^���a �����;������#�yK�D��Q��+�(|{�B�갯�T�6������Evb�`���67���^��P����
�+��nΙO�P�|�!İy�/p�q��Q��q��))���U��ݟ�8���.��I�R������3eYݔ�jG�U��N�W��x�������_�9�uS� ���Y7����x��إ��@��w�	H�<�y�����Fn��_ �,US����y�O��*�jwMw�KG��"6�vs��Z ^,��^;�^���|3W�09<�`�䮮���qS�Q;�ؓ5��H���y��!hW�Um�zn�������ʡ��Ā�4:��m��2
�插ߒ��n�9�=��ƈ��������%ઞ�C�2�	��][��u� xq�R���X�s�T�Z�Fx����e%�ժfs�zi���k�"�-�?
g�y���!ײb50.�Hm^�rNS	�{�ἱLa�'�J�F")����q@eKqf;fZo�i$���� ��ty��PQt��d"����IE�Z��w�
&���6��炊���/�����L ��`��K� �Tî��eU�C(1oρ1Q_��z��G���bC;6RI��Y��`G�/n�59���|����L�5��f�����6�:��8=��d�\�t��C�o�×W@;��m�~��o�4�;j﵅5b��T������V!\�v k�[x�%�Q�T��d�ƶ�����TQ��g�Y�ÌƧ9W���0E����̉	")����o���[,�Y��ƾ-ᛗӰ�4bKx��e����41ڠ��Z�ya�tn��!�+�2�횈�.����r4ě�UC�$\|Pϕ	&��]*�:F���P��3���BW�`��"�f�S,��k�jn��Ć����g�V��H"������$0����*������%��N����\	�=Wi�8�S������k��R�>e.qx��o&�ak1�FԠ�ٯ�6-0��8~�pX��T{g��Fa����ɱ�S���Rւ�c^�gPphYS�p
̿C���ȓ)`d ��v�n���p����ۜgQC���p�-��ny��C�����7���qv�J�lN6��6��dȝ���M�o���\D���j��\Z��W��Q���cA�IU+�����]�iM�sX�׼$�-���K��JXA�ѭ81�s�|���>���QG�.M�١F�4���L�lD9r��˸�[%�慱�]�0
-�7��k����s90 ��*Z׆&Er`�+#���-'@���C�rz�e"�+ŉ�7��z[�-}������܌D�6���<0���E����b`q�X��7�M,�#O9[&�U��/���9��/��q=g�l�֟��.{����ŕ�-A ��[~a��N0e��8��	��{Ϟm��1VX�Q�-��<�qY:x��v�������e.���Mѣ��%(p(�"�D�g?T��~�S�;�x�r�1�FK�3�O�ۤ@�j��eV�� (ϜK�W���LVPQ�!+�4�(!l�XM:sz�R/�1*��ZgQCc'�+�ǞV�m��
g�����W$J�H�\�DP�"�k@�h�*�
��ڦ'�V�&��a��J��)l��S�d�D&�xMO�,��J��r�߀���{�y��6ͅz\��wͩ�	�u��¹�w�c���^_�1��(������Ef�ZGdPc���Cfg�L���S��@��y��ʵn7L6�4�T�o.R;$|��p{Zʞىv_R)�jl<!%��t��
Oo�J���T�|��@p ���}R=v	�*�ҏrWO�I���A!$��>��RuA�����B6���$�`�*��VA0pѐM(�L���lYp����g�g��0��cN@P��<��	ƴ��W��v@�WM�����8|o1+y�G~�b�?#π�QU���=/}����/�Հ��E�A������|OK>����cH�%\8P�ʼ�T;�ev���C������o���t~e�r��e��Y� ��|[�>~��p:b�vƿj�y�]y}��`�{��*ه�/%���&�s7'*|��K���M8�ߠr�Z<_���o��"�+_~�,\z}B��ï�K:5��D�{�.:s�~M ��E��?iӐ {'��Mb5N�և��C�{��(3�^�6mF��ZMY��c�x�<YUVd�������-F�'6c�x��pؚ3\v_��Z���|���ˢ���7 ���>�?�P?�ӡ[�������/�����9��l��Q�v�y��m(C>e��)/+����JG�v�8=��7#h�y���H���m�`s7|�g9�o)*Q�7��G+��=�=�Hdz:F��7�̹��I��ѵp'��s�70:(�	<�,�`��`��9�uE��6k)�u���{~v��5� ��<�����%��u�|��M�����k>b�i �O����j+=N��A�7��[j���-����M�(3'!�8xf�9W5ή��T��H0
7�b��>ҺkFj��6wu����	�p����yY�������#vxDq�Iʽ��&:�b�J���� ���XXߞ�,�W� �ӥ1JC�=�S���_��A�o���ː���cE��t��[r5����)�t�f����2�P�\��S�{����jٟ�j���梴��&�MqMȲ.^�=��=���/G7fl�"J[؝!M �Nt,�ke�LS^S/8�.�7baʲw8(��͂�g��bZ\Z�yf=��.��|��H���@K軻Qi��9��AQ(g�N��=�򇕫�q��ʂ��?��?��e2�o&<�����H_38tF	�G��/��3�l�&bA��ڑ?��	l��!Y�(ӆ��eO�i염�s�2�-�ʨ�-�_t/��Q��u)r<	�����#����E�*�h�7a�Ա(�lo�JKD���}�0P�˘���"/+JK.?&i��;���/ ��\��[<��h xG����֥�ޭ��'�}7"��HŇr�²��G�&�]l�.#��{o���܂5�1�D�BX"zB��fl�c�ʴ*�{��]2z�����B���4��+Eyp۹X�m�hE���*<r|H�j���i���˥7��=4��q-F�X
�v�Ԍ�~H��߰��w�s>�[�Qa�.��n�!0EI�s�j}��QQ�@V�QƋle��.^Fp�'W�ZnsȳҮ�Q���@:-�q+��}h�w�V6x��k�4ޫbeOjT�m�x2��Î$��&gU��ܵZXT�X:l�3�z��s��G+���D��p�E ���% ��"K��G�����v�����l.�>��H{��`�Ck�VB�H�1��&x���[�P]
V��vɿ��i�1�/�ä%����9��K�]�e0����P�[a5�Y��O����;-g�������G�-��G!��`u�S�v�f"0n���'�����I��&��pk �;}`�t���A'��ѳK*�
3�8'(���/�<x��&_GR�aRZ��ha�O�
-��n��gJ��N_Â����J�s��b�Q�A�i���'�� M錭��'))���_��?��F����3��p���f�ҷ�#Wq�1"ʹ]ó˯�?���t�����奀�;�hQ��N��r�J*��ߺ�8�����b�$�jpn$C�α:06�ą�6��}��/�v_��&BN�A*�X|���H��{��(�ܱ�͏΋ޢ�g6�L����N��^�,������I���TQ�$�A��Q�|@5�%iIa�z6�.��`�|�,��I���;�R�"n�c���A�ZJT+�N�"���5?{�^q��
,�ū�d>�F�O̅�^�^#�"�Y-����=@]#U�8�����;���B	VA��g� �;JSE�-==/���DW��>���w��AL8uʰ/Ԟ�c�=�>ŉ`�	�]��������qDhx��{LT>��J?�����!@U������R��WIy��O�AN	lY4="z�K��H9ȼM�����y�{}\�/ȥ�0���R��*�^�D��s��G5=�q+.7S�\����J͜��&�`o@����ߞ(R��ھ�Qۓ �a ���ؗB�~�tT�}}H'=�-�~=�mx�	/�ç*$�������y��b	#"�uڊLǮ�'�.jגkʿچ�8_��o�o-!_�e�A�����5\{�n@��0��W��*�y��}�����3��I�	ɔal'�v�41����kk|����ԡ�;�[0��?�JF-��ƅ(u����y+,����0�,�9j(��,���IE
`g�.s�{w$'�YQ�
��<�����t�a���#��!	R������d���[��hc���d�I�$�vZ�Z�s[�Ǜ��C�#�����~��yg��ѓK���||d���LEpJ����Ì�v���\qO7<�@�3q������AD��I�I¯B 1i������_��g2������D�x���5���9]��0"��}�����Řԙ�S���K0�M
(7W���؄U��}B�Nq.i!��X��Y&����Zڧ�'�++K&
�_ϸ!"\�y�[����n�c�0�cF$��T�0/UXW�ZeP�������q�؜c����K��p�8*�N��m�a��[�����[����`��ie޸�wk6E2�XX�|i �~1�����|ci��E&1%��6 �֊�o�v�f.��� �4���U���?0��]EL\��v��6�Ly��s۠e9X�O���Aڟb)�t�"��0zddI�yB���cC���)P32��2�oX筻�8����"۹6@�J1����1n���S�=Md���8���0�6U[]7�\Z�||ͥq����ѱ�1��\sϞ����TD��V7�+��P_|�����)��'	p�5�H�C�w�m`(��7�*LOY.$�]Ct����GJ�JZ{'k����hn����\t";^�ݠB�1t8P�B��%�/�F�ސ�'̖�M7��┥`}�PCp���4����>k���4��6��q��MY�]�;��Ý����97��7@=	rO�(���##�M��֩7T�c��2>VN�̧��Vۼpؤ���>�'�����@Ah�?�/&��i�l��0y�A�ޫ�:�`���,[[o�:�C�'��C��K1������B�9g���=�b�w���z�MRv�)yeb�ũAΖEK}�z]�'�{ �/�����6 Ĵ�����Od<a�,�3�����K�$��;!DO�mUt.�=v-(��Yʔq�V���Yh�۬?�����Wv���D��&m#\M�%�Ǳ�,R����10�EU�Pq>�)��"M��,t�����l24�#�2���s����g�P�nmpwPQ�GF���T�*�:��baδ�0Ҟ9��;T*̾t����>�dn�Ulyp!����ˎD��sf���G�� س7%�s�R��X���g�椛��|oN���{V�D�FE��?O��x�[�����%;=ON1�4NG(��߼Gr/�<�1�'�	e�%�$��X��n%���$=��G�-<�T:	f��~���cz��_�'�����Sl$v�aT�פ<��y)8������h������a�4���vv�v��$���(���Q��ї�N��?�z\#���f^��_�V���:#3"�֭#e���W���t�� [�`���i�,�?:8	�ByuK�xS� >$�ĳZ�8KU� ������ƻu"x�s�Hu�k_��}�M����9ZWPĄ�క��)���h:��LHcf��V=E������y�����w$��d���N��9��\���D3�6�u�>t�6f9��ɕ�kJ�*����5�9:yL��妈#:���o%�0Z��40(+|���sY+9U�YI�P�}uOܝ��1Y�*�F�UX=�=��߼��"8�.���c�߯O]��UiT�,p-L�-�_��� (�h��kb��*��d�}�l�K��d6@��"�]{R1|A9�kw��Ȥ�*��# Lyf.���"�#��$��=	{'>�6��K�/L��j�f�9+�~<8i�I��q��S�L��5;]<6��5L�P�4c��h���<�`:*��Nn��	�Z���фxG뇦J9u+��Ix�����,ŉ�<��W쒑����}=锲B�e���[=��e^��[,rꉗ#Y�����O�b���[�j*q����7T�s��<����b����g/cr0�xdŪ%&��X���dAt�H�a��P �2+�H�&Ѽ�$�e�����K�Ș��o!+c��/,aS{���R���L;�6���)3�+�E?rgX�$PSYf�Ta巖H�!�\΁K UߦD*�Da�J�C^*��yK�N=W:~�ʌ�cGW��@�G)��E���E�7�5����s��Y���c�f�?Tѫ�Bm$!Y�r;�veE��� ��ʏ'ш¢ٲa��Qe�81�{c稯qVV2��go�]e�s������L����ؽb���/{׋2ZoR�Z\�{�70�����h�\+e�\� NNq����u�	�]������ ���_��O��{CG*�tf�P��Y�3�F$��S��Ίa����:�{0�(�E�uQH�x��K;-3�OV��YT��d�����IA �):���JV=�-$�K�C�dl��~s�[9v)u\ ���� g��(	�q5���F�H��{�Q���Fs@�S�	� ��6P�[Wz�^���� �E;6�o�W������k�D
5=�|�WjZ��'�§�k���'cL�c��?e�������C1G߁�pW��� Zd5췿���򺗦���0�-H�j�E�{���B"�[�a�Ϭ����$�r��+�!�Jn���z�Sn=ⴂ�K?}������C ��p���+J�-Iݵ��@�6Ov/(p�g�Y=c�sy��1��;���b�R�"(���乏���� W����������*ʵ��?8�Di!�ﲈP#��(`�uL�VoD�C��[怕�b��rA���U�/�ס�Y3���G0��B���_}7W�:����-p�	q�P)T����5436 �J�7@	�p���+��R�1m.pJb= 3(��)D��9� !�( �ټ?�H�����07��Ѣ:��&���$ �˯(�-�q�ZQ���	��pr�w�V��gT�#0�g0h�BK�Qd���8y�DX��	T��`A
��_�hYeQ�e�(�3����Ul�|�UN{*��g�!6������k�Sgr��L��|���9�CTEj0pvF��u$�㚍C��Ɍhy��� ����) �1q�5�]mE&?�y�&YvAU�����X�񑒂�%W�w���|u�7A�B��wZ�� ����Ol��p���qǰ�Ҩ����B/S�Y0'���к�)H���̺?�F.�m��m�HM]�)����Ggu[�D���:�%����7���� Ti����=uF_1-)r'V�Q,���n����D+~�	IiC�ԍ��U���%�Zaʨ�ެ�B�2�k� ��>�ѡ:��wm�mɺu����d�:��1�П#I���v��Ĝm ]5��������k<�O���z$��f&��[mƌb�b�{���X������xm����p#{�֭Y֬X�T��n��(t�)�����k���e���<I�O�t[Դ&��QcC�4*�U����!$4�t-z�39������!�?�w�I`�����s0������c���t'ovq��<*��
�D.0���|�ΕMå�<���HK���U<�v�K."*���K�Ƚָu�������$��R����R.sEj��̇Q�)4��ލ���� U�����f����lC���8�:-/�� L��4O���K-��ẁԀ[�J�ߠRZ�&&@Aڈ]�9���]5˭�NZ�Ҙyi�L����u����1y��KKR��M�v�2'���xh�>����`��0%3����ȕZ]u��w�UdjN:�P̇5�CN�]�:���EE�����m�hHe/���D�I#m#[�0�>'? �\ޅ1*z�ƨ��v���|kg{w�R�'2�����B��Ψ<�aw@�L+t�c��a�� ������`팸�T�(i�_R�p�`wJ��`���|`(V�j��<��+6�5�Q]h#�ߺi�盛A�r{��.�������[R:K$]|9�<7�_@%���SS��!}���"eȉ!*v�Ί��<ѩ��?F��x�;�1��h?v��@�_(Lw�;#]�8�k�}Gz���L��+a��ܬPM�er����T��wFb{�	�@�-�>���p>Q�E���0����V�o�Hg��B9C�����x�A0�J������	�HO+B���v�V'�X:�
���~��I�1���l0�����P�s�RD8�ͺ���@e���	ѷ�g��ɮ�_��#�C� ֵqx�z��8���4���5N_�C���>I�ʫ��3�hdN�,T,L� %}�#��}S�"/[b���l툤Ou�����P���"���#�"�&���w �`)p»�m�ݳ���DZa`���{���ڃ�H�� X$5>����j�[�?��8,c�V(�ȅA��e�&f�M�Ճ.}�SGC���jƾ��-�ޭ�i�h;��|�� u$0�;��l�C-1TH`����N�����r&�e�>�ze����%ǖ�(��+�ܥ��lsb���Z0��Pw �Gv��xs�����ZZة���6��q���^b��l�ͪ8�B1)��(������X�mj�}��7�����:��@8����}ǈġ��;>˂��T"�7KO�2/�[��mH���Wk���Sϗؗ��7��C����-F�n��VIrD�Z�)�S���N���r=S�w�[��2��4_��9S������n��N2�vV�Y�*E�$[���j�i����,h�GU�^�2�}�_"��}�q���,_7����R��n<���1>i��ճ�U�'���`�t"�˫�ZgG�t����!��3�8�@��P����ץ ��ݽ�@l�Ze��`��n�3S��i� jR&5�x�\�����Ǡ}�8*���������G��}���-,����_>,Z]e��K��U�)Z�\c4Hi�L�x*�$�3����# k�9Ǝ�����s)�`�V���w|\]��R^V�Yd��~䳆��ж�!��-H�i��� ���/!�WH��]�ߌ/��\�4��y�I���a) �t�k����	Wˡ��jg����>O�ڄ)���y��>�J�/R�^{Pw��r��)�uJFإc��I��O����65AQ�D*��V�	� P�T�(��6�&��=�CFYuC�W1�>!��H�>�`̐l	����ֹĲ	����>������(��}$9�����&�\s�Q��2湈xɶ��	��ɷ���h���ӹ�=�D�T�����N
��=]RD�Y4;�^>3��"df�i�̥�3��mގ�X�����8��-�q0��m+b��@�H���I��oP9�	�?9��lL���ė�|���+2M��je��-U�Ī�C��G2�6ۋ��^�|�֝��VV�����\���P�ۇ�I�.oe�u�yt`^Q'xq'd�J�ћ5��e���K�P��v��K��~���#��NU�\q��7�"�c��Ex>|�GfH͎,��Kn˾�� �P#Kq��uN�{��WW���CY�&b04R�k#�U�î�i��I{�<�|����k�o�/�1!`�a��瞞t��ɛ�U�.\�����3q/=���Rz��$�z������ �W�?9�h�HHe��c�Ae����b�iQ���w��6�� ����p��g#�"~[���e /g"Ou���9"�%d��r-v��4X�rO���Ϝ��z�l��%%v;$�������� פ�/��#���*�Y��/���gD2������� �|��W.)��� �����7i.iN�2Y�9��R��H�q�E��ͮ8jc�E<]Յ8^��moh``Ћjp�Jj��[%�Um�B�rv6�+�� ���v#��x���j���+���e����k���j ��K>CSW\H2�����ɕ���`����%���zx�W�1��+����!]ҧl�vN�?�Ar�.����Ҡ�1���`iqx�xQc^��S�����sr����"�<6��cJ�)�\X�P�Y�e�L����߹@w�a��FI1�}E�8}hp��7-"�C�ɼ��_7���$�C2�0]�b�=���Y/B��2��-�0@��P��s�O��쩱�TN'3B��CHZ������#e:T���r aO_ؠ	��F?��bc�s���K&Z�C�^hH�M�ӏ�F}y���9FHo>��u�9:*b#DF�zs�j0��o�u�<	�[�|Jx�v>8�S'�P�L�*�b	�+�˘�Nk|"Y�}��l���'2Ǟi�7.s�G�g�ub������(��(��W��p�ԏ×���\���ǩ�I����+:x%-R;�G0=�t�Z�q�V؅�7Kb//_���n�2�Pr!t���%
�6Lf���h����R�Ȭ_ȳ���{�Yam��?'���3�%��s��_�u�{Л�6t�iGs�)��L�n���΅�k��.aD|��,��_Sü#~0��Yׅ� a`"':�����Pv��P��"��?�_I���|�T-���S�*M��%��9^��)����P�)��UW�:s��P�p6�oW����q�9.�׻��C�4��1(��ʼ�Wei������S&k�+���� &?㈔�~����?�>Pe;5ڵ�\C�	C�&)�D�B��]���=
� �N}��SI���.�چM�!�c�9ol�"�;��I��S�����5k�B#iW�ʑ�} �u�+�F���=�+N"�q�h�u�E���?����(��~�2$`"J$����E애W�R.�]ɰ�7���e������*}5T�ν��&��M�ϧlH8\3����ƕ㍊6�S�暯T�>͊mm�^��]}$\����+���G��G��\)]�G2����W{BX%��W~�:�qﲳʾ�����m�<��z��Ӷ-$�*�Q�:Jm�&vD�W�%��N�]L��|�B�zA4�,N�f�26q�7�	�GM�6�.���`cIw��ٖ���d�XO]ϐ$"u��(]���H�-�"�z[��&���E�k��l�cZDm�k��Z�W������-m���9��m�����J�Y���N><U �0.�l�#� ����Z ��b 3�g�_�������X��|n�O� �̸�^�F@���@�����X�O+�^�~�����K&�JRp�
%2�\��b/�ˮ�`���Ɉs|hY�����c C��o��
k����w��>(����U_\�F��U���>g�"�Q����z9Ut�-)��,�=�Y��Ul������BZ�>�(�~̐�h~uZ/H���NHx���F����í���/&=�d`i�������zop���&[^�b��[��TWgM-��x��S�N0sd.��\��%��弪����D��,����p�g�I���t=��A���o�����s+��}�(�O<x�M���ڒy�C�U����^6��>�J����B�1f#���t�N*_7r�d��)Qy~H|�Ù� ex�}O���$;�r,�)�1��4��CxJ-��H!�����t��o�E�"�==X�� ��ޘ`�_���86�>��Ǿ��Fv�h,����s�DMkVس��f��)��2�g��o��ڢ��B2��%�	L7��4E(^f����+��Y悅�K;4�D�ّ�8m�˳���>7��0#�ih�%��-b�����}�5́и��r�	$^�X[��
E����a����*�u^�c7]W��z0�J]�[�/�Lq�Ž�xT��6m�΍�Q��knJ��V̸L-�f`�����[�],03�C�ǏF���C��HVr0JEv�:������(3�]��W����G��,�����? F7���t���R>���k�m�Z��oF��	`���`�v�3����p�)�j/t���I]-��3��t��������x0�f��=�ݚI0-4�g�j	-.g�Ŵϟ�������qk�m�:���l�A
�� �\wz�R/���j�0�CiH�!�#j�G.N�_�&����%+��m�- ��-�>�pB=1+i���B�CM���dTto`Š3��&�[���[�j��" ����Og@�ck[�W���=��XD��
�g�U��m�m�� P��D4
r�f�2����z��L=Ġz�r�v����#	���\����}5zs�h\<��2 �\�$o�ͣ������e)�~5u��K@O�j2��q�Y*��o#�Y9| ����px��瘆(�n|��Z5F,�e�ly��*�q���kB6!S5�je[�;�d�n�e������?�}l�<��ΈE���T��GE񊸡��Y�*�1'�+M�Zh#�T1F��z�G�TˆnKp^��J����E�\�{eg��fi���PzA�Y�cN���Q�/?�㷳��w�"����6]��5�WA�}��{����&-D:nۿ#OF��jZ��f��p���}��)q�z�#��Ed_�j�]V<.�]�D[4}vr.t���B\��<���g��qV��%6}�,;�5QZ���l>��^Hݣp_��,`X *\������/��]CaBf�!�R���_��.f����Z�W/
�z ��%3m�V��P�y��<�y�V��3��d����Sx�}GJ��b����bL���a�Es�^�,�����	�����v���lf��;l���.�g1S{ (^>��@�e��en�mr��t�]��f��Ӡ��_*2�3�-1�5R��}p1:���l���[<u��a�E�L�hA���]o?�uKq�n@��W�M�P�)�"OV]'�B����MxO���k�����٘��@~8X�E��}����U�"��I)�*ڽ�3ʔ�v��Ǽ<Gu]����v����맠�o�����ZW!Z^�>W�[#;J�^6_22���p����[�ՠ&&�~CՓ_��3��:�v�J&�y�	(4T"|��4�3���`mU��]�+'7�Fſ���Li��pQ�7�tE�d�A\y
[�����('�|��.����+��]�*-�B�'�`%�M%��T�|�+���ņ��Cd���@�䁇Qv��x�<�򶲱R+��=�VJ9��C��)���5��r�-aaQ�3T{R���Y[f� ���^��d�N=��}�=��vh|`BϠ�>�?c}߰�%}	��=��ح���gw9 {ڬ��<%n,�!Ӂ��p�S��╬��TN� �q�G��h:,�v��U�_����q���;�!��F�,���u`�-ix���~�h�/3��/'1�T���1���;A�G�HIg�T���J����Tm�a綠n�Ȋ(tx���Dv�Ul�;Q� ����2��q�$�H��An8v#,ܦm��%�
@	�a�/�[�b���<f�)�v�
#2�N����%��@x�ƾ4w��<L�Z!^SVn�����p���(Z�
X��ܢ҇l�+����r��i;����4���&Yy Ԥ���=b*7�i�F�8j+���Z��ݎ�hS!S��dNw�8��?Жx�?۳��S3%��RPwʹ,��R���s�� om����j�M���˨��Q�5k�|��:k'aҘI}7l�+��$��g�2l�W[�(��TAp���t��h��nF~���Lr�+��׊�y�N�O�0R��,���B�/�<*;m\&M����.�M�q"�9]�x���<�����-Sa@��I�T����~vg'�8�0y�_q'��k�,Z�۽n��5�7��7��d����Hab�Tp��n�9��k�E0g�,��,�m��l�p�>(�F�T;���;+�9�s�ûi�[M�Wˮ�v�κ=��v��^�O���8�eb�%��]�Ȋĝ2�]L|�ʍC~5�z��2��#��Y���\H�cW薵Wן��_�T�k�uohZְ�H��nV�=����/�f;a�M?j���F�|����Y�owg��I�Ry�lR��+I�EsF�5�)lğ�*�.2bd���zh�tB��3�a��������c�1W%������ c���g�*!��(5`
��99���pBr��?U����W&���q�=��Cz�PK���һ2�ǃ�e|��@��f�=�ly]��L�װ��`��W���]�>�
��bgL�	"�#�3���X�37{����� �bj��s�ꞌ�U��A�� yn��"ѹ�����0Ñ�Q9���a�0z���� ̙��|4����u�XO�֟����E�ύxb�9�0m
vzX������V�?�� �L5q�������*E6J�W��,k����,�������G�R+�*#���1����P��K4~��g������I����A�EA�7&�7��{��d�S�)��~������#��<	f����,p6J,G��=�/;"�P*C�BU2_j�GNrCe����r�d7*E���l<!R4u��-����QǷ͋��qX�|^���O@�r���'aG���pb,��swrO-����"80��W(����4�f	��f�E�K-sSM)���̷��"�>����N�?�}��4��cy�1ʏ��TT7�~�܁.����3����0p�t�����\����17�Ea�Y�W�֑����&7�4�+�种ȉ�y�-?��K�VΟ]�x��f_/ m�Pg�q���v$��ME�A���K�5BJ��k�L����9��Hy�����j}�u�ߎEK@6��Ljl�7���8���둰)�����#�>'���	����?E6	�(7�M�������ל0>��}�~;�R�Ł�g.hA�󰇕.��w}��d�]o8��
<EM<k/���T���ܫ���-	ʺ��B�Q�&#���|&]}�~�I0�3�o��Q��U��G�%ɵ�$�o�z7�Ρ6q�w�SoGJ�}p�0�~1#X0�*�1��Y\��~c��or�V�ɦ���_��P�����w\R�m���7�����������,�2�b
��`��\�N;�/�5���!qC�O;���#Ua�N�wؔ�Has(�d����wx�aF�V6:A�����M��٤L���P��(�X�E�wU���Cx��P+��a+]+v5�V>�Qo!L���ȀbY_�W� �%��2L���<O�ᗆgwANj��q=]��9�a��d�U��0Y�T�ˠ`v�����D�X�8�`s.�V�,��I�Yp��yh5����9�����(�a�J�A��qg�h�}n6��C��ɇ�H�`�V�I.��>,�	s3K�:Qm�Yg�!-7@���?�v�YLťհ��&�k�ZÜ�p�$�����L6��z��<
c\X���,���O�n��ѵ�ڛ���0T�+�T�`}���{a�R'�ꬶYTL�R�������m�@�S� 0���B� ���-�9y\s9Ԯ_��Y�J9C��n�|����=�ckI�p`,�,��規G�j�.q��:�[츼���L2�[!���4<o.K%s����#�Ç|������!Y.����N1����7ȡ�vUp��03NT�Q�A��,]�o�.��g7����$���=�Ԙ�=�n��긞����}�մ�v�=��������
��1�x!��I��m�;�.�Y�љ�' �'!�9oỢ{P��t�/.U?Ѿ@սW�_ЙN���d��V�&���}n��G4��pT��4��i�� #��6�	�q����U�i�����
\:�0#�(��\��V�.�w�?�X����3ԭ�?"H�Z�76ة�>r�����9G��=�5�'5u�̉j�Y_8�}f�J�`hzV�su0������b��j+O�mȔ�ַ��)Z$f��s�dL�-�Lo�jd���x�.�ܺC��U�k�1��=��I9>ʱ\ސ;���'kuI�,͑�}��	+�fC������$�v�2u & ���R��P YL;V���{�c�3�3~.sg��z-���-�J�gx�� �Q$(�B,����$sŬ)��$�1���9�|uqD[GCM�~D��y������7.��9�3��Ʊn-��םS���y���j�LtY?����{~'t\K���v�D�8j�Hz�3ȏ��<�&�l��;N� �Б,E�H'�{�[K�@=��k�k�?����K������U�r��3�oɕB�{�k��>�n%]�Q�{����Ź�Q⯚�{���q�ڏ��kːB����94�'_��Zѵ@<����L��W�i遠�(-���'{������X!���U��a���;
7��N���S��߃��g��K���<�3A��B�o���c���:FF��n���ĕ��3٦�-Ȣ�5�C^�	����;+"F.,�r����7�_��� ��ɣ>��ur�3id��aE�R{�{@�t<�^m�E;)�`b�ӂj����y�f���[`x��2���e�N5إƻ>�7a]���6�Z�������6Ŭ��E������ ۃgRm? ����񱹗����zHqQ!�Uắ�r�S�?��=��`��L�W���a�$����ϳ`Ќ��8�}Lh7\n��kw�C����������⃷��m����B���ֶ���͎{�ɚ���mnU��`�_LU9��I`MQ3���x�O�������R]�����.���GB�QM���e�&�a�M�P2os���-Mm�7���-�����#A��H����:��J���R,�T�9K)P��n;�J@�=b� \m,+�@8�f�G,@�AZ���(���h��V��M��"w�r�qW�e��&<���c����i7����0���cS2]3@I¥p6� c�bb�Q��*u`� ��)գ�K-�s�p����g��5����:����F�﷮�.X�� ���%!����׵9�]�spn�'��G��6��\ʩ�do������J	��!j�Nҵ�	`�?iY���������zP`ڨ��LJ� ���@��?QÍʛR��q�DJ�/��{qM�d|H4kS��e�ӭ���6P�? ��豕��Y���!⿄+���_�����3�A&��`6��,@���@���!r˕��bDJ�n�ݧp���.�4J>r۶����j�2l9	�ў��!������	�L���HcF�q�TL��t�^u��s��*.y�`v��3!�nS��6�!$x2ͱ̢���*d۵3	�ы-?�d�JA�H�����a�a�^����Z.A��6�>�A���gc�/.!�4%YPϕu�*�S���pC_k�\���%����gڑ{v���6da��m�����c�v#�g����6�͌�-�צhkǑj`s��a�tm{c�6�w��K�$��mPS뀵zY��F:jn��6SصIiP�u�IΆ>�45j-XV��w��%���Gp��(k3  ��/2�_�"��d�M��+���n:�Ւ�X�ٳ� ��N��L"z�x�u;��Hj��/�z{^5_��auR���l�Ɏ���qK��D��1?]�u�;V��?�w}��O�C��~�f��L�y�����==� �hCv)��~��U�����[YR��aV�^��&�q���!Y�!���6DH�s�5���̧b6�ܬ�>%Q�<�D���Ф�H�~EH�g.ٲ�!0k���p�Y�}f�������8�(����� ~�j7�ܹ��/�v&�T�ƻ4�����"/�����=�O9S��kc���:y(��B�w���� >������$&�{�(e�K���7�<�)����#�y=����k}��# e��C;��/J�� {�U^�����#��}�z��&����0�4��1�5�n��uy�� �e��d�L������_+�BF�x��_�x�C��+�#Ohs���Z�H��w�~��M���
�d�W�o�u���M$B��K��Gb�u� �����v�B	s7��3e,�m7����ʱe�j|��}�]�� �30���%�tm�`r���>���w����oQh�c���Q����&�,}:�.T�ڷe��MS�C-8��yZīz�F��&njh��-�.���[�c\��Z!/x�D#�R���|�"�$����m�b�h!�I1X�c�"�@Jȸ�q�f0[y{I���I^pO���&T�3A��N�>9���O*����}�SZ��jM��{x4�)N<;k2u!�[���W����y��+�UK�s
� G_����|�q�g������ǟ���G,�ոS��F����D�&d�^+Z��ʝ�^����h��\�sl��Km���wa��ݚq^����� ��@�Y���d��v�~B�U�_���}�0�T�f��|Â�	[f�g�W��v�2XU
�fƍVZ�c7�Et��ix`�`��8=�t�sQ�4�\���۾��G�`{�
�W�!=�G���l�����0ݎ[3~�8�<f�b�[�p>�R�G>XmbnS�d�+��A�w��
��B.�c\wQagE`U�de5�<7y�58�x�?q\f/\̖�\��GB�2P�+(�=�S�ָQ��~7�M"�+��1{�:tNL05ze�_q�Vl�����eLܘĔ$e�;�F�
=ϦtրNZTpG�5Qty�ya)}-8�2k��reJiP�h{7S`x!cP@mz"���#B3Wn�!�l�Y79���&e&gSl����0t���*۩���5���-][�}n�����#�\��G��f���}�lK_ЌP�cP��g.��D�6񣏪�dfu52g����ni�����4)�j
?y��,K�O<8xl���;1Єd�Dα�Mp�? �QX�[�I=�rI�-6O�w�Fv2�Io�$�1F/��C�l��n��~��0�n�h3�ڝq�[ǧ��t$�!;���P������!
ZUU3gT�r���@��u�z�B|��e��\.I�y�p�Q��O�bM��VO��p�|�%���!"���uŽ��OGl�'~yOd��}bF��X��/�
?,8���
�j�Hpޱ��S���u���)�@G2���ku�ŭIj�Xn>j� �7l��`�:d��T�T*��c�2����<�m��D��Z�Z���C\��z��'p�:����ζ#�2���3̿N�)�����SK�zJq�s>ڥ�J�ۏ�˚YE/�{!t�r�!�����.`O��2��S�v���(ZÉ��GS�� (��;�%���󏞂�V,�����}�<z2Nf�fs�ux���ؒ)����ȸT}���U�F<���|�T#��XRF2c|��=��*���V���i^��9Oq�6�-k���Q�b�%$I��@#m��u��Q���'2ۿ�12Ò��Q�L����^v�w�h��5Z,���cc��uX�-z��z�]���	qz��{NDR���l�;�����=�HA��L�<�+��������(�]�QN���nJ��QIգ�~�$��G�������=	q��N�:C����Pq�_aM���87����%��4�cx�k�9���%��7������W�|$�g�k.{FG�'���6�d��CfW�$���4��h�Č��i:"������&��4F�W�0�hĶ�P��WX�r��S��D�۝�β��"��zH���@W{�b&�	�HĐ�N'8o	�Р�	O��<�^�tQ79dYe�4p��Y~�'x1�!ж�RK��PO��+���֒���+7Fk��q��T�T�ȗ�����V=0����(�|���uE�25-�^|U����(S.���z:��Ԝ6���:%���.e Q}}"ﭔtJ(�7��V�W�od����֗c�ڲJ�X�D�!��U�g��B��lU[Hʌ�ԑ�~B`�`H�5K+!~���o����@�-�Y��Ħ[�L��\�_;�V�'�2@�6������i�������g$��
�tZ�0I-�
��*�~O4k���4��:���<s;�p�[\�Wn�U�.ئzct�ux�៦q�B��;օ`��]����m�EK�8м9 ^.�c����Brr�$�J����z�z&����4j�(P֌rR��.��.��f��E����#"h�?�a�`���y��3�%M�	��^0X7�,��8�d#�W:>2��<
@�k�m��5� �R�4E����hD�#�c
�йy-�D(0�Z�,MG��;�-J�j��?8�e�Jy�q��Z�Q��q�G��$��Kp��]��2���Ht�ٌgu��ػg\�Y�~�E��͓�Xӕ\C+}��^� ��i�7:)�;t�O�Lw(iz۪�A��@�������Ѳ�]ՅT�n!kB�M*��w�t� ��ͅg�~��(.��M+y<�'sא5���?��Z6x�Ѯ�<K鷈` �±�u��y�ܰ=�x��_>�I̗[�M���=�I��{:o�>-��b�8���b�UdI��a>�u�G&nݝ]{�Ѻ�L�tB�U͂�6����Pg=ئ7�pغ���A�XE�x��1@*XCX3��64�.<i�<Ǻg�F�:9eؚ��kR��ng��b���!e)���0#Ԧ1?��T�9V�p���7�3�
/l����Җ�#J ��<Lz��L���B"p��h�5k/�|kֻsl)wǗ����9i3���B�iiC	���󐑩N�9�qI
��4���;Z)������f���m˂�� k= ��|Q�h��_��k��c�y3Iw��s�*�~��$1���m΅=b�I�� g��F���������a��i���QM+�A2�E3W����S��h?
����{H'�_�j56�0哅��-�c��0�o���1��(:��pl���6�����X!�����I�T���)K�å[I|�~NMU>��q����~��HaR���z#T�b�V-�B7����=��Yv" ������b��{���;�N8�����@-�|��Y��n/"���ʶf���n@�D��R�`Lq5�C��ja��k`���[�+d^��´"�|�'4̽qG��F�M���	����IH��j�Ǫ�(�m
5e�<6s���k>�r�z����].�ا9�����U��o�t�9^o��W�7����`�e0))��a��&ӊ�"<9�S��+2C��ѡ�f �`$����˪�]�F{p�I�U���:l���pQ���qY}�s�؋�x��W-c�H;�Þ������/���q~�vp�n���̻E�3 e|���>(3?�<��������D|��h�.˂=f�i�I�HK�\O�P�GB���y�� �w@��ӓ�8�����?�N�������,�٨��"\��%��"Z�wǲ�bi�s.��=������7B�����}y�f�d�����9��h���r��I�|�� ������NZ�5�����NA�L5X,��	 Z�^�x7D� ����t�	jH�(�b9�}��A�  ��ՊP����4D���X)ڱ����e)�ɲȈ�a�l-�l���-A^v���g�#�Soû��\�} +^av%R��]��m&߈�K���{��<Aytyq��i�gْ\?C2��
�[�1[7�p�潯l;������Z:|��#�e�ib5+[6/������h�昒Kp�ك���A������@��"��_�s��>s/1�ۂ#���Ұ�B��I�� C�$� ��A�����V�
�����R�@"�͙�
��|���l-[��n?�~9�S�T���AkȄ��+ vok���Q{`\N��I����p�B~��� ������[J5_1�=hXW���M_a��?��9GA5����cU]̸��e�Ң�>���b+jK|�?/b�[5�ٕ�zf�K��v����L-٧�`�-��MV�8��֮,�W�������9�sdyX��Β�{�%��@4�1����R���M%MT#&���84lcN|����w�yI�z��s xUco��<�)n ��+�Sg�J�w|-,���W����pl+����0�b�%f�ރ9O�"ϊ�����! `��ٱ���׊�Ζ-/#��$�0#������Y�Jٶ�⋻��A��]�rBecB�承�$��~G��^	iO@�����6�	E*~魏�/��Y�OVݽ<mԁ֛��,�����,\Θ��\2��5�����<�W�� 	��/c(�|5QGsP���[&/�lC��;��!N���v%�ǬhBI,a2[�������R��NcH1L1�J�c�l��N%trt�b@�q?IV� 2[�����7���cꐐ][$b��S0�f1��g7��~'��;�:�0 ����YS>�xm}��_�a��'���-��HPo�.�d�p;N©N;������t2�\�V�%�?3��g����<��8�u�I��]��O��f��u5�=��j7 Yn�zb-$<Oy2	C:��[�9�[N�wp�4�C�3��J�8ad��m���Ƕ6��\w�3�j,���Z.Y Q���h� 	k?������a���u��U-�:9�1R�T�0�s�h��%�p�/��P�{l�h�������l�m�GU*s���ك>�~:]������ȳW˺0���� �����t�I�?2���C�[$X�c��^w�ND��jE�����]i)e�_Z�z�q������f:>�i�ᗐV�HQ"X��Y�l���u��Ök��w��Ы�S3��-�������Vj.g�8�ܼi��G?��cS6���5��3�.A�Iz���bo�X5�G��=����Q֖�e�~��/φp!q�b�a�H�[�%5�Ij����S��ʑ�.Y��Q"������y�'���)=��Q�¡���!mX?���[7b�Ƥ�ě)��<R���%��B֜Q^;E���]���(Ti��� � U.�D�� M�.�
'�@Xg�M~f�L��j�`Yd52E�^k�:���^���ɇ+�q��IPڟ:����xƹ���I͢ �e�@�Um��:闵e/� �l���l��|V�{X��K��r���t:�W0��R&�
^bεo!&+��;_�m!�xj#��	���wH�UL�W��2�V�Þ-��q�y5]��9��n�^b���A�x�[]Pk춢G����4_קּ��
����1+�E�� 	�;�I}?a	k����Z؁H�9��*��r0�d'z^z!�D�����&"׀��#ڤ�2lPo�mBג^�6����O��,X�=��J�ij��^3�����yK��ƙ҉6��7u�L�d��0{b�՝>奝=�.�����MH>$��L꼆����~���D�'�pn9c�!�Nb�J��lJr�+�;��m�ʖ]mXmcԴ��ҁ�Ȍ�N��!��� ִI0D�Z��J-���Vw�k:Y�L,��"z[ԇ����ѿ^�n�$&��4�ܯq�@�(e���e 䪿ggU�V�ZW�_$�[~����u����iy!�æ��9a�w���߁0���~;�UT�Z��
�,jKW� �A���2��3�g��&��^�Q�`A"LD[\�Z��ß�(�K*hA�OJ�
F��w5��f/�N�§vd`�pz�4o��/�Duک$Ŵ@����_�[O_�5J˪�'�>�ІM�V���.�}Ӿ�Ao�b��M��Y��ߏD+���q������2K����67t�E��	B���M"��@q9��&\>y�7;+�8��k���\KZ_��j`���)���(or����'�j$x?��=�� *�My��n@�����r]^(L�&9a=n��\܎j�Z�uMh�>�8��U��`���WH7N�BJ�����Cn�:�Q�j��i�s�xf�ic��c��(��71_^r�PpH��)����U��RH�t�1���������p�V���7�<9�x8�����1��d�s-���~1�?�A�dTa��2Bv �J����aڐ����G�W��`,y ��v��l�>_4��
�rS�p�tH��1�<�n&y�,���{?�K,Mt��I�;�����;.Z{�������&e�i�L{v��SV�W��wJ���	f��0456P�Mz��zT�C��ǁ�o��AC�:%c���ihy�⳼U��A���=��vW�y��<_���h^>���3ڇd���k��z���m��P�;d:v�����V̀�j���8�!��3L����s��u�NK=�:iG�����]v$hTpdK�'c�1������hW��9e�&��f���A�-��� l�����	 ��6�mtd^3�[��P"�o�M��j
��Q[�q���ج���`���lToGLXG��^�c�_��d��J�&�Z�=�m�@�fм=	���~aSp��=�C�>�J���-5��L0zp�����Ҧ��SF��4�e�/kQ�Ć��"0�h%�jxå�L[�!�5��|T�w��3،�X5#���O�#��ϟG%��cV �o�^[19Q*���;����s�������|�%?|�~��{��E-t�
�>,��Z���9�5��"�8-��j��:!�̼����I���ؠKe�9�������yK�T�����W��U-�5)�K���9��������M��7�_w�Vpa"rL1��eNtc3UZ]�y*�3ɝ?!��^K�m�ƀc��W$�xՁ��^�l-��f�>.�zu����$
K����~O�O�ZMJ&9���<��,���������U�d ��l��{�ɉpZn����/�X��c��`k�*���|�ϲ�~�.��N��9���>;��jƻZ6���8�p	j��c��8om!���s�����xpT�|�I�Fݫ�w�L��$��)�S����w���s�E��#kɥ�9���IL�`�2��s
M7�8M��7�L �:d!��L�X��0�<�q�?��n%�U]���E�P�3}�I�A�x��R�6W%T�M4�\�2�2;r�tWN�K����c;wB�`�]a����]��E͋��x(����<�/�H��d��b7�/Nj�f-��J�ʖoA���� r���۰W�I�9�(3���Wą�Rx�3�P+��4��X	���r���z{_�] ���6<RM�>ں��T!U���~!@�.�S�l\�BѦ�G���w�&j�FH�~�������q��Hy�s3��'|
]S]����)Q, �z�u1� �jV����e���Z*7�&��v��[�@�o�A��]��5U�O��[F�.�?.&�pv�z���u��^i�ۗH�Dz��+�&gDޯޚ Y~����`YE��k��8{5a|C���j�Jpz�HYۏ��@�^���ǽ[��d?E�/к-k�S���ۑm�"kc�'%�ܮ��F��
H���y�`�����,6���'ew�DW��}A��m��-�N���`%����^{�U�.���vn[Q���LɥtwE)R��96cW�A��%��,�e1+�5��gd6��Y��+��>�|�i��LIμ�DpY�[�)���cu�� O<Ȁ��J/�@���*7 ��v�.�̾n4��;��PP�%����tlgڽ�A�x�O�G��<�����҇�àN�P���_�5307�B��2�}t1_@c/��8_pE�ص���pzbL]vd+�8.�~�뮎R�>)�:������4��_�I�i0(��4
�IoY���2?\.|�:_N�I�г�Xb�����~�}쒊��>ɚ�Ar/B��SF�6@U�@K?�r~S��ͣb�E��K�0��y-����I�ynClQJ��f\MR ��csҁX�b������tu_����]㣚�
�S&�)F��ْ�����ʰ!���#v����~L�}�U5/�N��v���D���1�6�u�|�.��c��`��Utb�iy�^6����y���~25�ق|Dx#�3��Ý]��T�yU鯊ƿ�sd��L�����$�Qi���X~g��,m�}4�:�E����o:��q������s٭>	yZi��13�<`f�;#�^��عB
�2�<�{Fқ��E�L��X����p��oGhn�6J	�iҞɅ�}���n���Yq�� �V̇h�"|�7�eA�^1���.���afH�L��-,M��?����}-h�?{���ܑ6`3����ny��T�b���E�`z�1�41�_�S1U]{��PQ�8�0j��K��o��ˏj5}(``*@�k��Ļ��6�m�T��.y�kp/���.=�p�h�@e*�Z�����`���AZѹt�"r�9�/P���C�O�3Q�7ȝ_"@6=�[�鿞23��V���K�Cw\�R �h��j��9F��Sx�:������X44��bf�tR`�I�4Mv�w�At
h����'ů�<|ʡv��!&�}���= ⃓�n��1���Z����r����R���Mx�y;��SΉj9Q��,y�BU`n�,�h�I�*��B���˙?��UKǡ��ڏ(��eLsV����U2M�ġ���w;�*Y?9w�L��ܓ,���ӱj_z�E�O��y���� +�(\ 6�e@m���?�.-��H�"���.����w&�x�4�$ݞ��%�g�����@_`�Muc��"�e��u��xON��0o:�G��	k�^��0�����l]Xy`����K=���i�c|Q��f��,���ۼ��}�ʔ\_t��j�7��?N�֋.Q6͹�89��!ii5]���"��c�"#Svm��Aq����ڍ�Bi�ݛ�-*i�c��%�nU�Xe�ABV!n�H\!�qR`|t/z�5)�O`+ѝ�n(������� ��lP���h�c[>��B� >$�!�ۥ�eIح54�6��u����HDr�>d$�#�L�����qF].i�u�+N�G�A{+M $v0�\�d����<�Z�ti��Jjq��Z����娍B\�p#7�/������j�n1Ҁ��e���h�9C˜��T�)]��<�
���:���lQ�2�ay�L�{����D�\�ރ���R�Ao�d�I��/��]A�aJ5�/*�@"32 ��������c�[�A}���߹�����t�<�:%��Wc"��>�;	���iT��'O<y����e����Nt���TƖi
�%����ሦ3��bZ�Wރ�-���9h�%|8̑��G��,��9�O��Zs4��'܎,���2��b{P�~�ˊ��m�"��F����A�Oȿ	oׁ�wc�a�	�؝�f�Nt���
ʰ�1ΚO$���18���_Ϝ�&ᛕI��Юw���l�W�m�c|����Y_P[eB�a���P� d��.�Q1����]�=��M0��|=�i���K�u�u~��Ъ"H
�R�dB��~)e�~��wm.���(��၎��_������qHa�%�4����O:*�4˟T����TY����ܧP�J�s�*�
\����Ɍ,��
��|�x���.8-L �li�_�r��[�Ɣאts��A6X��#�%��~�5�2
�
��� ���0b��ب9��*���A�1NW���Ȱ�ƸT���󞻣o܅G>�$[��M*�H����7�w���:H�����N����J��5C��4G7�{�ô���mF�A#���
Z��֮��2:u�"���2���[e��w�O��֊�W�=��T���͞B�JWI�d�j�$�
4#�:h`7h�R��w��4��ZJ�sj��W����iF*#p�,��f�na�q{��Yy�����g���Xk(W�Fӿ�b�ҍ�����@�IK�������^[���S�UT&�v)��2:q��w[�g��r�L�=�Z+�1�b�ˤI+�-�Յ��w�N�ՓHZ����Rroh����˜��Z�ֆp`Z����@��괝������Uu��3��/�F�=<�A���9�~����(��Q�M/�n���	�?����&W��v�c���R��!D���k���;jF%����"�ٟ�ȸY��w�&��~L��"/��G�Z�x&R(�e�:�3��3�d&�H�]�d�|�/��	J|/��D���|�r�/��A4WVtP���^�ي�"���q�A���Z1b׻=g���dHr[���b_-s�JVq�î�Pt"��^��<�`f���'mNa2�G�v������������C
�Aޒ~��d|�w�Y��e��|��7/��3�٣		BK�A�Y��hz�!փ7�z��SZ&0��{#5����nH<�m�К�7�Lo�}(\�c��/�C�9H�BqP����H엡���p��K���#
Q�j��5L��O��ە�ҧ��(P�|	p{���F�����F-�Cr�ȶ�9p�xvqnPz�'���ڬ
d��t@��e~j2?�Dõ��
�RF	Qtʿ^օ�¬?[�>���hɹ�#����*�V,�V���kn4�K/o�1�fj��o/N"�=��!�L����'<�:$�	S����x�MƁ4(��|5"6�S��i��a���=��E�6`5����,\�JHl�>�P�"q)�=ϴg�I��K?9�l`1'(sE_��
����d�X����8X���?	~���I��I�<v^
��L���j����WT����'�(�a Sv?/�V�[:�Sx��૖�3�E1�\���O�mlb�k��*�����6���7�ϼ>�{(�X��9˨:��QEw�]��~R��֠]o�u�-]!,i߁�Fs"}@��c���f2����b�cOQ�WȒ����&"aLݞ���a���L�F~B����$�����1���K��l,�jx��bL�5�I��a�`��n;�����~i�U��x$��ʱ�~�?=t�7��� �?�Q�?;���qCaN��.�: �p�)Ϙ�Y�Ȧϴ�ͻ����Z&�[�ٰ�|������{��Pd#���k�ԮA�Sf���Ht�o��%d�D�t�� ��Z���c����M����J,4+a_��6�mA��l�Ufu;�X/ݹ^7T���3��^��\�����D�{ ����׈L��£6����{�ȑ�FV<1
�n��̯2c �jF+<l�u��6q�o���Iã&��O�	�\Փ��j��J��؂�1Fyߥ����:6?X��b?��6� ���pՌey-;������`Z@!U���Y���X���d�腗��"�9-�{3�5n	���`T>~��|��Ru�_/k2;%��`P�⹫��� � f����+�NV�2�gj+s�S 	NP��Y��ٰ��m Zw�$�ˈ��lq5!��m.�
Up��2U�V9���,T��|����ҁL�������r)!���7����/e���O������g�!|ɽ�L����6yNJ���^M�o����Ji\H���:��a���
%8�)V����\d�\�J�e��)��7E ۪��������K��\�%�m�q`u�%��U��q��a����Dmȕ�5����aN%�@��(�n*Ҫ6��uV	ޑ�鸺;��X�Ĳ�+���u�G�`Y=��h_��O>��E"њ�yp������5�X�o���p��,f�����@~��w��4��,9�a-��7 �\MV.'�Htm��|�.����Z*�o�-�br(d��m]��ӝ95�V?�%ډ+���@��C]�#.���i����؇���G�j@鞨���Z�H.\�#ϗ|�o��餗AX(�,&?4a^?=���/Ǳ�ٖU��9D·�b'fj�GQ��O� ��R���yP���nQ�U�=��STʈ9�W��L��si�N+��O�O�%�Pz�O� &z�E#���ra��ՍLч��{�������6��ϔ4��R��!LA0ߏ� ��p��K6*�/gtrT�%90#2o�S��C��Z>���_^�"7�귭5�!����#,�'!Rҙ�O3�q#�Y�D}pO�XnsP۵��8�0�X��<���"Yݖ8@b֊j$%wO�ǥ�l�-<ˉ8������7�"bMy��-��1P9ux�H��y�{$�_��d���%�P7[1�-���LR��2��0:K�%�sJ1N�Y�hp;��K�a���I�;2/��g�3� �n��D�43־G5Y���
&:==�	y��O���/֑3z8�n]㮰 4�La!���4�K�G���-����3kX�uJ��p�7�X4\t�J����P�M�Gi������0I���Lak'��E���a�R�;'�z�k�����js|NC��u���?-7!&T`Tg��Ӱ3�Hnnd�ܦ�P�x�"��z��x��v&�����Jf(?ET���6��ވ�-��R�f��#��H�\�ɡ[��9�>.�*F���5g'*8���z�&�K���)�ζ�́b5L��:�O��;�;#U�n'�G�|#M����
�怓!�8�;q?�s���Sa󹇸;���Dp.����!��4|���+zl̍�*�����{N���<�2�Y�؈��Nn\n6��w�璬���V����OOF�I	�j�L:f�+l7�i�q�����V�@ۑa@v6x��=�/nkQ���$a�����S�S��@ ��stcaf���Cd�[c�;ŗ�gf�?I��)���T��W�ڈ�؍S}I�����1�E	�:.��/��[�����2��[a���Ar���B�B��ɑ�U�������ʱ���Љ�v���Q�OJ`kt���k^��MF�W�B\:���Cn�s3X)�C��`	jw\n�u����`ڠ��(��*�O5����\SFu�/6in��B�hE3_5����MB�:��s�X���E#h�9F"�q��X����K��E.�5��6�G_�Q�U�.�h��u�����BS�9��-nҞq]��=�����`/�[%O��wc^Q��d�,��z"(Y�'G9�]���Y8᳧ܲF^��+0&-ȶ6�|���z�맘@Ә�.��/���zß%y���������+�)�f�})���w�����|�Q8j����C�2U%�I�
d�-M��A<��ϱ��X{�jb�1zj�r��*��rn�C?�lܺ�A	�Zu$������q�=G��l�V��Ǿ��9�nC��znĆC�h����hk�a9�ǳ�!$��]�aM��W�a�g҉o�℧�M��/�a~M�K����~#Bda&:����</���$T��#P�P��b���b��j�m����{}KNá�Oeĉ�Y�>���O�&Q�"�����Y�F!BA��=�L�}&�`�vHM�D�s��o� X�l���9,�i�Ƹ���x���t_����9o��.��׃�4.v�g��1u�^�AA���2_�C|0l٨�[<sᩄ��z�'�FL�������<���E�9�l|�L>������K�(���g >�J�� 1�ő�q��P�ݚ���W��d?���BDsۣz�6�	%ٍ�M��~h��;_^9��jXc�/�A뻈>�O����1~+��mq��)y�6�lw�^r�0��d�-gW{���GHT��(���%SJj�3a�Qi�"D�	����I��$���$���ұ:1¬k�˃� ��n߳e�p�f�|�۲�%j"?v�q����r�;�VN����L�~i%�����	}��Ճ�V�u��)��vB�H_�)��������s*����O�n�?pA~K��6�&�`x����X;e��j.3Z��d�_饮O;ְG�,zR(����2KT��O��v{�a�8 �O(�QL� 1 �e��4"9�H=ն�N�ꌎ;�k�n�*md�v��#�AR��@�MD#���:�Q�t��9<6�k���)w88g�R"ȁ8���Wϐb4�{��������
�ҩI��'�S��s "Z�5��ㄶ�y%�fi��a�n�KM���O�Y�4a(��Zy�k�6�[��J(�>���<c�����ϙ��D:c�c� ��+�M6eF�=-�2��J5tR�4�G�?%kK����|��"�Oy�_2�~��Z�r��u���Y@�L�[%N��j�L�5��U���H��K6�T�lw�������$�K�_�/.�� P�Z�i⦓ɫ
����,�}�̈r8���|H� PӜ^�h�5�k�.���[��._H}?���漎4&�JL$�����ƴu$S�DأOu��r�#������LԲCkߗ�g���'$4�/g����֭(Jbء*������?���9|/�T$�	aR�S�#�p�Wo�:�0;��ޞ���k�����Æ�"'e�+�3G#�n�g�����m���s���U�"�% ��t��;�=kUE�z&k%��0�)����xr��uBd�ĐK��=�����)J��Ѽo�?��'�Ni;#>��K�ZA����*�ZS���[��������"�O92�r���YU��R2
1��."f�[�s�I)�T���lR�Ǟ.�`j��.Hg_W�*�B�{J����iT�P�N߯�{�� ��)��`�
O�ȣ`96OD�����uhMt����n��jh"�<������)e��-78��nֹg��d ����ӴN���5�AZ���Y����6>$}à�,���f��:7q@�=ϋ��l�����c�߰�Yq@���Zd����i��`�1�Ʊ"����:I,xhc��K�^t�*�]���CM�yV%�;��}��W�E-�y"�&�ؔg���%�
Y�~��wk����K�*���C1b��S��yvd�=�&G���w�aǠ���M�d��d��,��*�!m�
TGl��_]�P m ��d0�$��W_�����/0�4/`��7�C�T���L�%�2��J�M�Wy��*qiri�ڳ�N��oQ9�@��Hxν���T33��^"�s��݇���� S^?h�W �B_�n�/�hH��}x�g���r�J����kH�=n�a���9�`ݩYJ���.�ƶ��#+9ZL-��$��9i�؂�� q��l����t,7�|�����/�k���skb�&y���ˉ��$%���e&M��l x/��ڸ\iI(o,!(�{3����#m9��~��U���A���j����̲��I*V�h>�"�����G�~�/�+L-Ҵ.1T^
�
��Cj-��B:<��%����Z��4�a����+f|�a���mW��&Ⱦsx�a�SiAV?A�����'�&t	�Ý�bE�	s�	u0d��t��բ�~�5:����Xjˊ7ar�R�b1�i乼R����r�)��ǬO�&]h<" �⣋���z�����l(�):�}�m_)�&rƘS}�-'����t�+�ڄ�1
�4TzJcA��{���]$i�W�uh���B�����We����2�j�*�3�V�����A�ӟ}5ߍ��K3�g֭�\E=T��0�rX�C��"@�`�x�5�`�t`����H�/ӡ&"�){���MXkɍ�����u�i��֜]�$/����^��e��R�B���>�-��Nƥ�$:3^�h�yѰp��5P��|�n������yc���[	1l>��;m����%��,�('J�c�����؈��2� �27{J�)�߁�*6�Ù�|�HI�MD���T��'��?�?�����+.��Q^���(�)�>�/�.����M%�\�3"���ci�f�*��ѷ@&�aƉ�l�b���B�\/F3���,�]��ê�lF~�X=�v�Dt,�N(PJe�C�6�ӡ�6$���+i;s�Gr��FO�7?�����!af�;���F�"i �[1?���j�
��k�&�����>ieXr����<�I^�ĳ�T	��+iL�Tf��G��>~����A�DO��l������e}�$�!��k���J#q�3�������} ��K�>]�I�@�`��J���Q� �r�Dsw��<�oJ׃cZl���dTmN�7��M���/��ȵ�2
1��Ny�%-fGc��%�_�^����*՟ �-Oj"韚�;ܔ���.G��Y2��!�����iDk\���I���uN��P2&��`»��39]�<J�ۆ��{���q12���K\1���b2�2�8�;�_G�D�okݶ/�6T�����e�"Q�uV-@e@������	X5kԇ��cxX����#[�
��˵9����?O���n��)[L�t�}�I5�:;��1��Jz3��E�/�Zs��fG���p�nL����V�.�NwS+s8+����G�7�Q�<&0���6�̚U�9u	���s������y|�(�!fR�%OG�(��)����9�������	�j�� T�*�z��/�G�9L����ߙߦ�H �w�u+֩�O&�J�.�e���H���-��-�Vٗ�칼��p�=� �'hs�	��Lm,��Ƥ�B��٥��\�5W㢲���]2望�,?��@�ȅ�\�*T,k�(���q�h0���)�j�7ڠ�|H���Ą�(�����֮��aĜm�m�������,(�� �gfBCE$�,���ꙉg�'�N!�H�E�٤2�Z߼u��:V�M��������
^�^(+� �2���t9�,��OZ����E״��;&�v�D}��V���F%������c��8\L��Nڇ�3!�L���ݝI%�m^���%.�<�1g,�{HѪ��+�d<����J3��cM�ZjN'*
v������i�RIR8LZ��F�������h�|~����י�&��c4��
*Bha�����TKN�.,(�^G�f8�8���P<.p�7�ǦJLh���5��2�آ�E6�=�b�3b��w%d/h�3�[y-�Z�xFۋ�}9b�d�E�n;A#�L_�eϾRo�t";Ք}>sg]yjn�7
�Rd�+��Yp���⽎4q�VC�����w�N�߁F#�{Ɨƞ�&A�W�����c�i.O�W,H�*������	�{cO6U��)% �>E�ŀ1|2e4���r��=�Ǎ�2����'_Tr�=^�jg�ݸ�\�m�0b�D�]���Q
y�

m�뀘w�<)�krY<N�-r�J\o\8��8	��������	�y.ưz|8ȃ��6��
�1�6��D)aW�I���1���I!��1��C(ϳ�2�Z�a�����ȝ-*�U�pδ;�����9�u��Gd�41֢V�*�%1���j�L7F�%���q�k����u��7�;&#��1�V�J�@���0�=� ����/�����1%�E�)�l�+�+���з�����v�i�����TU�VM�g��y�M�u͔Xb*])��X%l!���WB��b ��?�"AG�B ����I�^�h� T�c��3����4KZ�b�?�б�V�h3��~\���'�[�.�����u4)M))���Pn��̱n��<^k�U��ENNs/����Ծ�Ɉ-�����_��&�1�i@� 0$8<%C֕��촏\���k+�V҅�SC^��C8�~^��b.�u�<��lb���d0�V�H��ز~�����wyC���*�k��Ts�c	d�n�C��x��YO�w����e�V��v�;#�3P�`�}$Dʹ
����6!�znȳ¿%�����.ovί�r�Ă>��b9bу}NN !�Aα�-�@ ��ǖ�H��c�J����Nq숭����������(��/����:p&j�bWz�9�KA�����nss��#�vV?���P�]a�Я�J'J8�7�ⶴ���8~	R���
g�4���)5�!�����S�eP9��tԮ��>�AK%�r8���9N4.
���/�����)������0�^��M�c3�䘧vYt;W�C�H`)��]\�k0VK3R��U��h�m" <D�M�z���5�č�fgT�?#Jeh#ŏ��^��/~ �9��:臡fnT�!�/��ΌCxUo�*h?�*�]}��n��߬W=˻H�\l���zg���#�-���xoa�\&���!��@*o6Ϙ���e����7��@��E�0�裾�S�9�p#�K�i�_��D�/vt��\C�U�F4� ����8��˷���V��M(y�)���l ��j��@�f�w�G͠�ie��B�50�z
� ���d�cz�h}X���e�!m	-K:��#�C���36��	���(��_5�8"u��#h��uv�#j��v�C20�DW��ގ3��,t�:NѠ� d'��z�e]_
�aG:��c���2������iE]UCO�E��ɱv����n@<�ܖ�컾�i*2���`�fz6M�s�L�����h�y��q���V��|��:s�u�s�����{�cbm���H��8n�<6�9�WAZ&�x��z+���3J�PM����ɽz�� W���
vU���PmY��É[�o?�����Qu3*P��xE�����v��DPC�s��.'4~��=�/�\'�����x\�����*��b��L��	�Y��#}�#4�m�Es[�(`Ԍd4<�	�3Âf�G�x��M|C$�mhئ���E�s���,L@�e��V
xF%�eS�C�l;�ն�W��Ƀ��h�����l�D]m��ojPʐ>�I�X�BI�M��t*�Fc�4c����z���9��e�n��]:�Ո멼G���`�����L�K����fT%6��/+�ۡ�Q�/z%�"��mC���w�G�s�_�>����N�(�.������L�R9j^�'���G;oN���a�ɇ}<F�M�&5W�Q�Yι�y0��C؅��Td���!6j�u�ve� ��3$���4��Ʌ t�~(�:А��XF��������,Ĩ$���0�H���y�=4�$���qyWp�w����b�ɶ�}c�zOЙM���"��l���F�x�@��u�$5�XOl������c%Uo�I�s!���c������!�pÐ(<l*�~��%�Yin+���~���&뚿��\�A�����LK�MPteڅ��r�X��JR������Q��R�o;Ai �h����"�đ�W��V"��U��Zs_��R��569�[^rR��Ȉ3V�*�V}d�r7���EYWg/�� s���أ�{#H���.*����I��Z��!"d�r�c����Z��_�����TWA���OM�Q��!N��
w���w\�ho
L/š_U��#�EHVC�{�E��q7] ���Z��&�����f�S��ϒ?��kX�18\[��/�İ�c�=�������h��.ܯ�SJ%y7:t�6��7,��
���}tO�`��e$��\!�,�y��ZU��9L��ʥ�}��^2br�(����A�s)>�{�9@|�h�f��m}G�UҺ�{u� {w�|�By��"���e+��Lgkp�s����ǖ����,����n�z�!2+\��$�T:c�a^,rCOV��֨�g�~2ՇS;��vE\[�����Z����M|����Hg��e�+#_Cpi7-0X%c�d�b�r�Ll��`���$�-q�[��'����F���'γw	�L�*/�%}Q5��\�t�mx��%�/Pmj�S}X@7��GW��^���Z:�q�;�R�9�ڕ�+�.4
z`�HUf�T=�tݸm�n���&z�	���d7���w6�1+�/2i���~z���(�N��ȩmMx���_�J�y|�����+v�?amnث�Q@h۟�Y��+�XN�� �+y_^�}�S��M�����}%}ܚ�b��E%E�=b܉㶥iF@�FBI��,�D6�2A+��r�B��&�#p�O�q3�����1e��ք�~�#��ѮNEv4����B������u/`�<�"4$�� �,���鰅/S��%N$o�ìR�v�"����F(����S�X�_�dO�ˊS���-��Ԓ�v��.\�r_��������)i/y�k�:*����1b��Pհh�xd_V��D�1��0�tqG��p0��!�=�pI�7�����H�ؒb�G��� ���r�Oꙇ�k�)�֣�����KFfp�5O��!)�5�?�EPN�����b2���[}��]��C���.�
O}��/5I�m:����uŷƥ��������+��Y��N�xw-Cu_Z)��W���6�)g<W����u�y�717"y��z,q|���H�%G������'�h|�RGo���JdX��))�W<�+�����ӻ��E�j�@��%3z1������B1�J��h^���]��/�?�鍱k�sȚ������}�9���p��n��N�J<8�3��!��Z\��q�4����B�-��Mv�d
Y����XS���������f:�f�=�t�$m�n({�u�3�"����s٘n�v�E ��%e��c/q�#=6�j���d:�O`C~]�?�ل�s���Gg�!��"sF��v�����f�8��y�c�2X �K�(�q�4H�-��1�^4�t}��2�������7�J���PV��w[�IЦ;Eۖ�}�T#|l^R���j��;�w�B놁�A��$�� �e�ƴ�WvQ�k��0K|��~��
���E����M���uZ�"76��{�p��l	���/��и��:T}���bd$k[]co���j���9sZ�uc��9�M�:�!��'�%{GM/{��}�5*�(�,���Y���ڙ��O~�'3C�\���=@�P>�fQ��*�(7�o�)s����ۣ��h�yy=X�XR�B5DG��/����Xzn�km�����# �B(�2�:6�o��!��g�%[,:�C��80M&�eZ����O&+�PO4�Κ�c*��xo�9��)��T|J�b؁�>;H9L��Nkr}9�>�?�x������{�9�Ǘ[��<ƑDA�!�xn�&��y}:���|#TQ: �z�-�����}\~fE�I>���}�&6pa�g�32��	�_`��eEA$�e\%�4=ɝ����Ya��
�%� ����� ~S��8�DmF���_v��<.��X:�ab=�"MqM�)�K1/��ODd�]Az�aI�
1�Q��ªK����t����E�co˸�l8oCɟV� �y 7::.=Q8��2�i�g�v�}���b3ꌴ�U�ϵE!��7���]P�4�cM�S�=�E��ʞ8BG=�}-ޔ���Z�
{+"���^Na����H���c�Ή�A)lf����Wxv��<p� �	(Iθ_E��=�������o�4�9J�e�
�G�_9���A&���1��Rk�я8^SƈlZ�	�U��ŉ��^��V�]�לU��� �����ܑ��ę��1�Fs�n�[T��/�O�]=��dc��O�kƓF��6��ث�n�Y�^�ym/�X�mt����}~n�����<�]7�v��D�&��8�dHJ�l7i�ewFZ%|w���I�<��F�YE�jт��g�N��!c�pZ�\ *7�+iӲ�/j�w�%�~^�n@L�oh1�N
�Fv[}$��mɲ�ѥ&t�~����w�^�N���.�"~ȃH���������$�kf����z#uz�>����Jp�ڻ�<0�����H[�������]|�D�t1Qz��3M�F��^
�I�9P��*�P�OV��2d�z��!gU"8�%��\x6V�~n]0HP�X
��%G�:dA#8�҆�Tu�.Y�A�N������������L�Y�@$6j,qP�lis�&�`�������������/��-�X��#��s?워N�;��<��y����5�$�ǉ	���i���#)߄x©M��q@5i�"}��)��*H��[Bl_��DC�h�v��������[O�,����%�1ǁ��"�푕�	��q^�u�v�L������>h?c|Í��C�mi�XO��uІ��G�k�q��4�Y�n�)�{no=HOã��J_d�u#�?^/�I�{b�)�8�1@�! 8�w�W�nr��5P{�&�M �����t�������
�P��&>'��r� '(�I�����q�2͍?�'g��c@���H�i�J�nU��Fqh��4���4H�m�����]k�:��,�;:j=]�c� �('����u�����U�b9�f�j�4j.���:8�{��2��G�:���a����P�#Zw'��?5��!��!�ih�����ϧ�"�aZ�c����m7�9�to�**�K�[��H���'����,fj��J���1n�m�C�.�o͝��b�b����v���f��(�����dZ!������C�V.Q�:?��O������+��B�t�7���wx��	̠�$[E�)�ZD���iW:ʓ�ggz}̝�|������P"t~>�����bN�~ؕy���4�a2I�?.?�_8P������"�Ԩc�(��Ϗan��K��'h=?�m� ������ ��	$9�C���5�.���<�8#�ڜS,{�X� �j�Ĕ�o��F�k�^w��3�.1�R��'h�C�CcPL¼�p�暏�A��Kz?�_�2-;ʜ��T2@ Bk}6�FA׮����Ș��c�F�>��Gp���0ͺyH�oem�C�{��h�!�U�ي�s+�؎�H˩�ת-�k��D(n.Zֆ&K-�:�+q��>���Qg������g��H>�ܻ��t)�����s�`w2���i�T��-�ֆ-��ݷ!}�e�4��s��B��V!X��J���Wbq';k��\�.�W���ao�@Z���)����g��*8����m�m��Em���AG�ڬp[��6��l�0Ȧ�㫕���v����F�⿌�����;�9Q�Ȁ��\�zG-���i#~�
�}�w��HUPnJV��Q`/�yCX��6���47���w�u�>�^AXt'�3����?����sS��G���ଷ!6��>��mir������kax����M��4���5�O�*dn��<A����'!�7Q`�J�d�@މQ��ڗ���5o����8(=	&<C��f����L(��Ne��+܉�P'�+G�<SA��	]�Ӫ�-���)��c�T��d�m�1#��!�6s�����e�UՀ��휈U	0Y��_A;sKy����H�V:��3�����B\����sʦ��Y��]Z5Nl����٩��c[�U	�.��w��V�?�B�f|y =�h.��̾![xm�:���?����H$�"M�v��و6�.��Em�]+Z�]���.�x=5�(-	�Ǡ]�Yf7*� غRy��;��V�G1X�aj�Ѹl�n~;��یZ�ebdr�"=DZ���B^|�p�Ir��V�1��&L�d��Z>�c�T��j9v3��ۍ�%��Qc���`�P�`S��4�h�L�j�W<�k��L`�� #<���f�7�o�)����GRs�r�2٬�u
WY�Z��G�O
�<`{�]�S�.�S��;�^�g*�GT���d��EcfYd,ט���������C����4Ÿ�NwML�}&ME[��s|f��Vw���pӗг�۬A�;׏�o��3�s�Np=:/{����	}�@7@��O&!�� G�"�A9���c5����X�{F��ؘaKWjNc���XK�dƿ��S)�g����JT4�+Y��=|�TL[:��/�q�y��5��8Y�f)�yL�dd�l͚�:����x�S��ڊPD�x���BVY5͟�6$:�sB8!Y2�  =�`��Oũ&!kh�S���`�S+�l�]��
�`���i���:xn�9z}�
פ���N��C@h���M�3��02�z�@}Z���Ӹa),F��L�I�:6�W�'g>�K�>��>vĤ�	�ߎ��D_�hV��_>玽���q�Sy��w�߳�3h�@��=���i�x�J��L�{��/q��r6����)k����#�d���,�i��%lԗ�0���vt)�����׃.�c{h��-��A��Y)S�pjsS�RA��Y�:h҃(�ZMo+�.`85t�h$�]`6m��^�<�,)��-�I(-G�%B��\����LȤY�|UXK]��x�Ul��&'�
=M�k@�H���N�d�_�9!<��SdA
���s�{~�ք���m ��/P��]�`9+D�ت���������'��I�e���K_E��v��j�m8���ۭ���i!3���2�O��cDm6����Lg����dw��x"r�9��S�f�C��=� �3��2 �r��5��%6��bC�^d��%�ɧ0����Z͠uj�%j��u'�xdn��τ��3�z�vu���#���h�n%�D6i8���#�LX���d�J�ޢ��^�#�N���=1�x5G��u��h�_������aW��C�7�cV7Z�Gr����V����e�8s=�� T���Y���>�BPj_�v�':�/p�ؿo�qu�X�p�]#��b��]zDva̸p��8� �C��:So�&B����ǎK�� VT�ά�r�A�X�{�a �7a�χ����Vn3�uH��*���U6h �a��da*.D���f�n9���r�oZ;��$�*-M깉q�� ��i;})����]{��o_�	�-ciLqg�o2٨�,�Β�̫G3�_�\,�3��#�I*����0vr�j�_+��˘v|*�gV�����0���7��8��W3t��B�c�B��t�{�#��7�U�^� H8nMm�Md��>�U��>��yNn\��d<�<�f8���{<V�'��V���K$$������� �5�����j��hB���O�o�����m�в^��Y�L���e\�hY+Ee�8��攼^��P�N(��r@�{/!������=K�O�8�u2,��	B�:���Ý���Lc���7z��1��o�c�2t�\-e/vnщ���Cw"�� ̢�k&�EG����i���6v�#Sq�n��̪�x���S9j?�\�V�X+Z��ذPG_�{[�]���`�,u�.su!, `r�b�i�Kx p�m}0�'���I��5	��O-Y�eH���|X�#��4m݂����f
� �xE����� ��RZc��9�b�n��xoT9�vH|�^�;�r'�(@U�*$���f�[�7��+"� �U	�l��p��}�,R���$�a@��0<T�� �����>��p�Ƃl,X�.w����c�2n���q��Q�{���"�
]��B5P����q��$/@vPܒ2���K��Sݯ�os@9mG��1�6`���bK�T��ʜ/��6�.�^��Q�b���+�;Oi��Y���� �:�а:Q�_�ã'&<_����>��� ��Ε4\��3��U��� �������^��{��y�blU�#ʄ��`�_M�w�>%Y��� z�W��Wg��8�,z��.��C�h*)xG���ݪ�}U,��V=�?P�W�|�L85>������&���&�������%��ѳ�{��n\u2쯀]w	%��"���Ы�a:�M�q���:��/���kT�����.�%�f%��g�@�~Ԇs�5
�h�~�z���]<���;��Q��*lf� �P��,��m�<%EW+��g6�'�4+�`Z������k�u���B?���0N*���V�.����j���[��^���#���=,M��8�!��/����}��і ��<��(_�+�ϫq�XP�p5>�w"Q�()Ц���s�A-�� FL2�u]�[g��1�g~Wς͋t�U�M�E�Í�≹�8�]A����<;�!~�t�4�<���S�N �	�V�K�O
	(���R� �H�@/����NI���kh�"̬��Ѩ�#])h�Q�.L󙢕UW�l�F��3��w�lķ��	���]G��qz%��Gv�ǉ�d��܃�TQQ$�
�f�,��ES����w��z���3׏CG
�1�G��ǭ���U��n|?�۩�����z\��<w&�j��8{.�'�U�]{j�P؝��a`���&�<�8�q>L�?���kÅӧ\�{J\�X8a҇Kݖ~�l˫]x^�Y찘=�BC(�X:��};z@���P� .;c�����x�`�]u\�(�12J��0aɫ:2�uӨ:�3UַuhŁ�m�b�FFq�� �',Ut�/;Ҍ ¸:�@7xz#?�wYN�sT�QI���%aAB�:V���pp�k��]
jɔS~�l�������|�m\�6q�����r��>dG�N����������[E�\�����#�����~ͷm �#�V脖��w��++'e]zm�ۉ�� ������:����-t���7�(��1}|��ʄ�eM��6�qy2T��^l�d~��A��Ӂ�rTZ���V��w{���@��]�I�����P��*��W��Ѭ�[���4��j�?i���0XF+%�]4�"P�˾a��|��Z���l�wm�*�}�0J��g�r� P&�*,Y6��_W>��v{����f���5�n(�ֺ��:�I���)����.Um�m1N��J�m���(Z��i<-�]���ڛ��(�jV���!�A�{�Ig@:��4����ن�(l4!K�X��0_*�	���Sˌ(��k�
�$�g	�*?�\�x��Gf��٧~���gM�ԹC�Z|���"�z6%Hjpk5��`�16���������iPq�5�1��bL��r�X�d��>��i��jK�$u5����p�+�|Qc���=�-IJA`,I�t��ݿ��Nvn@��J�jѩluk�=���f>�t�<�z6ڽ��v��B(-f�v���/\;�K|:�~��[��9)S�y�Z����/to\+R4 j�~*�ҍ<h���0�Ty���¿�3@(�K/�A�,��*3}����b١��'Yh����~�mߤ�������g���T��IuAid��~ǳNF��*NT�\����gɊ~ʇe]���z�6����z�x,��;,�|
D`�/A�8���=$Ņ}�/Z�a.�AH�A!n�@���ᓆŖtx��_W"��#���0�\�[��e��UW��)E�sR�E{��~�P�C�>�r'E�f����LH�t�G���Ì,w�~S��b묃P~�*�!�WR�y�F��t��U�1)J,��5�Z�R��sg��q���M�n7#�R�y.�+x|K����1H��}�o�
P�A(Jt=���m���nzs_tխi���k8�a��tn�F�&��Y�k����_+��T�b����9�y�͠�c}�������O/9��sm@U�Ky:�Dg'��Yd��Y�*S%���0�⾗�+[&	 W�M�{Yհ櫂��ȿ�X��bT��.m\�o2�g�KU�z�-�*�~��SxM��0.mnh����f4��*K�&�M̡���DKgg5*�0F�u��|>2�a煳i�fo�}5o��1��T�-s���g+ݭ`�M��b��O@ڤ�!	MMc6%��pM�;��r0���9���.5R�J ��;��Q<=\R���[�ů��JT���=�!ġO�6�A� �DkT۱�}��� /��Ә3��(X�� �x�v>���̋�c���2.`�3\$5�^!�������9�'b�a�e�bQ���$ZD5�����mu4�<�P�[%0�8V5PԦ팡�|D�X2�gX<n�����_���!��x��N����@]���J��Y��Ǻg4��.m\#���;�5���Փͺ���l�U��	���"�p��?�)��Z�u�6�&F��^��5���� ������Zp25S��9�e�l�-+�����A���&u����0��$�=��K掠i�)ܔ(�T� ��j�h��c�5p�C���6����OI�6�
!Pў)x���c�8pZ,�*Q�/p��_���:ؼ�a_IY��B2d՘�Y �uhR��x��7����]Q?�\h'ߪO2��3����,'P���/|�E `l0��e�5���h��ܷ�y�[�v�V�TH�9�e�¢Pj[������H� S��X/>D��-E��6�'=�w�A5�i��f9Lދ��|������{�4HAc1Wj1$�l�%y�.ٗU����X'6ڄ_�5ų��N���ac�r
�t��f��0���(џ2�XN�YչْM��{��)�$I��ߗGXD(l������0��b':��J���/��*�5�m����vp�y�UyER�xz3Li��M���e��M�ڮ|Eo�����}����S������#�tvX2��@
V,���<��օ%���]�_r�(����=>ߠ��U+��
&]D����j?��r�;�x<������t�[RX=���z�H����9���>7VYcuu���~e�P�Cr�9�.�<Qɥi�7�V�?]Q��m��L��:��dϫc��`� ZHV�|k\!g|����ѦS�� ��J_`_�x6]�3w���՗���&�3A��_��ů�7!� ��c����lNO�zөz";������`]s��G�hY?���ٗyO�("�0�mÁAR�Ba