��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0����_���3���eĭ)|u��XXp�?b��&� ë����
���#�SDY�91��C�K�Q~�j����Z�����q�Q=t�5��r��g$�#'�1+������V�iE9x	��գsl��h�H���>U%ڠ�}�����O�������^�B�����ʠ�i�����v����w�vr�mk�{���avL�ݿ �gx�O���X�c&][����G����PWE�р�lԈ��l�ͬ�W�[�|?h��rt�	*|p4����;	�dN�D������x���qܣ��}���Q��?���0�ˉ��F=�!�"��p��!薬|bNhiL���H4��Ԋ�|���);mr�h/�TN.}��K�-H���r�P��i��3��1�̸��-7�?��v�AR�Z�؏�#x��N���$��C;/��2~��I��}>7s�<�A��hA��Y�>)�f���M&vW�|#���!�ltF_�,_�V�ӧ��]��O��y��}�YB�ǰ(3j��@��J�Bs����cWG���!|�q0x}F�oY�� [�%:��`���)T$gQ~ B�	��[O�W��gg��$k�� (��g����q��9.��uf�z��2�^v&ў��o_�k˲�>��"�HE�9c�8P��[X���B9��U�����S�%4�rf�B�G;-�Q���z0���g�uʁ�N�7T�y��z��;O��H@�d�g�A ��!�v�IU���e3�n���/|�Z��m#������Ƕ�q��P+��A�_�tk��	��0����@����^J�x�nx%>��`��A�����f��E�<�M\8ŀ�.8"�0հ]��������;��y��*��<L��Xn�gG�V[g�s�k�� ���Q�����%�Q�;���rP�9-�d�T˫�]Iّ{8��*���%����Ԧ'�����7)�>�����cF���C�%{=��⥻:�pQ0���ԓ��OS��z>f��Z��$��A��:O&M�'Хp�e'��5m1<�O����N8������b�:�f`%�b4����شl�-j�m@vʕY-X�Uh;A&k�l�����X�
�°Y~����^���R|p�R�O�����0_�:&�b�#�nR���_�@%�<M������,خ]{����1l�d�04�
��pE�u�G�T�: �@D�������4�q�@M�`Mp1<W҅N�wmwb�_�`[�^t�[/��Zxg����+���XD�a��o48Ga*�I)%����u��-*�!��zM�M"��^��ǲ��	��O�K:�$s���hL���m�=� 2P�Ӆ��1�(�a:AG���v�t�#8T�`�$�,�DAZ��?_]�i�WI��Ę����K�KC�a��l6�)��Qh4�����KB�"K�����~��Y\]�`d�S�*��ǌ��T�KW�mk޴>t�{�.�gz�2x�	��"K/[3��i�X ���RQ��5� $�����}F
}�#�����QKDB��6��4��1�y�8\�'g�g�{[�~[R�H����MC��YP�O���3�f� /��E����_��y?�A�2�_�b��	B +�ޙI�p� y@[���DY�I,ݿ12�A�%x�I���:����$*z��g��'��t0���I�K����;1(�:%�e	n�L0LŵR�o{&еC%�X�o�,�@)𑞡���#����%0y F����:�,)ϕ�Uj�^�d���/�%&aY��II��"����
�'��	�lӾ�C͜<���T���Ul�5Y[J�ɍ���
��/�E��)������l/��o��KW�r�����YY�<��܉C))���<`��}�B��>&��!ͺ�������P}W��g��$�����r��(��]쌜��l�f<�A���<獵P�;v�a�����R��=%�쵤z=��͋���B��q�ϺSpHWN咽�q�$�ha�Gݷ�0SMʦ��%�����Z��u��7㳯�}'��
�Gk��w���!�v�@ L�h�+��V��R��:�*�"TDt�f�ò���YG�87�c����B�!����(V����aǭ8��[
!�3}���j'��(�D3���2���t+0/�6�<�t��S�f}u���p��� �ZS�����$�8[�7L��+�X^.��'�Q�E�sOS��"�r�v)2�{�e�����������G0�2�/���Uwu����9	D�s�����-�6e�c;�7��V�%y��RlT�"�"�W�����C�Z�$�--	
��j�f�h�w�)�B�$0)^��*[m��ۣ$]�ֱN �x��73]��F�y�I#nMnJ%X<m�n"\�uF�w#k���_6}3DD�FX�I^�d)�����h
�+�	��ĆV� EK�w����X��5���4�7�օg�=ؼ9�<��C���Ĳ+#w�KI�<�"[��h<���w���D�6~|K&�`� �%���A�V����p�
ՇW7_��J������"�"ƙ���{�5+����;��W�t��^�9d���'w
_�b�w�
;s�G�I���I�sB��k~��D�zɂo��M�/@�$�?͝a�z Y8���W1�@Ou�C��aVѥ�	Ŭ3#��g�U�bn���<�ĳ"�w�r�=�¯��摸н��9~&�����%���`)%;��'*@���Q�&���H�e\��:6���rf:ߡ����_���R�[�]�79�W��!(�^�0�%+���,��d[�23D�1��r�cI��W�db�+Ö�W�}��9�)s��h���8]�\�Q�7țy��uЂ�)K:!�ނ�~5'�ݢc�
5Hm����(���� ��O]��ܟ(k���mǯ�66�jB�79�����* ��dx�Au�3j'ݔ`�#����矍�4�~��Ɠm՞�N{��)�G#��ՑSd�,���'`;���}ɿhg� UW5$m�v�2�5�E�߯Y
v�����#��O�=b_���
���X��փ��&�賔��ڡFk�����"�+JK�_������ÛǸ����%D��	a0:�@�B����]�I[xs���Z��oo�!�]�)�9˧�\%[hۜ�5��Kw��ZN$�)�P3��JgO�,��J�b�<Nc@ok��I΃��_��-�ߛbd���@�JH4�Tk�fWE�����I��<�P9�>1��pp5. p
�&����s�Wh趈�?�E�&}���:��h��\4�rͬ�h�RX
>�Vv�d!Oԙ����z��hQ�;�R�%�� $gٖ3o߾�FA�E��R�-k�T�WԎz���������5T�F�ԗ�����(/E{��,n8��a�̇���E��A���j�/�`��g� �󷄤��Z�z�e݂v ��0������A�:�孧z���vT[l�@�F��KK�a���rb5E��i�(�n
s�_JiG�̈�Y�|8d���yJk�I�N�W�ձa�6	m��TV�;2�B��Y�Q]�cq��MW~��/�k�1�������aT�&-W��KC�M�l���,��^���b����n���-W�B5�{�%����8��K�O���5������wˆ=�n3)슰�.����4I�����jش۲��:! 6|R^�86xÖ���-��M a�b~�%�Y���>�G�Dټ8s5�� ��`	{t����n�y�ə�}BlW��zeƺ���V�V�l܀����9Mņ���0k��6�(��jy�AvEB���}�F�b]�̐�Y��#v�b(nv��i��A�����ǜ�T|\1Pb�5�Y0,����Lۜ���l�ƬE&�l���PÔ"u4��4H�k[%�z^�����"�O��v:
��c=L�❷�;L�����U�õ;ՠD��L����,��r5Amt[���Ȃ3�[rj�l�ψʬ���	��yp���K���@�HI�T%��q
�^��6o��bp��]��	>e1�ڱն|�äA�+mH�>�3�Zp�%R���/��R+����5~Z�bo��x�ީɔU�:+hRŒ��&��vH�'|o���~mPlzK����ՙ_L ��Oҧ�In�&���i���9F('�v�����&������Go�XB�̟�ګ�OA��x�4��Я�by=�(p/Հ��%�!#�za�DE1���'�"�[�hV��ņb�)����Nf�Q����]�m��!���,L7X����U=j9�NLJJ��c�jQgܵ[I�ε[���_�h<��:�%�~����@������Ԇ��?:�a�	��u�_Z�n����̮�ks��"��4cN��r��6J�E����	g�[D��hk�;��KڿO�:6}E9N�&�=3A��K��A�k���~�//���ޥ<R��v�Na�P��7�rT���Jm"��!a�� `%��6��t_�ƚ��J+{L6�a� �$�˹�^�E_��S\����C(FQ��^��Ř����<U;*c�����=�a����Kl��-"L��f�Z6'�t��ҕ��^�rC,	�jWwu��,9 | -����M4^�`q�ۑǧ�
��{�b����)��[�V���J��~'(�m<ĭC-�]�$����D�s7ut�C=A� ��:|��8˫��� �a��^���zPh�`�]�Ʊ�?� �Qb�ܒy]�"�U�CsY+]�|�E*Έ8��܆@���\Px-Dw&�q�p�%7�N�
G"ա}���Ƈ<�;����Rj�G���������w�ŕ'N��IL�w����jj���6sm$�+<#1yy�b��G�p.�)':/fM�NzxoJФכ/���c)�^�}�h	��ң��~�۳&¬��H�7�Y;��c_a��l��gQp��1����g����3")��j*VH����k��esK&	������wI� qP%g��[��ܺ��0nqR�·�(P��=3i�5�wPh,~�!
A�+컖��M�'LA�R�b�&!h�5��O�گN�7�����C��Y���
VK�:��ac/�gd�Mt�f,��z�!��>x���A�G?09��$$̝�֛��)�Jblo37W��mF��h"�z��fl,>��;���#)N��A�t��E翹��+C%:Y�vW��F�j�Ŗ/{�O	c�~�S�n#
ō".�ҭ :�r�M�?Sڨxu�F�0�J�#�.��rn1�SV}�7N�|�FեN�hY%�+U������S:TA�O#K"�$D�֡_((���pٔbݜ�B�������2���J��B����J��{��2C�66��9"�t�$w�J@ΟJ}~uŚTL8@g�B]���L��R�X�>ˉ��k9o�B���Y�mi ��2Z���Y�c����u���!.���%��D���m�����}�� �QLd�X�K��8ΪW�$q��V�&a.,�{�I+�B�ohZ�O�1w!��a�����^|�jQ��"o��~ݑ{3*?���[ q*(k���M�����$<C��E��P�0�X渚>��ED��r��9j�y΀�V�<	����VC'�tI�l7��g�s��!g�SL���-6�f�~k�cD��˗m�DZ����l�pf.E���ȍ"����M�9�@�u���>C<J��(���<H�r�`���l�:��82��Q�<gm8dA�u�7���'� �t�o��y�����ȅSI06�s��7����͡���hiFU�u2N�C� n|��{�+S�G���CO>-�,���q�_�/�����H������j��D�������p�0�\l�y�:Y]{�+Vͥ���,N�w�}��#�?cP�D����Q9���#%C�	�[���5�b���3�J��Y�Y>�Z��@<�pޙ���!����Y�l`���΍���`�Y�kD]U�<�+�7��;n�Q%V,�RA`��P����w��BU|��
W��M�1G��.z5���Ǘ���|=h%7��n(`���''�f�ᵪ��<��1�m��%5���x��0�H�a�YB�ɠ#k���1�,��.$�8S��[Y]|��V�l���䉝���b�V�1ќL�� �c�zc���)4S/��I۰sed�fm�j���S*5�v�RV<ž)%Gb�C�_�DJ�-�5N���;�'DX|����[/�͟䂨�P�Ύfu��_,@�]���暃� ������<3ɽ�A��s4�����F?9�A��i���t�'�sU�ex�(�G�X\���R6S�Ko�=s��iմy�yH�{?�����	q65M'F�3��s�nڙM�$*�*��晾ehc\6eŇ�A�$���O�����l�ε|����ς��00^�w0�Sf�����զ�ZOH!��J�ᤁDeV6��B:���m����+xQ|�ƫ����<��!%�BFl���R|� H;zRU��/�b|���W��꼶>%bH���x3j������~Hڈ'�U$YQ�#X��}��Hp�٪�4Q�΃�Ê���B⿄  ..�XB#zN�+��M�kh-�,P--�ԝ�����i����!���V@�~��T�'�6�B<|}�7-���!�b�]?V9����i�7HB�h�|�:��������A`�
�p"�wt�9��^��1c�~���8��'����YxI�nO�Xu0��{0u�!1���<tC��ӽ�Y�VyGP�.䴧��D"O�x�_���P$�k�E>p��WH�S褭r�գ�Nz?V���<"����f�oR*�>�W)�2�����F���$�ǚm�3��|vI��넝�]b��#@z՚ex=���쬌���O���p�I$����n0А8&Q
w��B:�)����n4^��0�(�����\��-�EU��	\?��ήP��xs�ěR)��E@��A�"O��Q����go-�jr�kϯv�,�>9��mn#| ��݌���I�7#E�w�Oo���*z�O�0�ć4r�p��i���q1� �P�mUۛ�eZ��)F	aps)��ԓH<h_�_Q���������7Ӣ�t}�D�2�8R!2�����_�З��l��2vʳ�$�49��E��ܯ�7�A����V����v�k�s�O�>~Z@�[`a�uD��=h�/�ge�6����N>aڌɦ`�s�3�8V�?���˥���f-e0uJ��y����ba�=�B���aq�C�ٖm;�ذ4��K�!Iդ�G'��A�]sd�0T"^���-\���ͫ�6�	F����ɄXĩt�'7cJ\6���'�� �K{z�V�'H��<�� �Cj��]�I��V|?��8�y�65wj�m$f���hͫZpoRl���8���P�~�D�R%���O�zxd$�><n��i�p�br��~�Odr5��0虒��M��uö1Ǿ�����V�"W����}cʮ(�F�6�Gw�K&���z��ԍ��dd����:ύ�`�]��֓N	�y�j�{�se�ګ�K�Ĝ���c��V��G �&pa5�*�M�Oӎ�C��{�t<b�m�60�o�X�6��X����rϋ�*z$@�;�{O�=��f͎���$-'��=s�r�l�R����I��ɒ�k)2����:��w�o����!j���bO<�g����X�=�3��S�	� ��QeU9�p��\��P��\r<6Z���� ��aK�ƽ'=���>����w_J����mb\�'�-䄘�����?��޷�Iop�l�����<�Vu&+���jO͑	"J!\%:b��$��4�X��,�C��~>��5H!I(&b<[8���]-VN&����ۖt��-.���d��� S���>F�"��m�˹�q&g��
8v����6��qN� nh6�?<�ad��Ua��>�=.Z����r�\
�i)���SE�~I�������]�����W���Zq�+K�T�q6�p�)pū��[qMH�/�/O��Dg����7�f��ܯ���N�b�vI3݇g'����Fn�賷`�VP����W��sFx�I�rǵ�<�P=�.�w$p�fQF�/�j��JR�?UL6˘�ہ�z$`R�����!���Δ��V�����`_�󒕄��,�N i��<P��L�',�?��׻��|�	͇4���r!`T��9�A�[�&�J�?Q�I�dp8��7�;�ԍf�r�>��� ��T��N���zi�r/�-yȤd�P���<��(6 dL���U���b7��bp'0�'f��vd��t�b����<��t7���� 5i�N#�[ҹ�!����O'yw)��a�u���������62:CgI�"P!��[��k|j�9��i�-��x?k�4/�'��X5�9�R�؎#�p0��<zg���Ўj��YE�����r��(Qc|E� =x/8ĎK���	2�‶�\'��"�&��.���.�Z_������jʎ�,�']����D�T6����%��?�WE����i B�X�M�
�Ā�ı 5��m��"44�B#�c7'Q�wc����'9LQt����e_��6�x
F,d�"&�s�\#���Jk\�ش�ִ�"�{�,��ޕZ� 6�W��t�8>ݑ�@��7��6�7;����68&	>j@���娊��a(����u`^5E��.��y��iJ����rk+��d_qE���W���y��Uj	����uq��������w�t�����߿^iH���gs�(����+�)@؜O5��R�#ᝒ��BJ���/T�Q�ue��qPq�t�*/�e�pp|]~�
0�ܕ��7=դU��L���>�_$��%��)=���IBB>�m�aZ/x,��1F��c���p2I]?�f*m�Os�f����]K��O���W^��ܲ͋`��;�~��կ�c�b���@5�h<�䩠0Q`��?�͹�5!��|�_�3�6	~?<��.�D��m��~�w<�kg�،+U5>�$@�'�=0��r8�I����Q�g��Z��w!�N]�w*A�i����C��-t�|�����]���D_ߢ�8��鈕\��%ț:`5x�*� �l!��(T�r̆��j��5Ԩ��Y �U{�JL9��d<��O.�cђ�=�'��$���gG�>�>:;�4@(�=O�h0Խ�=����I�ؼhI�#�����F
'yi!&��8�xoA���e��1�Bx���� ���v��Z��� �z�~ʶB��E�6��\�n;B�����<�'^-���j�eӒ,���v�2Ӏ��3�lN1H��C,P�Hv�3��5tz� 4�5/�f=R�:NJ��M@P\Dn��X��T����45��w�9��?�jי�0wP�6�ݣ�S�"�	�y��(�O9�޼��)�{2�G�P �H���dˣ��b��=b�0���d�r)�!z�Sf�<���~��(Gh�帥��p�!���	h��a�D�Y>���F������W��Jikhc���w�ȚV�L��e{�v�F��n�g��$�5|�(���:�9Q{/�^��i��+Q�o����J�-)_��O�Y�K���߯\V���v��~��3/\�<�
�7�i'�ȇՌ󜵳nT�u�~l����p�ЙJ%��*����\t��6ͨ/�[��l��&�"������^:+��H*Lؖ��1����_�o��z��!�3+���/@h�w�Izr ����
��a	[*��	Q�|-B��kY�����ux#�#艡�e
��"�/�&V�����������Pt-ZFzr��؍ϖ�eC�)��o���sqc����)c���3^��K��#D�|ţ-�r��Ig��@*#�c�ز!������d���E�w��)Ù����� d�7�`Wnv����ژ�=��^�,