��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0���p�?�gu:���@�6h�zj����y#]��DQ��J�1�_r�=U0Kb1N�`��5\ɾ��|�k�p�I�Ç�ek颪�^2�軬'�R�$���p�.��o6
�/!@f L���2NB�^����0��c(�l(T"wo��J+@A�eK̍�Y�	=�)��=�@V�6ᒧ�,���D.Bm�0�.0ǃX�#E7�Dߡ/Q`2�p�OE]�|t��v�je�Jm��'r�h�M)-j)tR�6��n�'5(�߱�ԣ�:^z���e��wXXir5�KFb����Ld]�aT�,�o�����zm}��1���_֥gi,�#5^	�:��e�'�8}B�q�4՝q��Cն$d��˖3��4��4Ɵ^���gܽ�Ɲ�u���>�����?Q)0�T�"��+( ��q��E'(Ċ��x��Ա��I�h�3����>�˸�g�]�D���*{�3�j�H3*�L�gb�| Ep���41y��®�b
����}�ح�~LI�,�^Nt��й1�6���� C��L|1e��w�d`5���&?b9g���P�������_P���qU���b�&���b�ajS0�i��#��9.9n`�R��7�G�;�<.M[q����u�1X��+�d��Ɗ���K+�0�Da�Z@��݌�����e�{�D�dkh�>��7�v�Q�e� ����r��8�0�ZNd1/a���ٕ���ϖ�ڹ���9Ţ���?S�/�LՌ�+�����g\S�eG�)0^R�6ɟۏ�����A`��b�_U\\|��:l̀���<|fje�7�
7 `"{��㡾�d���7Cw{��Aă� w�f	�7O����ee�a)������{%����0�LZz������(�,Rs?6M`M��Ivgg�ٹ����/�� ��R�4�#���8K�cr�R��H��г�^x�A,�B�@`��49.�n���ƻ��!�������m�\�E�Ҝ���^�l;��}Jw#��2��!��|�Q��_��=m4�id�͊�#j�F�ѕs�-o~Ӑ������šJpT��!W�ZNC�c���#N@��i�����1���HN��M��Mv,�[w~�+T�����-�t|��I�! �+q`��M"H�:Rv�D<e�\ʂ�� �&[+�3�M�0����� �*��b-2��qN9��T��P�g�s5>/u��.�g���bX��X_W ��D��S�$���$��it4�UYg��-#����t8`�����M��Eԡ�zҙ��/xЯ��q)""�^�+�y�Є�q�¹ ��΢�w#�Ia�3@����6�jd! �����5@F��d�k��t47���!���L<� R�}����E���lړ����ƓUE_��M,���D��/�{V�XUP����j�'Tϒn��˫%�%���s�Į�"SB���9�zͥ�0�(-15�5���%�>��p¾ہ\D~��4̝��]�9/~�<��&)��Fv���������zE>I��A�yUcj�_�^�f�p�c��͏���f�V����^k/���:��A�hNo�l��]4�Y��xQ�,Il֭�t%V�auD�4$�v|�u�AeOiZ����H��y��\z�¿L]��Es���2C�j��&F0鋊�Ǒ�w{`wc�v8Z2��ZG��tUH�s$��8�O�l���(c�c�R�=��/wh��'*�hN9��e������^�{�^(���j�ӞQ�� 缳A!���g��/�����3��cvwv,D ����������д�1f�	J��]��HKJ��ZB���$���c�Nڧ������X��"������1/�w�mW@H�LQAt��gg�-~�QU�?�vYJ��Z5�.>`�
nԈ���C;w#M�2Q`z�@�=�Uj�5A<K��$�4Q��(@`�ޤ"�ޓ��ľ����P�[#�.�8Q����]��C���$c���j���͔VX�����[�z�ӧ����ӁX������<�����G��d�a�X�9�`�JHċ�*ЙC^Y]w�Bf���R� �W��⇶��tQ�ؐ�b����!iN=w3n '3k��߬8�-1\�Y.���<�a���F�.� �����8�])���S5�X�o<M$u�Ґ�àHUj�X���q�k�sB��9wh�5�ѫ�^�h��I�P�����"�g������a��ׇ�5�>#�L�GS�����`�l6���$�4���OQ�5�ZF4F��)+f��~���Z���7���x"�[g�%��~+��h��Ȼ,%��4�W�K"�s��R��αU	���og��yR��"ˠ$��oޚ������[u���Q9W5�Y-���
"7V{{��(�/Е�˄�(|lN�OP�md����!��P�	4 �%8볇�M���$���o�~����e�F~�9��b�LG.6��e/�	���p�P�n�4�	���$>���*D�O�����ES��� ��r.k�yM��l�_R[�XR-�':������ε�]j0����=���_��v���ci��)Y�ӎ��]cv��:}�>*���{4"�r���ا%r����G��B �-zg
w�}n��F2և��
��U����j��OHR��;�Vk}�I"�qc�y�B���ь�	���|��w�>���ƙ6���i*ڜ�n�۸�A� Zߋ��$��z�?��=K��B����Ȯ.��wo�C֬9OS��T�*�Gi|r��pM�p B���fW�%�5`h\nk����)�)MX@JO
��Wo$�Q<� HJ�\����9�=|6���=t���5C�:i�fQ�Bw���'�O"&�
c�����%A���%ؠ�u�LTvK
���&���۱�daQ�<�}d����k���;�@��[qz�}�6�����E�c�������2_��I��~�
�'�n��{�w�����-T|a��x�Q}�����F�L��Řq�� (���hRؓ�WU�`~D35��&9!��)#�!�YT�rg(���A�$�9mu������~��0jC��+���*��v+w���D��I9�n.�)�ιW E�&�����N�k����%�k�p���i����,�<��
:^KK�e��Yv�g~c��G�'[�Q�	�J�8D#ɛ���j��������pB�Wp�=TIq���Ux]UE��|ZD�������x���*�ۀ�fE�sꢢCH6s �[Нx�qԏ�:�Ԃ��ӌ hY9)�B��`�GQ�il	��f�K���?���i_��Rh��dO �t�����]��=SևS�̪�4�y���ѯ�%�Ǚ���B��-�����f+���Z��.������G�?1�b?ƕo�TLH�+������w�6�f<w���7�-�<ǖ�!5k=7i�L�l=�ӝd ��7A
aM4��o�5��N�4�|��E��N xUW�+����Z�W��B�X�&�����%*�ZA�F��(�ؔ��`S�Z��5��B�i�~�����"��&vD����p��p��E`ar�����4s��eNc=��Otr������¡2����#��o�`/�H?�q��h$�FB�`���{��R���x{JD5�w��ʨ|A�T���䆂͆�Y;�N1�Ǹ�!��p��5�J�m�k�����NԒ(̔��Y���=��$"�Wp���ƸB��Pڙ����ۏ|�ۊ�rT?_N������e$|�8��s�8�Y�1
�l~+;dc���ÖT�f]�`����햩�"�Ht��&w0�5�l�y�������߁�Cqop�m}���S%@WM41��3&��Z�J˛������v�?���H $�W��@�;A'�Ue�u�Wl��'�A����d����2q�iL\�����&�r�ԓ���S���5�H�0G�&FD���VLP�ڧ$х,�@,�8��(��-ֺI��qJ�����j���}z럿�Q1]Z����z*��C\��(�I���(����񳾡�x��5d]X��x������Hs��9���U5�6}�i��η�)y酏ԑqY����ɪ:s3�]�`�,چ�p�U��� �v/��lQ0r4��N�:-ͷ[n2
���䬉�fc��\W�;7��Uf!⃭��wk�V�����|�{{!�Һ�B�=hHs�}�����Z��)�*�������Z3=�ՋtDb����ӄJY�e �X��w[�t����	��,f��T���H�[&�!�T��27��30��;A�:i���@��q�}i�X�jkm�U��X2�%�o�Km���ϼ�q�nmΎ�O3��Obg�����)���2?�15��
]@�9U*�������7��3�g������t��l�TI?r��Z�f�G�����x��m��^�?������~R��Ġ�m&Xg�.�ʤx�o��{F�R+�%���cFJ�Ć��v� ���Y�a�&���_^U<�6:JR��6��_��Y}�{�e���\ޔ�(�Q�Hx��Џ�k� A��-������D�5S� Z��0��)oǣ�e�M����@��)<�+���!��;� �x��v�KQ�Rܿ89w(�31K�	��7�Wn-�yx�o����	f����<6���_+T�v5��o�4xr�ϊ)P �x�&�>';���UJF�
i��,�_t$0+8냸��s��(���t�X{��W�6�N��� cܞ *8d�4�\J��*�a<}i�[g���4����n|F��p�t�����qoES��ss悆�y����"�0ç��3�E+w�.�kE����\�,��,l�����Q�É~�ԅA�y}�c��-�uk����.�~��)�w^�����g�\}^�- �J��<��"��A>��	N�f8I����?=����θd��՟��A|y��ܫPi�Ňo��{�Vc�M�՟+�4�l�J#��z���`�Gw4��~�,�:{��y�RϳU�bLĵ�iZ�P�T�Ĳ�u�X�鐙�~��5\�ρjܹ����_�y�ƌ�:�W�J�ץ�� ��tn�u�ѣ{j6b�H>U	@�k�����3�����`r��dd��.���Y�KA����`���ۻ���l�{N����
[ �u�hcۀL,>��e�z��#����c���ը�Ū��x���q��j-Tm�P�ޖ�1n�4!M\3.4�И����U�;����ibO�/Fqj�_��j(*�V]=��<���eA��s2�s��n��h/��h;V_��)G�ǚ���O3��8m@�r(E̙��M �@��{`�E�=��1h��j�G�a�+z��<%�2$7sf��%�w1w�`y��b|20{rq~��!Ol��6����ݲ���]3����+Y���J�f�H�֭��w:E14�����~8�V�'�O_�,�.C�����tQт(-ǩV�	���^:���	Y�|YB\`�v�~�J[~�a�3����������v�x�gb��S��<�!yص&���H�T���d�#�nޗ���T�`����,�G\���ٚ����!"(��i�c�ݒы,��M#�2�=���h r�>�a���A4<<=˗�S�>(8_vOc�ToǶ�RkP�!77|� 镍�S:����X��3�� �-�:3�E���n�z��{�kS<6�R,Q��wӱ8N��S`�[���e��T��KO�G�tm�����u_��sGna���Sk�fe��p��Ն�$�6���*��P���=64J�M��1�bu�Xr�_!��e������pM+[ht~LԠ�UZv>+�Zdu)���j��8�K���:C�I;;�iCS���!�t���1<�U�Y2jX����ßb�%��e���M��)�Zd���΂
"�R��E^}kIPI�� ��E)���� ����VA_�l�M�&�7e��g���"��HǄ9�˓?N�Bs¦D�2��]y�6= ƣ��njڜ��s5j�L����+�l5=�;a|�k���~������	�Ҡ\I�B��u�Ft��:s�8/�j?b����R��{��%t����o�n��������jrhUg�؎���,qAnQ5��L]a>!':����6ԗx�W\l���~Xajr��R�!��`��4�PA	f	��ڎ�3�w�\�@)��k���r�Yĸ�,R��2�{*,� ���;j@��_t��T��5��@O���ña�S��#'�G*�@$a���_��r%V��VTn���T��rQi��XRAr!�3@&4�];6�b��lrB�=?A���̰�#��Sr�8�Ǣ�zu�p�#�÷�K��	�oJ5����1Y��3)�!�̓F���c�B��50S���6�U�^�O\�Eck�tf��Z�L޴���KŃ�cf�Ȟ]�����r��˵\	D�3����T���S)���=9qnIC�xayb�4�C��_69�u>��|��AL�	��lu�l]K7'q� ��	NgFc��̎��m�J(̅�u��}�G9b�B��8�"�["Ha���[w�:F7���3"s^�Z����S}���*c\����}��Q�&��IG��
�v-�l)5f� ����YKW�顢��1�������f���E�ꐢ��@��(I�I=�FY� .��)�as�O��b�DI��iZ��+�Գ'�z|[�V�#�O)��OP�Ws܊W3�˼)=�OI�F#��R���!�O�c�G��{��g�Z�DR���͗�||���4#�L��)��Q�W�=c��!��Jz��g;h��a�P聯�%��49��Q����jH��6�{j�nχ��`V(�A�	;�!���!?��L�J�g���9G�^���>x>c�!�Z�#�����a&�M'�(6����_u�Ж���a��@#ٝ��s�Q@$�Zz��G�j��yŸ�b�kV,��.�)ש���~a����1gs�9SU�-�>=�-߀�{�~� 8��� �|D1&�����=i.��v��>�B�`��b!8��-Q��{��Ϥ  ������V���ү�^T�pu��$D,� E���A��+��*��3$��gL@'�D�N�lPj�d��?�>��*i��W���۠��?��Pd��(6��%�"�g"N:��<@k������x���zYd�'�S���8�J�kbfY�v�����+J0�OSgJ��C}�(2��3^@�g�	ʅ5/������X��/4f�%L�:��]����+ɓ�E��BSWT�	�A�ӟ�佫?��TWx����)�p�_�-�̎�x��*�ּ~ʈ�����x���r,55���y6����(�(��jnyi�p,��X�(D�V��]�.t���5�%�$�_�Bε{�=eaK��c�Z{�X
=���YU�|O�\阖��&E��t�_�5�gW���,u�4g���5�3!L�8�xB=n&��RuÆ߲%����c�\�PB�Ƨa�	���sy�> tx�uו���I&R7�ؙA6n�{�Q�$���4�[���ܻ����Xl��I(��a>B!ʆvZ��q�'r�g�I�K92�7O#�^��N?�cΩe��n�|A&�����_iӎ���ɲ
T����\���ϑo��[w��Tʧ�^��F`������k�W��P��T�S����Ɓ[��y;B�"/��:� �Dhxri�CU�r|��<��N!�̥,�9S���,��dj�~�+���_�5G7Y�_H�:<��8X>���B3��x�v�-z�Fac�9�2|�?���c�����L��<��#m`x�-������`�?��"/	��Ǐ/+�4�8�-98�WZO���i�M��_7A-�V{~�L6�2-Ђ�⨂��3�d;��skT��!Q�{��<�+̍U]�2���9%G�=m�T�b�楒���� ��}Pۀq�	�Q#�cbCWcȡC��qZ���և�E��۴2i���~��R�geF����`��3�?����c
������5�<r�U�l�6˔�}����p��d�B�J�J:�d�	t��Ipa�炀sYF�<R����n#}��=?���&}��G����b����n���1��鐋0��!%������_��lL-$*h���?�F}�<���L=P����u�3d]���
i<Ъ�89��Q���;J���_vL�nu}9f��W�9�W�k�F�tyz��q���;/��ȵlxEDS��t����Sw�w6�h���;���n��LV`0,��AbS�q�f�Ʌ|�ç�r�,��l2N��V��R�jC��_�	�#���@��?��!�)Y�8�t��eAo�6� ���=���>�3_�譲^�o��Fe9��u�������;�u��p�iz`�-1{��~$�D֜:�Jp�xU�o��\���}umM�@{U� Sr�u+�e�-+@Vq�˥��*�?��@�q��	�-��mTʯ��j������׍�2��/`����G��9������|g�����J���Bk���^���w-!�B�E��I:S@��?��F H�޲x�v�%����;޼�h:�hIf����a3�Si�Xۮ��Y!��8ғu�+Eθ�E���ӹ:(���X30���C��p,�DE�_xԒ8Ԉs��Fµ��z|��u����1�4&�=4[�^S�r�Ȍe�[x��R��J^�|�0F1va�`�ČA$1�z}D'�Ζ)Ho�7�j<~G����54A�X�#���^���"b+�{�8Jb%O�-*_ I�F�&a'��^���JL��Kh2�XR�{�����H�ݔ�b����x�����-�8���ө?�ʨgB�@<����W�ִ��WU���%Y��Wp��R���3Z}#�;�̼�Q����	K�;h��������R7Q#Y|�H�UC�-gr �N��!��0À��^������`�Z�A�/{�CL�ŝH�a��IFg��ܽ2U���;}&Lm�|МP*	�Y�0b���|h=��BP��(��mV�Yr}T\����5�Xd�]��:'v��[E�lzь����%�v<o)x�o�Μ��I��p�7�:	P���d��ͅ��I�X�+ю��ڄȕ�@��6������RX|�aN�A���×���.ͥ��p��qJ���0)��kE$+	�>Z6#�i'<4��pBI���t��-�0�5V.��jE�!��Rj�]3;\� $Ti�[�>��+����
J��oh���Ⱥ�����C9�9��>n�0X�C�#��}V`��)*z��'����:m���a~4fi��o�%M��������<dw:7O�� k�������|Q��h�lwK7:
(�����(���'�K�x/�Z��W���hU�T��6�K!'.|�80�@�b�F��V��@��n���Ў�e}H������ʱ�Ga����������s[��N$Jy��;.�;�B�.�CF�x4w�L�������� *�8O�P��L��Om��#����e��& �!:ڤ}�'nYM*�x���1�)x�i�\�HA��S�4���� �_\�A� :��=
K+/@V�B��Ô?��h�9�+�w�"̵��D��U/�mׂ�gʺ�bP�1���z�Sj,`T=?�Ds\0Y<��e�T�b �����VBl�qłn\�6uu���Q�E�1³d�6R���B�k��Q���������?���8|ɬ7z-�i�Ȕ
�`�o���Gtaz�-���_�b�][񱑑�4t�*6%���xI�����˕&؛7����JR  ����CX��WƂ`\D�8�>{���P�IzU�2�E�?N����F`��uK�ͦ������|���Z��I�I�F)�Xe֛�Ӥ[x���-z7��1Y�1#�'k��-w47�)���"�!��]l�v���S�Y3*!#�M�݁d����h<� �J3�ܗN\� <"�
fx	��u�'����=���F|�:�yS@�[ϜN,6(N#t�'	���_�t���S�/�e#i�e�ّ�.i��m౒�Dk�ȹ���'30:Iٕ��S���[LT�{�3sE�>vT�n�w,!�^�a�VKt���&��l�����lRLQ*�� T��+�c��sVQ
)������������_�U~�/?���U��;�:��>�v��I֩O��.ʏ]�~n4�_�ﵷ'��
�J}�M�m�� ��Ƥ�3��9*�~рA�g/�?�A)�{��Q�*_�oIG贾��sU�s��d:5���p�~1|�c���"�������ܑ�'ħ��@�#�1E4'ȕ���{�����pcp)�1)��{���?3��������]Z;��♁��#H)6��)0&*����gjVg��a��nL܌�D}����s.V5Ff2��v���r98���Wi��X2��PG7��\��a�@l?����c�����@'� U:9�a��`�Gׄv����Z�j��0�;}��D!�2P/�0��Y�ĵU����&���5�\��J���]�J�>|g�1�~�<���+sY��IC�X�=��/�#�)�Mqz�߭_�F+�N}~��}���?G���㮦O�NIs����u����C�@)Ӱ&S�:�3���+Lp��_r<�~^��\��U8d��y��1f�ҕ�	���Z=�i���-F���"��߹=�=KE���넴Lq\C�jL�L�Tqg����s�t%ߘǓԟ��^b6�~F`�c� ��1%"�� E��%��=����y�F��b+�G���^�������=��h���U<8mAל��0�%X	�3�|�V��A��L�'�Ԇ���.�*
���nSL �v�Iy� F�H�W�4JQ]���l��Ǿ���ф���*]�������K���ۋ�����a��a}�"��?}1���(��[i{��'�[��;@d WO	wz�C�+?��.��
\��#�O�7{�* �#�Q���i�/&����%�WE.��?y!��n��ÍI����CEﶲ
v�!5	2X@N츸��~>ɉ�/i��)
�_Y�:F��M�nO�m-�'M���D)��3	g�����D?�a�/�,�4%/�i*���k�h�����h�"d���"�P�c-~TH����ZRc�$�LTpû�"�R�3�׋Z�n^��W��������4�۵�g��r�OF]F0��H��O��iG�1�zQ�`���w���J�*0�}P�=/J��de`}����ȫ��[���v���z)/+bƈ��IIu��I}���3��L�_�p���_��P�@���o��۠S�Ө���&�̤�{V	�K"�e L�����B=O���7�\aICR0Y�6� �$�:��%Es�����2���t����C�/p��KL�[2j!K.�n	�l��+�->���~$�N��[l���é��$��VzwV�T.��l(�0F��-�HW[�`�$"ȍA�A*�T���e����4�ƺʩ&�
�`�SE�#��l�R��aVnӤ�tQMӬ;�ը[��K*#x���� \Sl�ƕ��|P�`��Ej5�V���&-��(� �G��	��w_?�C+���o����l�l$�aB��� !m�3������.I%!��ͥ�gk��P�K��eaVl�PDCKV%*(�k����,�ҽ*(��(��lmt!���L����U�~ULX�\כӲ���DP��OTxC��s�� ֪&x�6M-���;�پ4��t�0���4{V��_�?p[�]�x
}N�R���	�Z����5���$���Z�n������§M�}���^��ԡ�O-�����d���Cw&f�av����n���>���~%i�wse�u�)o6�3��HB�4-Q"���A�)k�N��NG��P����	�dj�ي\f<��P!��x�^�SW���u�ܚ6�H�]�c��N*��V{]��إ��
���Lc��
V_���(��E�}Ѡ��T��A�C�g��c�7��(<���4� VO�ÍI�$�d*}��L����/P(SM�ydk5#j�x�:D����g$z�Pɧ��/���k7�h�t.�l�`��=��SCL�cu���M��!&�ny��B����4}��Zn܊�� :Lsw�V�fQD�·�|gjl��!2�זjܭ��b��h�����z�l�y���/�2�N��%7d�Χ!��_�ܴ��#:��-��hPb���N����|����Bּ�%��O�}
�����iTn�o9����RiU�g�RL���<h�q�x$]�����_�5S���/�E?iVR�Z55؜F����,�ίݦ�̍�q�6�bB�nB,��@��1/y���:@�\��o+w�܃ɓ1a��dh�(��ΖΖ��W����,�9�ͭ�RX�g�#�|�h^s�J�5,�hJA�Yb���������2�PA63ԙP�� k
қg�5�f�g
��V8j���蚻�n�;��ߣ�\$3�T	��l0��]�3}+�t��T�!fY�� C8� ��t�V2y>�!Y���4�Lh����� �Cu��^W�K{��鈴�i�|�f��U�9�ſ�=G��Ό�$ϥK(�+	\��Ck��˷x)���"^�/��i�jE~д
Rw���+���xFFԵe��}����8aERG�\��>cҷ���G�W�����🜢����t	�\W�1�[�3� �!��+�r��2S�r�Ϫ���Z�;^�LK�`��[]P�rl�\�e��h��������I���X��Ț�P�k��iZw��.���<�X^HE�� ��M��#R�s}� _�G��݇<�3O�őu���k�Z�wcp����M��r���g��X^�_�pp;���q�p�F�����+�.6�{7*�[av�Y|�3S\+��H��0,�sק<+���e�(�	���=��.Y�96���:���BmS����m@ћ83�S�b�7(���x�&��X�2K�+��9����vc֓�?Nɳb]�ɸ!�� �6=�:�v��>�gM���v� ������yG�H(�xSkk����юf{�������EƜPs�t���-M��	�6O��8z�����*�X�IN3���}}��+�&L�$�X6�q���/��Ѯ!��]���%<���8)<����ݳ�@��k���ώŶ�P�	^1{�5}�{�Q����r���_�@�po�͚��E�����<��n�b��"_,�@Ɂy�b�W���Z��J�
 �~�z���W�n'��%3*�1Z�:9?G���de������ �WĬ2&rid��E���5��b�rb�*�G�:hNj�AV؉�X����CxyO�E.en��ڧ�����G��ٚ
D��dBTQJ1=�3mZ��!�S�/���i^�p#� .� hH���j��9	�T��6|�����1xC���=�� Ѝ;��
!A���/����#�8O��Ě?%�WNX�HP��J ������<V�`��S`1n�`��p8{�%|.u�d�˕���@�n�w�����ɱ>/���HyJ���k"������M�RW|���q��\2*���5������湷9���B��u����z��S7��K/w_/p�?�,���Ť4&�zP3�!�?+p3C��zN\3��:�K�I�������u��%"5@t���X�?���.�r^��KT����>\���mD�ÅK��BD�Z�l_��/3o�2���ս�g�ք=^��+bp,���O����n�-��O������sW���A �����X�B��R����He��X>r`�.����A���f@�Z��c��iy�0f/�MQD��62�9�.��o|��U�1��c�d@���c�l��Y��.a?4~a�N���.#)����4x�S�0 �0)獹���I�4���;}2%���"�첲+�l�sq������$E�FT�u`�z'
����l�4j���a��J�n1e	 r%.Ƥ�����`�O�o)�!�D̭n���!�6�B*�D��"�Wr�����7e� H���l���FcOs@�i}c�1�Q���j
��!��^ʩ�(@�Gـ*<� j����p�=�X(斵�J<��8�G*�"�0i"O"� ���U�?��䰿pmcVÜ"Rx�J����w!�)���0/��@�{�{�K�E�{=T�����Hх'1&G>�4P.H��3[�A*�
�?Ѥ�51�q'd5(�I<��g�S��$7TT�OQ�]{Gڙ4tÑ}�/A)f9 ��dd��Lf�sxl��2ھ��v��f��8�Ŀ�h�f����9�D�*K�6=a�tG���M~�N�}�w����&`8��|ޝd;(�I�)�l��Uu���=��F����+�́z��{#P�ڹ�g��3�N���'���C�kJ/��Ż�������^�ر�(2�VV��ՊYڵ	�+73��hڲ�3�91��ϴ�
�<�i�.5aBqE{1e��mg��V}x���=�y[[[x��X�G6�����:��n�n��3��r;��HJQ	u�i��6'�ja�	G� [��w�<~+�@\�!�q�m��L�Z�@�G�x�-W��x�%wԜ=,銣�����&yK��w�@��Կ0±i�[��v�(�G���e	�I��у|�]\Sh�:���"���N��?3x/Y7�R���Ͳ�Z� d��ѷ�0 U��B�Ke���|����U?l����}Y�#�-��|�q��h��&�i�%�"��(h]}��meF�q��H"�3Tm&�K���Pc���W%��	(���a��-'�'L�`�~����ge���v������C�ed�Mc�=��i�p�]��T_�b:k�H��R�����P�ip���Y==�O�6>�L�u�R�/�_�ސK�w�?�`(�S���g	���fk�Q��O�נ/�mp��<�c�n����@�p��B=9)7�$�PE����Z ����AoA�7��l��Y�TI�I_��G.:3�̧R��[[�N���C��a]�57��Ud�>RP�ō��,١�d�H��U֢�GBI�Z����R|�����z������;A3�C�hz����S{>�7^��cyU�<C��]���sT*�9��Q��H�:e�L�XMު@�/�37�M�A����C����F�0�0(�'R��{9���'���t�u?qM�s�L:�J>k�5��Ɩ��j�%Eߘ�ggka�?�&V����Ij��4&z� ��Or݅2^�;���1&B��yr~af"�^�����ǡ�C/��l�.r�w�����N	>�ai~�r��G����-gĵr������ Sn<��X��M/��5�>\��H��i�i�up��I/�F/y�1I�_iw@��
^7���.w�"�@�o�羴���M�	�H��#�\����8�$d���H�6,��r��'�H�fN=i?�ק�3>� !>x��� 1r̬TpVf��5��{TJ���j�s�.��Ƽ=6z�ߵ�w}
U�;��)�7���B�?�y��+�]�W�0{���T�5�Nԏ_h�0��W
�#M��<���׬]�	e	��񺶩{`���u���A���G��MkZw�[�5?�pŪ��e�����^b���	m�۪�3A��J+	�� 4�G҇�R!�a+m3�9:o�T��
��5*�1��:H�P��S���-.�z��=�2f��B���o�����_=	c �Â��J�8?���i�Z�y�*V����ti�oVw\��[�$*�-��MyIS�' z�:q1���&����"�����o[���4��^%	X<��D��aiZM��a�QD�+��lQ����DN+"N�A� x��Lν��%�6�ϳ�H�$���+kAݲ|���7�1� Zl�'4�n��0��
f}��Nw`\����@����г��=�#bu�`?��o>P,f�&��^�=h^O�:]�iHUK�U5��"����cd�\�5�mZ�����Al�w7�(��=H�=�/52C��xWN�%��_�߾�s����+���I�af��J��l��M�]Ry��zmޓ������M���,���n�Pv�������dd-ca���	|ѡU�H��<!�'��2vh��^K:t���,�a����\���i���F�'��5ٸ�g���S�$�Z�7�b�B��c�R�;3S7%}V���|p��o�4\wq� �1���?�g�
�c��������@�m���Qɑ��=��%�3?���
2r�( W͸�*?C��ox@I�z�]�s����`~˸�3p_��c��ឩ%��b�{\6u4C����ײ�)��N/��J��oN+�U�Yt�p��jTl��y9�&8�+����_g=&����A��|�$��æ��Zk�˼��� qA�1l{k�[��xJj4쀜�Wu~mD�:���f$��v��GoLL����0�J`�y�z0#څIv�^�hf�K�~�ɪ}`&>g����^b�|�[�c����:���e�P1��I�����Ѧ,��Ћ�7��ˢÓ�
f.�+:e�X�
���5 ���& ���|����Ȇ�)Z r����>�_�i�x:��b�6����K)~���O{[!������cQOM����?2����c[U2K�a����� ���B��w�-�`�#�1$}l�0�����h/�#7��5z�:u��[���ϋ�Nr��N����B*kb^YRd|beY�c,�<�����'��2-7؜h:����KG��r0����5(����P��ئ���Qb�+x����U� ����Af*̉���F�����nQ���j4��"���2��ֆ�p�z�'�,t>�}$����w%̮8�����NI.C�+I�(��K���B�*Y-ǡ����>�y���'�oؘy�T#�K�֗^@�
�<�����4z"��s[ƿ�YhT�[	&�,�xV��\�G��GŤ~\�����\�T@n�_�ƚP����r��4r�-3p�&6D`��
�x�����ޤ�|]	f�k����������$�L��h7h�KS W�k"�3nc�W����^_]�����6�v`��x���7�,��a1u��"=��pOH�Eu�ӂ�� �h!)���xr��������x=Z�#?��b�[w���V�}�\�qq�,!q��nL�V+�a�W�+P3;��'��^f�@^����dF�+ئ�:�k�{���6��Nm��&5r��"�#�jU�y�)��,&(H���,A<���s��F��c�2 �����"��6���[]ɭ&�s��uVp�C�AY;AT�+��Ҟ����E����&���^�V6Ϧ��v,��p��1c�	N����wDR&��Yɜ�E���V�~k�0�͂k�a_rHFܐj��6��Ut7B����Uu+����+��l��9ܽL�g	�6m��ꭆEj�0�:�~@�m}K�t'�*�u���O�!3�+n+���N �e��0XJdYg��2���Bc�Eu̓ݷ�"W{&�&W�e�܃KIo������T�)�g��3���D!�����7AloD\tV�S�E��
����T#�{~��:��yN?,�1(�ޙ����!ۊolw��lO���ª6O�lv�Ş�c���t�,x��lD�7����~%������~+��6����%�¨n>�w�x=_y�66 "p�Z{�)��yE55"Ȓ�E)GA_�>µ�T!�a*��U�5t�Y�XI�����>�Nh	P����`J��^��&����V������vG��9�"�����?-a||&�f���EpRL�H%�7{��>�%4�)� �p��uG��Vcݹ�1>in<��m�<�߁OT���f��b�C�z��u7p�Q��g���_r���ltg���`K"��D�l� �گ"p��ݬ�
�BR�ě�˚��\�EV�2#�?��b�\��. �=s���l=�d�}�K���om�������vT�6��|;�_߉��ձ�ķ 7_;���DKJssg�K?��@r�֓�@�+�0��AV��t�Z�-�*�u���8��+�O�)"�V��+I�����:�0c��z��_JTi�@Q�)/��lj�45 J���/B۹�px���Ht'���4oOZF���M_MCB3�}1^���TU;�U;�h�G�Q~\Hd�� T�B��>�>�ngѻ�Oz�䴗��t-3��?�~���Ϙ�|�gD��}ϴ����r�B���*��;�Js1�ƭ�6�$C��Y8��<d���� i�)��ٖ�&���6-�K��
���X��5Q��	����@��gݓM��ѩ���=x����Mx+�\�z0�e�+�н���O�F��$,ͦ���M��S����^�8�e���z'q���M��Ԇ�@�˜g,:�t���sSN߼Ψ	e���En>�a��*L��)��rR[TY�����j���0�
�FL�������F �2�����k>l-��C:��ʤI~`�y��"��-�ޓ�y�$���}��Z	i��O�`!������B��}��.@B*OzY�[WBa�Λ�LĽ�e�b>}��g��G� R��!�	�X���v��̸-��#�H�Q��5�`��J�W�h�A`c�ч�]������	K��/����H*KT,��D�=Z������.c��1 qX������k�Zo����q�	j���T/w޸�0&�a]�6L�r�}޼�ڇ��{ePN�x���Ք0U[��4HME��E�d%A2�6؋L�r����vԖ�!* k�d���HҺ���g�Y�~ww^X��| ��d��ƒJv�#�<�[���`��3/�5�<��	�t��'�@�7����1�1�=�L��f?��ܚʝ�[�a������4�;�*����H(��Ǥ�]�J�j��ԓ���ڋ��s��g�tYL���ˇ:��yo���Y,1���,�l��X�MJTtO�$FS��(1nF���=�i@~�oۧ�%7��%Q��gM�H%0�|����-�{J�S�F�y����g���B�KAS��fA�#ʈa��4D�t���B�ޒ�1�i)��g��l>_��Ă�p\� ��S���-����&�|4������N���	�,� ��A�2ir`�ha��M#KLX�hN���d-H�������->U<��=O"X����R��a_��{��qB��C -�'������=��x:?y�u��GZ���>��~y�P"��z2�Ne�%�$�d2_��?]vN8i�hRurU����\�|��{�!��k*�:�ה\-���?fJݭ(����׊l�ŝY�k Д
��N���CMR�v���B��O��{���0s�7;D����)�����컽1E�
�c�U�3x>l؆��g_�A��$�2�S�BCP����+n�%5l�����C�R '�h/�a�j����a�puU ��)c�)�=���U��Xp��&r�#g�^�~��x�+$��(L�X��O�q�bz��*=��$�=C[�4I��GQt�g�mZbdɟH%F���İ4	Z���]1�=����;V���{�Sv��[�w���S���|b	=� A����Gh�}��ѧ��p�_L�nC{c�n╶Q#�\��傆�c��i��7��*�)s���k�O���e�W�`�6�97��~�[���NͲ��o�.Y�RY��,�'×�����{� sN	��v���P��"c+_IӚ8��\��:��a+(�<T��������'����bL<��<o��J���,�3��c�SO?���{2q|}>�d 85�ֿpz�g���̪�2��-�A}�u�<�20s�b^����BeF����LS����ݜ�ᖺ��[JO�������5��ll����<���)�ܗ�!(��s-��4�S� �H��z��IPb�0-B
�$���hNf,S,�ų�&*�c�P��J�Eǔ��0�k���P��?�b_�G��&�r#NE���ʞ�p��~�RR����RϢV��&�ܜ.�3��-��/�Tc��zl?��R�a$Ϫ^.���H�v�5�}�`�;�(z��G*v}���=�j?a����ig�%J&>�:�^��ssR��Z�m-'�݋�6�_��n��cS�WI�U��$��PO*�SF$�[�*�7F�;�$H�-ƧuLvjO�x�'֤+2v�"���h*	V�D��@r`�0<�P�g%��ӿ%�h`U3���!��3+�Nr9Yu�x	�(��`5� _;�� ����x�b�4cZ5��d([�V��N�/� q�>������0�P��}��F�K_�/y��gr��� -��.�]������h�l�I>̩��̷/�r�x��~���v���u�͆�)� ^���]
���_����#�L�Y<��7^D�h�/G�}�n���#�6^����ش�C��7˂Ub>%���%����'/���s�wT���ۧ��w]�dMIT��X��ڴO�
f��_���*J�����z}ןUЈ�>t��*����&_!u�����{�7��8�*L�-\(�!��Y f�	��;9�'�o�{2Kr6���&�w5��gf����}m+�I@��ϥ&�zF�����t�����}�$<���k�N��d#g`�$)��-9�>��nS=3=�G�(�[��,�`���3�Y�]Jʋ�V�kG��6�5M���S��W���ݽ��5b�ؔb����]n����t������;l�̟W|5��>M�-oz���-�Of-�X'�&!<3�Uf��j�Z��m��1�ɳ�Da�m8��(��2�U����5+��JX	xf�ǭ��KBi��S/���yh��r5?��P чT{���C��ߘ�N��&$����e���-C���K�i���[>�X���W�C�e0#�|�G�
��T�	#ڨ@G��l��A�p>Oޝί��R/!0\��z[" 	�7F��:{�uv�����;�Q�h�LWw4C��9�j{B����{���3��aMU9\���8Tjry��z��fK?��'P� ��ڴ�Ȟ�<��<f��v�e7�U�$�@T��q>x��Qn���~t�}�-�$�A�vXT��x%�p�C��h��PT�>�O�%��1�J���,�]�-�!��2���sN|��S:l�Ig� ;ԝ��\Rp�֤�X�/�蕪��6gUTz���gj�R&^�ҨH���=�nu�-�7=U�hTD	r
t+<��K�g����d��K���:z;[�Q�E�[s�f	��s�iGU�t�㲠d�����N����>�W��r�P�<r��3O�q��R�>267<��%�P��q�YQ쪉�\$G�mӂ�	.&o#N�[�fU!gF��jD�"����0K�[Z�ܱ�o��G!
��6�ŧv�cX��T)�'��@�02�M�9U�FK�O/uM y%�1;Yjsg��c�y��ֈ�
%��ņ�i�������By=?�� D?��hƒ����r�݀���Zs0��_0^ƚI!���k��u�Vqao��d�`��ڐ���H���o���XiPpd���Uc��9>����uc'A���	��MvhMT�2���bHx27�Њ7�:RrZ�ا�)�ʸC�W�1�Ժ�����ӟ�"I��?<���"�5u!P�L����H#�`#ӓg3��S��ϥ �e�J	�����'�:=��:.�H1K��^r���3FԌ��O3^�e���j?��6��>U���%[��sE/�b�-���yYz�8R��{���Nm��=��X,b�%�/����T��̻�<�5q���ե]�9���W�S?�T0J�,�Q������1��3���}Gi`�e&[^�%]���q�,�ٶ՗�Vk����X�g�G��[|�J�	�f��eV�������~8x�ʤ�n��� �g���i43<���=�X�%���x�$Nm-��>�2���f�vC�P���I�o����Z���r,�S��
7����M�F*�����^�*��%e�$�tL���I^�8`CD �ط>����B��Ǿx�Nt���Z�����2ޙ-YH��O��l5|�@��%�*�lM�y�ڔYT����X���O�@,�c�5s<")�
3G�n������8Z��A���mp;z�}(���H�t47��'�"A����S�TQѠ���-/p���J���V�j�F.����,/c�B��,�|��h�S8�՝ǾnԬ� �s7����M�,$e�n[J�]�g�����Cv�Akv6��ز�բ����t�?�٠$���8w��Ĉ����g�;`���ݑ���IfKg��F��'b��͔��H���t��n��*�W�	ɋ4�1����������Y@@=8��lt�ڭ�����	��E�TVE��TC�H��v%Ve�3۽äpH�a����a9�Ҽ%}FLy�"������K���_w�?��;���[����f��{�p���]^�v�6�Ȑ�(zz�r��H,_S�<˓y�v�Y���'s�Y��繝�*]M�WeY�U����5�Cg�	�c7
g[�[;9+g�e�fP����d�� �]�J����L9�L�C�C�6�R�n׋�aU��Ok �z��t����R���d���z5f��� �\��'��d�2��}؆��:ݜ̐��W�g��G؎bw�8�$j+a�*���A�_{�老	�C��
m����`\Y=`]Zi{�\O��=�lL.`F܊�,������� ��@m�5��u÷~#�=�K��턡�ٶ��12��h�=�Q>�:�!��'��q�x����u�T��Gh�
���)��OLO���4z_�^�F����0�F�@k���2�+(':�*L�z�*kƃ����yMV/g�]pX���K�}mM�S��u��[2�����)B�t�j��B]��(���?O� h؝�>�j�T�1}�2*�f#�𾕉�Mu�,F�^��L�򐯧u,�%���7�H�B����ic��]2�yӃ���������6l{gqZZ(�-U7h�[�P ��i�`*H�NE���~�7;��g�牅���^L+�x_��X,ߠLF�O;��b��~+�7�A��.%��O���
�6`��������
�m�v���9 =��Դ��}E� vđa�b�T�	E��O��B��;����6Z��ᕘ���T��䡘ɤ޺u�r�� � du���������d�ODx!V2���أ�h����\�*�	K�.ӳO��c2���2}Q2{��mM]�'^*�-jR�'�����*B�8l�{L���(|I��w�����I\x`{�X��aXE1�]6��ɮ�Q��Wm��� ���攼������(�tn���I�2�F?:��a�[��������x2>��Lg�ګ��A�G쯰�cq7��:����V�P��]n�烸}?Dܷ��>/�M�~Y�� �@��*� (p��F���q��#5̲ �P��u���wn8�w��p۵')@���;�¤ e��ΆvR.[[#��쓀#!?�"!���:?���S�h#�s����:�|s���9��HW
-����7�am�eX��Ŀ�#j����P�V_��h�K�\W���\�T1�&yB�q+�� �vB\�.���u�yB����uf�mp�����eq�E�&�Ny��� �vؚ�żn�)U$h�`9�N5���uB�M�<΍������5�h��1c4��]�*�cΤ��\��"����bm����#o����"�wF��Y�n�!��������p&��L�P~R�4��sWI�<�ҝ��]*q��q|�L|���6�n}��N � 8։
y���u:�M{ܻ�.ʫ�~\&a����`}]4��'� �?S��:��A�s�����GRr����h:�>?~�;��;��7K�`�/