��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0���C	�i��E�~u���Dc���
�#�X�y�M$����<˳2n˾�)�X�pG�J�Ę�|�3V>@�u+ǡ�ўQ�� �"���!��I P�L;-��\(a`��
�[ �+��^���ш^˝BC͑e"��eSjQ�G�9�#���Ul�,������[B��fڥ'�d;�՗�j�F,��z�uġ���:�&�2u�(�1 � Ұ���uutj���sp+:m�/�6gܚ���O;�{(P�V��ȅd�bR(�b?Z/}^}\"!��%�/����������1N�&U�*�x)�b�{[��4�늣����WJ!p�a]N���3���|���Y3��6f|�рʢt]��ZO��oR]%������įГ���j�	e1l����+	��p�tK_�������GH$DC��U��[L[L�6$�<y�O���Ox���m ���C����y{UK����=k#/)-��O��������&��w�.p�5	�V��lf�.��� �d��G{v����3ۈ����&�m�����C�K#�[�5L�R/�! d��^��Bsu[����h��	�}��{$L1	8��.B�pe~�S�/)`�^&q�l�d��[ �k�#5(���¦��+s(�+ym�5�.�o���f���?���A���1��6ҡ}L,��z�e=�%\1�Wp��M�ī�����{��A@i(M�:����ZH��73=��!�=��[�þ��~r��OzM ��	ѯO�?vQO����-	��>��Fb,��F9q��L�����MZ�)0���$p)k}QR����z����OGʙC낃����Ib3����7���W�bsO/	@<�;�[��Њ�Ϗ����㽸�aU�b��#6D�A�;o���oF�[ѝu~h/t�M�ڸ��J��y�:����i*����}4]ih6qd<Ҥ=�5.-G��,*��4�z����M*L�# ��%DOSp�}+^�k��k�ArpP0Y-ZO{���h�z9jlFP��NT�Kd�^td���5�����ʱ��9��I��W�La���*-n��b��A������!�1R������o��^�ȩ'Ij�!�G����\���8f��Z�'�s�^�Չ�<>��χ�Wq(y=5�����&���k}����+�ֆ�:�f������
��B�0�6k�[,�5-�L��W���V�x���N�l�9��t�]��������x�����Llùp�q����i��Z�����=��A<�;�81��e��*��o0&�?�6���A�բg^���6���'���p��� �O��a���]=�}:Tx�y�r�nف�������W6.���1�"²�~��%.��,�:�;s@����Uش�7�[�0�:GU_�P���(��(��~�9���~���� �l���5�������S��̜�P\\];��C�f��/�x2EnK[9�b"�B�3ܘ㨈0 ̇�qlS��
��{b'Lj��6]_P��������r��i�~D�|�ǲQ=j5#��b���K��A�m,(����o�5�(�|����I˞���Ph�ϭ$�ׄ~ٶz��t���N��zR�[��)L�;n�,9��c����U��8̏��˧u��
w��T���6#Ю^�F���ўwts��6P��]���\@�M���J��ɔ�@�0ĳ��;���d��W�׉��u[�\�[�@�3���@fS�ǵ�L}N��![�-)�O�Ǘn�Z(ʕp����oqX��SB�k�F§F}�IyOx�Cz!8j�qO3�yAȩ�eu �����\i�*-����ZnD�B��2 ��n�Y�\R�˶޿~&&��^�=�����L���S"I@s|��� ��0�S|�$JLo- �:��ዹ���۬�_�;)��Zr2��2d� ��x�U��c#c!�#i
<�Q�i���L�|Uj&ڙ~�~E-`���
�&��X�U�+�B[��VjC0�.>�����YAj�9���.��Ar
TO��e�s�ͱj�����⢩=�����$�Y#KO�ß��N{F�!�=�[����o�Az�t�؇���/�t��'�@�&��]�� ��:B�~ �j�:5�֚x�2�4f8'W�~�;5t����l:�/��o�����[�KkSq�T�4�r�ڍA�fBz(�c�+
#��,�Y$֨�
ƺצ�y�	����KV����5��U���ϥ��y�_8N>I/�0���2�1��A�1�OV���h �^��4=�;u��ؒ�����IPj.���9�(���c�)�u�_��9���j<�vYk.9��ÆJ�Q�;5X�Z�u9���]LD�%�ux|�pBh4���3�w.��X�e����ra�DG��J���:�mq2YG�`��<����^�H����}�Wo�L�N��`�	D"��+}1�n��<t@*H�ܷ�o�Q^�<��P}$���U�JF�h�㽖=�ԯ)�Љ�8_N�}7z�-^�Y�4�����gڠ&2`�FT<����H����:�^k���-�S1HM�@��c���JX�bY�Q���Q{�:0L�i&�����x�pU��#�&�k	y�QT�(�~e4��=��'���.[�a?�יs���$�Vc 9)}���pw\�3z�mj������{.��D`�1-��ԕ�M;|��7���Wua��p�vѫ?�mSo{�hyn��x+�G�k��]~@m��qQ�u���$H�.�6�@���vdc��A=:��*fР���gIk��+ɹ���+|j����g���<+p��L���Px�t~$�G(����O����<�,F\�{Ft�Q r%��*�o�o؅����%J��aZNٗ�b�e��
2w�,�۾%{ru�	C�~h��%�ɋ31?� �}Q���5�I;-S��rG҃˟��4��H,4�p�F�)���DO���:�3�.�4��|��%��z��lC�*�f�)�� ��8��hnĎk-�*69i*��
�`5��#�`���/
L�k��m���t����%̼�!;�1>��1�+�s|����wl���Ձ��4@0��jT����:�Ҷ-���tb���Y%���f� Ѕ�"�)|a���E��:`�����m_aN>g�S�0�l��p	�䯖��t�x��+b��\��@��7|{0 ��A�-�ړO�۴��ӮѲ������A���j;U��^^������Bu�����Mq�M�z>�)�@X&J+H�< z�l�k�K7��n5]� �o����\%�5�Ŧ��G��V�4#-k�_j���9��������[j�������$���ŶZ���B��"Vt4pA�NX�(V��3��7�QUk�,"�"��3arEq�jN�+᫃ē76'b
�P�$���=,����Q?d�P2�Y/qiF��Yבjz�ʪ#���ٷ�!7g�8Vo��X�w�)8�O�y�$jw�>+�ZR��-�ڥ_���
���؞�� ܏^�p���V�Lfjm��e-D�`߅8��Ļ.�\�I<�z���w�vi���r�L�ت.o�� }<�Z��ߘ�ŝ5Z���ah�kʈ"ǟ�DHo�A^p���u��շ��9���m�j��#�|u��^j
�P���0�8�p��#��[�!Vc=��]��.ݗ�v��(�Y��a�I^ʤ�7̟Q�}
|Ѕ���]V-ɢ�*���B$��+�w�AU=����H�CQ�p��Å�o*ƋD'O1��K�8�ܜ�d��#n��̝ #�.�,�2���Rߔ�@���Rp�����?���sp5����	zveM�0\x��v�B[�86�xW��2��SN�q�6�:�9��dr��s�@��$��hH�"�v�p#6C��5s���ŭ@������$\ծ�8m�aHj�1��;'�&FL"�9<�{�kI�_o���#�Tެ<�,�t�`�F{p�t r�n��0�:PR'�*���J2�����hJWP�?��A��*7�ǴM@��w����йֆ��|��n��W �LH�B3�[;	����%����/������[~{�j)I�z
�@Pq�I������Qe��;��8ֺ���l�ۍ�I�p�j��ɍp��Iۄ��E#m��?��W���%\ "��5�96e���ȧϪ��8ڵ�q$��mq��!0,	@��V�	B�ݒ�I0I�zFԐ��_�`v�\!>Ob�U��7����me8�u\v!�?��S!�����W6�O��'�'9������bs�:zX�%&D���� S�g+I(�|����8���.t���|}�_���%�F<Fjgq���B��3�@m��rz��տr�4�:�$�v���˦ ރ�A+����J�&gK�T��w�����K�c��a<�\��.��k��Vm�?R��.聲�F�Pzͽ�����{���!�ïv�d��<@�k�b<"�Z���<�iv��c-�h�"���t(A�l�l{l����bt�x�K�G,�U���*"�����\�;b�-܈N��p�[�O=5&��Ļ�}�5�n�'\Y����f|�p�"�pi����+f�3�O��Z��bnH|�l,t:p��'����y��kw0W>�ױ
�+�e�����}"�嚝:#�J~�;AO�ҿ��*���fh",��Oc���č��9�D0[UdĒ�*��9*^);)y���2���s�A����=ag:� {Q� 8�+e�(g��K��oo����xq(����q�W�Muь�)�L�_���\����>y�i��`�&*�3����6؇{�sG��#�Zݱ�����}��K�x(��x�zS���N���G�~x.g����)eU��2>�}�����Њ��EBe����g�e��))^��T]�<p.�`	̄���2s,�or���� �G� e�Q�<����d^hs����bu�2"�9:Z�R�Ԩs:��#��rc-,.��[��d��� ~�Ǚ��i����X^*�ދF0�=��0�>T��"��ū����q?����5�+C�g�[&��6�oC���t(3�h�<^��#e|�Q��hs=��#������{���8E,q^��@"�OzA�I D���%���#�-����"������>�9`�(� �����d�t
����u3b�L�`-TE��O��O}��Ǣ���	���Ɍ|^uUMRwCbLv%+���< T7%ϝ�����jĿSh�ޚ��ʣ0�f��et+�GV,���&�a:�F���fY�z�aF�j�˭B�>��m��/�����0�<rd`�I`\U}