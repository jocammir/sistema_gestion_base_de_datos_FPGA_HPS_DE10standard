��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0����_���3e���ӌ,npë�;^rz� �zx��3s�%�yu�gw��Ѕ�Nͬi����PH��>W���U�[��N��2ЮK.Y�[Sx��MT�HG>n�9����}N�veǮft���"�7m��gqk����|�¡U��������D�����[�0;��%�D����(����t��>O�|��/N΋ۀ��P÷���U��������FߡCZ�X4���*���;�MJ�-sBc�z�ѫDfH6Ȇ2��[����Ȇϓ95OA��/��~��j�4���m>��x�(JǇ�D��p24�K�y��Ag�I�|���J����ȅ�}狿U̬��|�GR^�z����Jq�A�W?ۍ9�����w�"S��<����y�%��Q��V<7pW��|�Wdi�6�$�@ԏ@J^�l�w6�a�"O�@�y/��k6W?'߻���O){�x�ْ�m,bc��*�l�����8�6o�K�*�|������/�M����f�eۮ��ao=<PRGqUjb�r��z����уq���P���}��Z�?a�̕��LQΪ�lW�E�R�m�(�ӕeI�M�~��O`�F�<{�a��)5Y;����I�J��r]!�FNx���"5{��A:�������	�ɱ��t!!(���*��G^���GI����J |zI��d �BG���:���V*�7y�)+�mVe�Oh���,t�FW�t=��
�Gr�#�����c���q��iG�5�� �`o�8��ҥ��q�ԣ�:؋+���km�M�FI��f���|�tR̙��6R�u=�G�����Ǧ�uM�nfI~o�]�]M��)����B �3�~4!&���_1|��Y.�����2��[�zuZ؜��>��uN�ͧKN�Oz)ú^o�0��S�Gնh8e�ś몕qE�0tW��n�� �C`�w�t���M��j���g��@vrf�#|�凷��,�2O%ȕ��Vs��o��/1�rz�o���`���68�Wڈ�� �������H�}��HAª�:̷0$F��o]�nM��z���_c�%��uw��es\6��^v���}�S��f�j،�;�� /�\q�x����n��'���{a��4�x�F��n����bm�)�7�d|k(R��3KW:47���~nɇ��&g��Ǒ���7�=ɾ��4{-�re�>CY�bi�@^�A�šJ��|�/6S�#]=��|[V@Pz�hQ�;�� �^�G�b�4�ht w7֪�J:䪇:� Fq/!Kv:u������牕ljՍ!���-�+\k�p��{�h�y�D�i��c���A���o@��:by�J�����y�]�пW��mj�7��)��tj|�c�^��f'�)T�ī�5�An�e�P׊k
��S�TV��|X%{t�w^���b�&l|�?�>�0�|D�&`�qҨ���%S/�ȣ�& ��Y{q���Eo��������]��$�'z�/��zR�`�7Ur����0��5��%+�(C�!�zuq6NPe�΃A���O;I�d��#ni��#����!Z���h�\ט"I
�͹�N�4
��1{���t*H��ZQx�WB���j�j�ej�b�b�!�H�-Y�]YD��C,�z��l�K)dl�01�L�R��B�F��K =�P�f�[�oH�*MX����(R�y��zy�!#�Ņ!��D�!k��υ�3vh�#[,���K�Q(��w����fT�$�*{��M��O^[�
�xR!�ޏ����3����E�A	"RC��]7.Z�y�`�� ���r0s�$�Q�&�d��/8(�$ѵ�N0���R�"g�b���1+��;�j�c ](%;{s��<��z�{m�"�^���A�e��iV{�\�G�\u���&��f���d��F����|�f5X�^` �͂O=���g��.��K/���y�=��m��*����I�浆<�|�̔%����g�f�c�+�;�1D�3�&(�͐6d<�V�����p�����ս����t�$��"�=%B%�<�=H����n
�B����)�*#�I-<�G�J��k�ɐ��
�����@+�ɐ���e~�5}�պ������� �N4߉�A�QQl����!>d2��uB�����l`����>0r����o7�
�G�eB1��Be���z2���M�0�Ш�+����pZ�REy���A�t��:�l�4�RU�G�'���Kb�m��=�������vN����Uj��-w��P�`�U�����*(WI�T�-x�z�8w$}3
3
�� A\w�j���#�р4�Y��l��7d�(������c��xο�|-ec=�<"�y}�M��x�ɠ�Mϙ���E�].b�N� i��߄��
pB��Kv�=�1<1RW�-�6S���M����cK|h����B3�C:���}t�ܥ���o6���]���flo��ߣ�F7����j��8�/��t������
�|��SR�hK����K��RT�57��t�d�[��:c��`n&�h#�w�F`�3*)�'�Y��<p�oEbހ��� ZKhZf��Q���GrX0.l/J�����^��?d�/}#{̜���}�xrM(Ue�荼�L8��ї�Jd��zm�/�^NRR�昆��&*�Ō���r��Efc�t<�Y�J�<z�zy��*�����5I�7Q��k�DG��#��ͯ�`�&���8��Ոl>�!D�!���)�ᅃ�>���|]��O^
�_ `3��yܿ�6V���E<'������
�νG��Ϲ�JG�鹠_ ��i��l>�¹&`��&Ū8��|��C�؏����yQ�Ww^�LN���2 v�W�K��S�M������{K�s�hT�3:��� 3����%|r�.�=A<� ��O�[A��[S������9�l���]0u�M~���Ь+�r3ۄ�do�P_�D�8���Fg�N��J����m��h~�R*�4�����s�!�4 C>���NH��bV�dj��6�u�o�eN�j?����:�������ٱc��ԲR0}�^���h�n$���#���P���AvD�͌�	_�O(r�<��Qx��m=-�J,�vU�6��nܡ����^~�m���&4%ԇ����F�I%�H�F({ �7�=~R��I@���4V��3��K8��p��DpL��]y��l�qk^u�\58�1�lq����y3ڧ�4�r,�<Z��;�G4|'ΡW��8m�x��0(\g }ݛ�{��{�a	��"`]�	���L}����EQ�t�^�L�&~�h� �����%g"m>A�~)�Ɲ�����Y ����Ρ��ҾZ$u`q;hXiF����U�8�v
�)İ�I�y�|��X8`�t�$f���g��ބ���rB��ɞ�Y��!#�}�O�?�g�U���=���1T��(ܘn[	��a�}�<�wPiHoF [.Sݣ�dL����$�'	��JbJ��8���6仫�������rA����R߰W�>z�X�H��3��p}au��%�����5��T�&�=���f��H��)������O����B#��ܨ@�ߍ"��N��=�w�>چ`���HM��iW�3�Rb��u�	y y�4K��d����F}�ϋjy�/ҕ����?�ԅW��_���N��g���/�#i�6�dZid��b�+�ɥ��x��{�����`K�
n� ӹqg��Y 
�����2ؕ�1�,zG|&�KYo[8�*8C�e���u��.M.y{w`V��~��Jq��0�/�j�f��qh�� tǥ��U��H,��� �N��p!�����0ՀeÙ����D��v����!�M����T␋^S��]��t�]%��:�}��ܝl��QUf�w� �r<�a��7�}�'�<���j��䫼3V�T|�������\x/�kg�W��7\d���K4�?s�!ۅ�������1����_rȯ*��K�Q����g�%)��Gm������[򪪪s&���YT�g�N�=�"y��{y���]y��v
��$$��/[Ҽ��/C��!F� B̪�s�*Kv}��'��󲘏�����'�,�B[dXP��~ﴘ�������]ř��-X
���D����m@���-�!���4ia�����n�@�y�=b��Yg�$X/@k�oG��;c��Na��<�Lj$+��n�{�[�G�M}�5��̗c�J���1����ѽnK�$��٭s
���G��+GD�g-�
����O2j�Hҷ'�0~׎!l<T��E��I�uA�����������>�ܝ溩�M4p9P�n��'�x���zN�x~u�?�!@ ��uS~y�:���P���uq?�_�����QH'+��(/2����������a�
(>��Q��n^���gj�� =t`M�=|Ծ7�!�)}�顧U�	�ꡛ���Fw{�`miJƏ�!�.���t�P��'�u�Z����4����Y�A�f8������L.��mWG���@������DXrr�M���:'� ׯ�-�S��H �^����V�+�7��C@V�
 ��C-��]ߢ:�*J[V�)ÙC�^�Kň�V���a��Ѯ������1�(=	v)� {��,���c��
Y�+v};÷�}�!���h4_c�?��"�^�ʿ&k�=Y@��;�wn�oR�_Ydj���v���y��Co'Ii�̘c):^Z�+�A��N9���Ŗ�m�E_u���:�nnjz9bM�x2W�����5��?�:.r���c\�bO�8����T=�Q���ϏD��-f�|�J-a�"�ɘ�.��N��`cԶ��:,��P����(�f��E��RcI6.c8�/��'����[�q.x�m�-n��,�tDI��'��	-Wj��ԛ_6����ď����R���;L��k�p!�W�Ra��2{���X\�S�Ǒ#��Ԟ(�o���]��
iJ:[1u�7A!�poB���Ve�"��^ӯ`0%p�0p�'"4�{\�$y���N�·M��3)՛;�+�%<˪��'[�ٍ����;��_R�掋�{7�7OW�wd�n^��?A�w���J�<NA�j~aRv�i����[:���L�HY~�x���-DY�4�A��>\]Z�F���S*�d��c�I�=5~_�e[�
�/���C�~�>Bm0sb�9���%�k�~2\�|�����Rm:��v�2ȕ }�K#.;vYAL}�&��ZZ���׭�cl�m�I�T�MEa�B���ݪ`������|��+� ��^J���V��,$�kuߑ�5/��vn�,�IX���0��V��8�����'���%<6�maW����0H�y��I����� ��T\��zJ�����p {�{]Y�P��Y�^�ݜ��z�`j�؉��Y�v���	���w[쨳$?wi��U���RM�Mu0�%���m���Hs�TQ��"����Ip�O�)�i	s��iJ<-{��U}�z��o�3�lR�@֎ T������vQ7�]��ߒ`��Ƚֻ2I����oq��߼Ԇ~yD1H���/��QY�;��l�e������{K�"��� �Ǫ��qd ��x���2'�{xZ��.hϓ�6ˋ~��P��U�F����b{`���Ga�)��4F�|�!�N_Kڧ�g\`Ә�-�eU��_���Z/;6�$�6N��c�1�F��mA_�@(h]����R���W�^��Yo���=C�y�/F�0&��}�X����.��_�r�P�?� ��uyj�f�1_b���Hm�"��>~�A�������ޫ�K�����z�w�$)���p�@�R!��'1�����HSE�!�����Bе�f���ɟ�Q%�
����s.b� 
��z޶�a�`�c@)[\��[�Gs3+�Z�������4'J�j�M6s����~��g��Y�����Q�l�w���~�7�"�/�6T�L�%@��s�9Im�?uq����e ������O���q��䗘���J:�]1�O~!����O�ٴ��R��V|;=��^��9-��Y��˚`%O�����_��j�`y*{vϪHѢ��	K �J�\��s5r|.�2X��c��3���E�$��h�١�Wea����~_�p����S��+��`-��T�����e�q��r���O��x�	�B�S��3N�kڝ9�֧g,�h/Ǿ�N����Yx8��u�A��$�#�9��启,12��LD
C�v�D� ���"�U�2�e��s5������_]�2�S�.��ww��b�E�3Tv%������~#�*��]
/_狜`�G�i�I$a"onf�9f�Q��`H��dY��������$Ah�c�\�͸M����=�s���5�@��E52�����V`gͦF�9�i]:����N���ٚ�#��1��1��c]��d�k�呗�RD��_i�-6*16
׶�q�| �5�-�W������ 	��0˾��-�P|ᶠ)i����V�	gS�����=LiK�Μ�n~���2���������� �i��k��b�D4K�7��wćB�2*S�h 7��t�=r��$�\}ɡC/�P�@��[^H,]�h�$��F�ϼ�9>9QD9��/��]�za#;��[^�=�3\�j�^�2��F@od�VQ��Ǯ*+�H���y��o���b2	��n+CgDTً�+$7fQ�X�*�#O��%��n����#���������v��g�ɘ�m�}�����ȼ�~|��沓���+��+$��&bd5�o�dJ�T~���҂�U���lgb�HPA۝}�q)]�p)i�5�^��8�s�6	�
�s]e����>�= ���iR�4����'���K�̌��y�0{��rb�O�'�c�i���aY�2����r��q�� ��	�S-�t@�����q��Pg�"~��*�]5�.l��T�!DzU��[}D-)��s`�^���_̠����뗖oN���Tg_�/����p��^��rz����wX�$���:�;^�L��c���o�w&��uJ�[w�{5����;�#�@�iOug��Yi�^���6�ڻ�����zG���=s��������ʘ�ԶD4�*y��Lci�С}�5��7��6
;r'���kgg�`�����D�A�0�@�0t�g���Z"]5�����$oҘ��[��ɗS��p�g��
�U�1�:@����;��\�#lL%<zSwe�\��ؒ��*C��a�/��
#����N>t��G�\���8�%��_3�%8)�}oQ�.
�֩�m�z�(�e���R���5 33���{=|
��c���!�IҒmP�����F�s�=O��8�m�nH����Dr��e�m��!]�D���#�����rO ���,��Y�_EQ�A�lS�$�o�i�A���G?B0������&�w=Ze.CB;8}, �J�i6�k60��N��(��l"��(�qG�������HܧT��:��`I�A�86��2��|��J���k�p�=�%T9^����Y8N���Tc�_E��	�?ߢ�'KV @�6�`@���Ó�5˻5�<;~���{Tyrg�łE�������©�pP��Tbq5��eu�Mp�N�=*>��s�ᢗ�w�{(�^Pn�/i���������`E���s>�p�s�_x�8e���f �]a+�.8˜�C-��O����J�%�_%��4֠�%C�Y���`�_������+io2�k�� � `&n�[V���]6��`Gd�����{�TP�>(��,���B�8�����)UAB�#�y���H ,��E��d+{	�J��H� �,��>�h�&�q�5g�d�[������d�s{\���*ĴH���-i��� )��(UhIP�[_L5AEEKR�9��Y���<lߟ���nҢ���`cϨp��de�u>Ai&���(wQc���M��,Ա6�����[ҙ�ƣd��`fkg�c%�������$�Kqy,P~]�ICy턕�����W�]^K�^YBs�Q��j� 9nZ)G�eL�3ף$��b����r�aT�-"0;V��4�	!���i�β�/�m��&S���Ea�����W��lǯ���QywZ��X� W�u;����\������L(��,�����d�Y-��}	�n[겨��ܥ�a6uR�b�=�`�0��@�.��-X�Hy?�@�5��ʼ��:(La����.|��$�Ю��L�����d�
���a�^�_�D\���,����C�F8ͽ��j���{�����@�*'��\2[�Բ8����e��?���?����}�~��SNg\�[�E�|�u�E���.�!�AW����������5\����˃r�,����Ղ�r�pM ��N���En�5U�<4`щ���Gϋ��o6D���Y��c�"���n�&��5��I>�7Q�I��TK�#q�_��m�5�!�`��b�Z����S�t��t*	�&d��%�������[f�2�v�����M�o��j���h5�6ec���{?�x�y<^�m�,N��֕)�����h�RVP'��;�nf���$W������W�[��wpI|������n ��^z�<P_�p�ױ�Z�Qۤ��ы�745�a{�1l��O�W��C�\�:0��
3fGb�"��!�I��gE���0O<+7��3�mT5��VW������	�ퟰ|?G����ĽQ*��c�ܞ�����q���.}p��
�Zȧ 5�jb��\�hT+,���u�a�适���|�?+X���h�2&��u�;�᠛�����
��� �59d��sw0��7þ�y*��oý�T�<��<`�5{�x�E:�;�
�8Ee򲀤I��ۦ�a��r��+5���9Z�.X�Y��][�m�a�y
)�x�w�=�pm�\1�X�f��=�v�}Ĕ�b&����&��,v��������#�w������H�[a(/!d?1�#qگ�紡�f����J������RIZC=�Ä�;��=�c& *.+`ӅGaNYb���ȶ�R���:X|ڠ;��L����5:	��@���(�O+� 'J�J.��7$����LQ3N��L�T�bϢv�wvIU�G�bjۇ�Thd��&`n�c�4���G5J�����Q�)D��8UlvOum&����eN���V"�H����K��ʡ$��7�/(X�a��m��������<��P$s6c��R��O��1������څ�����{��8�Q~����6lc\x��i�*v��4¾��x]0NC�ۤ��y�q��Wᝯ���OMЗ6�ߤ��=q�]z0~iJPE��y�O7��vA�6f׹�*�(��8A������*bF���=]�{���o��Ǖ8W|;SZ��!���<�sf��[�����<�a
ֆjpU�*Pf_F�լ�EZY+�[En����%�T�4����~v��ce[��&Jy��	4-�Bz������;�B�5���4ˁ���=�iKߝ��w!���|�P��?[�6��o3��4O���5!��08�/{�[����?��	���!���o��4��}�,�m�};�&�R�&!I��f�s}�I�e���� A>���*��nr�;�tiU��C��w71�A{��ԟ�	�t9T��]ǌ��{�(!z.+9���A���n�琮�w���u;E�oE�5����̿e�Q&¹��$�0�S~���毫pt�ȯ���/z�������ʀxg4�U���(���'�hK���ǳ��*@�F[+�(O�E�]��N¸rU�¬����0�0����C�XoY"T2]�w��<��LS�=v�k)/|��~�3��`V�@��.f����l;����=�0�?�tsn�L�E�U��(]�b�Y�gm���B�Nd���:��LK ���,yn9��L�q�2���k`9X���KQ�S�Niט����R�j