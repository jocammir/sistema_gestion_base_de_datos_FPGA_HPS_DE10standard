��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0������x`Y�sc���k���`ޅ��''��J3.k3���đ����}�O6"%C��f�ق�v9���"(�d��i�c�<�]:Et-��=h��Yp�)��1���03e�uJ��ka�%�-K��U�^o-ޓ���[[>�ÖaG6��,'��W_D'r���'w���G�LRD�?�:�N̮�*�/ߟ]پ�q����n-��!�<�UhQ�b�#�ŶgI��i�ps-�Η3��TЧ(4�������r׋�F��w�;�ɠ���9bP�{��׊�ÛӇ̂�r���q�@�k�S�H���-{�Aj��sW�v+1T|Y�ԸK��`2>��8bub��<�7�P{J�b���|}��b3����_( �][���{�Ȗ*���^)  p��k����b[�ax`:،W|q��̶�F~����e�]k�o��?����YU���
���>��S��������P����؍@�%�
��(ot�1�LeO.�ICg�Oۗ�G8�bSJ9�AÝ�L I|?��d�b����`�2����A��LnŒZ1pR˟�C@Q(�~�Z:�iC6��he4�N4��n�!�G���M��jmF �c���X��	Jmſ����V�襰�Ɣ@���`QHE��H���ʦ��yvvǚ�!�B2��=�=�ӧ�i���7�`�q�r�А��2���c-��.�"���_5�7�z�l�WGa|r�fͭ4�9vb��t��p���X��f�ZBȊkI:��!e�n�|A~@�c��w�ч+��\?
`r�}�tW�B���
\��gj��Y^��7�+��$�{(��	��;�gc����n���+�	Q H����Ý�w�VxpX�v��@��do���4L@��E���퐦�st���b����6.#���a�
���"���
,��
�k&���A����
�Z�_2~ؖ.g\�3+�4KD�y��wj�����,Oݒ������["���K�Ol�և�a����g�1�2⍭9�Tj��Z6���M��I�����N�|M��oO�ʆ\��J�k	�3�QnU�ޤ�/�&�,CfBx�|�xI'$��^������F��H��ᶧ�hW��X���g������'g�͆@�̂�w��lT�cA��dXz�*2»Ҵ�wl@�`j�=�Ƴ�g�G�G��x+���!� ��וU���wؑ<6x��LW�m�R<���&�����y�ٖ�\|���cG��G��ǶP�b�zE�evR�Q?!5{	#�m�=�6��$YQ͂5{C1�n�7~IZ����=�N���#<�ű���d�����׼#m������R�����>坿ʒa�v�� ڨ���l��:,~TF��� ���z,����\^�AfC]Ҋ�{�Ӣ��)��WNbX*�A��w�Rl��[��y�B���/K�H��On���}0�R�*�a���v��reM&�l%޲�-�C$NK�1�d�S@��wfS����D���X3���f�DO����c5[�$���X8��&8�r		XcJϪ�z?�����[4d�85�Ɵ�#g�7X[3�U���D��
�Z�C>G�D黣m�r�4��4}�u�������`� �������H�ݲ��GC�.���!O�wn��iw�� �9�v�'����{�d�s7Ȱ��{e��s˷�����T�������.���I�K�hcݠ���pԉ鄍r'y��y�tl7�P8X�N4��|��2~��e*�`��t3,+|��e0�pS��c���lk�ϧ�JJ���I������HBNB��P���+�()�R��gʼ����ް�]� \��)�<G�σT��/�m��L��'�E�����<v�"��5�.��*[d-�ⅼCn1���8��,e���"Ž�����_��W��q(�צ��G�=
�mgR�kT�˷������c��t�(Ё����������H.�]f���Q���~y��.HF��Z*?/YjbՔ����"?@Q�S8'��B��x��3NK��-�L�5�b���Č���l��֘�1g�QLS�?r+�f���pDŹ1���e���.�F�EB��:ׅ�-���������5�\j��\��T�l"���1{��Z�jԯ�+i�t�s�}ڧ���\�5��l��Q���
�.�YQY�.�T�V�\o�%�9�%�t�w�����C�Y�Li7�#�0V�&��~BMw5z[�ǭd�}��F��҈ P�%?��k���B���*�%��@��L`�6�������`�寭./n�ܲ��(_�1���%��.~o"���&G��	[e�%������RR\�G?f���f��"�C����}T��q>���k÷6��=�Y�����1N%[�\�W�ƹ'Č�t��WZZ���Z��m�/U�=��Qs�����ZS/�b���L%2J#;l�����v�_�ա^4��ϊ�/N���A�s����z6�����˻x�	��"���8�Q�I}(�R����������ĩ�6��w��f9���鶊����y��p��s� A8���;`�h���Z��F��e��� �y+	���oN+���&y�3s��wM�#���~�0kb�ks��HƧ�f֑W��Ce��Ї"�i
����ڴ�)E��*뚋c��U_46��^ũ`��.����	$L���E3KDSG	�Űa>����Em����$�ӌ����}���}.�~gB H_t��p�ƻ��I$W ��%�4A��HI��dN*E��+�k�p�Qm��|�_�h� ϩ~�A.������N{�����l����ld;z�M�P �Η+Xt���v^�B_
���ǣ��^��{��J(�^�D�0��o��ؼe���5�@�2���� %>f���:vH������A��P&vF�5���/���%Wa�j'_��}g�w��x�L�DWM�h�,k��� ؏��%�*{`/G(ǟ�|����o�2�25,m���#j7�&c�9K� X!�W<"�,�� H��oQ�����F�.�u���
��&}N�h9�®)�s��j�K�4�~�T%wY#�������c�0��"�5r��^;�"U���^���B�hs��jA��S>��ص�X��T�r��+�*C�������H��'մaݺ�5�r'>3�Ts�ƞ6-mT�W�����Zq�Ey@��@�^if����|� �<cl�W����`���,�7nQN�E3Z��V*%B/�A6#Y(/����Ү3+Ne�((9 �g$Ln=�OR>y(X�ãf������v��S����9���9�o9����O��X����O��Tq�k����Á�=�F����E��cLL�d�apg�|��r<}1��}>J�n�4tF���Y�٩#��(U`��"cY���>��0v�?�N�.�o	����[�pt���t:��)<v<�M>�t��g坺̀.GZodb�+c|�i�tJ�U��},2�KwF�����������9'�´`���'Q����Je�G��|> )�
#����(娢T���험z�&O�X�Ic_*4��ʂ�3�w�W�4V��ݤ�*4K)@M�U�(��j	�D$�+`��#�Y�B��t![�:Vm8���v�mK����+����T��{�oZ�v�����>�����A��|�b2���J>�3Yт�V�/���̣�n781yޡH�Hˡ
�Щ�����[\7��&ͱ{�]3�ۯ�"�z؆�p[���}�vϡ
��]��D6���>@���6щ��^U��s����=m`ß��	?d�&��b~��M�&<z��/�$yo�
�3��(YC�U��
B4�,H��ǼwE#�ǈfB����P�n�_��P���,]��Dג}�b�pB|ܰH��?M	�h�o��8T6V~��m���7����T~B4�3�?tY 8}�[,��,4�b£B�K�C��/��-sՓ-HFӻ���#��A����#U�xVZ��*L:�벿��v�� �{y?jU�2Ї��WwB���De9�[(X��Fk��ӴR���aӠ0sX �V�4a���]f��L�Nqw��0���X:����f�m�WBsB
��z��qF]��o<Q���_�&9�{d*�:�����ׂל�7U�&�h��FDͽ��!��5�7-�a��O9	��=�k��	o�T1��2;��̴0u�qI�UX �n@�\����p��gl�}��p�~jkW!�-����&���P��Mo��m�lR�mG6d�
z�fI<h1K��*NS�-�r2�4�b$�c����^ɘZ��h�s�RB�0c��nݣxy�ӆך�'�ޔZtK!��F�V��Y���a��Z�D
���4�{�?[6[��J�c*.a�� %}o�#��/=6x���x`�l4�c�ꘌ�Kο��7U�9ǳ3��.��o��, �j���_��Lk�/�Y�oBy۰�Q��G�D�_��xth�eG�"T�;�P��_�b`��*�o�=Z.�����f���?ON�ߠ�H0�
ˌ���T@�
r�I��~	�{ն��/+[$�OD�B���~#�]����Ѷy���e�'~Z=��w�
�X4L���~3�@T�~�$���d�r�.�LX�2�Mx�r��=	\�v�����Q���?o�IÆ�KMi���I&��3���e���i[*Dic��b�v�f�^�.��'P��0&�#�6�X��F�0⿢9�M���b�o�NM3�[?�^!�L��nK$�*�ݭ�3a��I�!��<7�c��F����e�5_<_ G¶,*���!��vՎjL�D������8��"=w\��3FGj7�JG�
�Z��7#˷���gQ����W�s���h�,X� �[Xi���:�%zU�M���i�d�-1�жz���:�q���h�ԷO����0nB��G�2��U������O��oB���:�7�m�zwZ��SP�J�6܈�c�0�tF52��%��Ah8' Mx�=���{����/@��0IƇwݻ<<Φ�R���aY��]���%�3LG��]�02E�Ƚ���Ydd(n��͘="gfWqwa���ܑ�� �'�'�S&w��r|x�eI�G0_�d7z@)��n4cC#&6K|��ȹc�M�.{U2ɫS�uJ5�����D#ճzI��
��Ӿ��q���Xѵ����������mbO��5 �L0ʊi�������s��F�ŘHS��o��"���CT+f>s\����I�!1fŇ�Jq�s�\]V�Q�<2��=����}6��O��R��s��v�B?���R|�gJt�m�n委R�?*������[�O<�T0`�]�s�0�Bixr���p��e܍vI��(�
Ի)9跴s���l��bj	�+�YIH�b�Ox�}g�D��S�rQ����)vg9N?z�'��re_(�?�ͭ���z�������ꩨ�iu�}�G
ټ�w5��4|w��mk�EJ8l����������13<�rSh�w�v�j�$iG��*uV�ܮ)E@�E���l�o�ơ�Bj̀�wY�ċ@�����i*Q"f�>��ÜƵ��H�A�B��f�^�?P�x�,_u�LEt��������j����h����0�@�Q��>dr~��q.���63��oW�~�<4vM�)��0��E�ڋ��8�Z��S��� �ĭu����T�'�9F\�:���f�(�<�:���,��8쟚��o�� �,T��r�Р[;MZ�� ���D�B�XF�٨[C���J�B~��i?�8�"I�t"�7�qIX���c�����8�N�Yw�s��6άX��h��'���YL�����<�&i%Q�x�v��s���a�d�s�W!��E�P�����sc�tв��}kU�;]���Q&�꼚*ՌP�+�d��Ink۶9�Cm:Η�͖���_�c�������)�nx�l�iB��G6��U�jF=
U�v�L�[��>�SO�?�{���+K!�w=�%@[A�4� ѱ6�����k�#
���b��ܝCg�Ҩ�K�Q������M����"Uׇ��yr�"S��3up#�\d���&�I(�/��)����>%Q`���[�����{��'nQs�'<�)�����ϓWD�~�6eǅ���V�;��1���k�6K� �ң⡈��AG	��N�}5 ���Y�E{�03�=�Yh��L�w��C=
l+�e���bi3�8���ŏ꣖A��'��r�XWo���������W�2ZD�5��f8�M�.#�ߨ��o'��4v`��SgFG$���|`�N����l���N3���Ȏ+�rQ��@h�t�J���*��|���
����q+.�"��������ߤ��s{��z��	R;�|��D{/^˷�ZQE�:x<���z��86'c-\��dm��XE뷔8�l	%��]��NX�u4���˩�oйN1Pb��� vU�H>$z2G����O��l�!Vr��ׄ��1��b�I�����)��1ǎ���"�>��auo���H��j����턫�J��+M�gP�%Pr��E�|\��B?]��!�@�B����ާ�f&`s2w�d>����n||��/�L��n��O����G@o0������sr|Hk�|��@��Šz�_׊X�){��G�.w�<�ۊ1C��+� r�]���١��򤎬�B����e�0PV���9gZYjgݩ��6����EOD�A�n��-�>�6GM#�#N\�(����UT6�����@;�`*��"���Ja�K�l�hCb����W`�l.ۈ��wA�L(�������8ͲD�s�-b3$ވ<`��#֐��@��
~ g�=�f��Ȉ�9�Q�Q6�?(��G6%*�;��<���Y"$������@��"6������Omu�/��a_t ��L�~�~|4�Inia�U��l��G���3�;M�?93�k��~ށI��ΊÆҺ��]��U��c+�[�XYLnD�w��H�(?Bcz���Y�X
�|���/������XI�1�H�ΐ�O�2�{U�C����7�8`�6ހ�h�3���YE��xjZ�+�xx4�Y�����-�&'ⲕE�C(X�>�����4�z��Yi8�K-<G��0)^x6;~�R�0��&<��n�E26���s+����w������6�e�d�eH��$<w�3r-���|̢���� �G�~ڨ��*�qie����s&�ǜ��pz�V��2�����9.���<��5�b�,��R�0̒�wΧW,�N������\�E�P��8sd��6�����^+�⾯N�l��©�[al�0��Z�El>�g`�ZbK�P.��+`'ݖ�T#��
_��}6�5
�AkR�5-A�gy�X�F��#�F1�j��`�����*o���� �O�r�$��LO�@��t|[hk����K+:5�D��UϘ<ҵK;L�-E�t2���`�x��ϽՁ(2�������4I7�#[�ַb�}1R�wm��ϫ�ᬰ��a�T,i�0'���fZ�wn�V�;�th��P9��[�� �$��^����?>�Ь i��_�1m˭Ʌw��"�+�@ABϦd�
O��*�
D�rF(��*sT�U���4n̹3��n%�6/�&�;^����N/�Ѻ]��_�FR�#42�?����ZSBO� �*�;p��l��r�ػxu��F������7i\PK+����+^רa��:�Nݗ���C����䞅�Cॼ����?�]��Yo~��E�]�ȸ�N���;{�Q�Yz�5�//4�*)�.�]���h�4����-�w�/�gr��Ϛ�by���S�Ζ�I�r�S�wE���a��#�o	nED��O�`���{~M��G��Lx��z*�ͣ�v��V�;ש��.W���1��Z��#�e����Bm�g
�k�S��,���/��ޕԎ���a���N�ˍr=�9p��ķ� ��h���Gj2�M��r�)�cR����&��n iR�1uCeOe�q���_nԷ�dl7�o�`IX�#�s��Y<������%�3�~�z��-��̑S>*�ϡ�EV�f��}6`u~̙
�� >{Iw���T��^���u��tC���˖Y�w�ߔQ�c�L,+��<Qs�du��r��O���m�WbsdYۯ8�&��uѢf�h�X�?�-��7��5�r�+����˗�qu-OQ�2��bTP�2E�n���l?Anȋd�N�>Ā�+�[?!@M�-��e�k��a�=J����G�P���F�� �ZV���Wp����ݘ_�P�GpWZKc��"��cI�:�6Y'S+�P�D���B�,1��A���KPu�j���z�Y���_o?�����N�nF��+Y�B�"��#p�`�{��F7Nfړ -���zN�bdN��V�/�Q(��~"�޹��:�U�M+ %R�6ǹ�C�MsˋxdV���|��l�>���M�o��*D��"<
�?��E�?�\�56����P�I��,�s�����#����0W}��VP��)		��%!� R��i^W^���ړP�`@،�s�rc���ft�x��v�!�q6�y�em����6�n��E�&8I�a�<c�zA;�E��PPٌ�B�;6�������.�?G�&�@V��Z�z�Y��C�y�.����}�P���`� 0���<�-*�����OH��0uv�F�2�9�m���+E���ܼ����#2�A���@��;��X!ԜJ�V(k���ؕ>
�}N���9!R;ʶ��U�6.�����Y(�ǻFg{:^bk��"��zVK��ޣ|���G�
��P�+��Y��F1���y.R������%�ن���*�Y6鮥tGB��
�u��x��7F�;�*��c�5�J3A*J7KU�F+\�S.������,2��3�BTX��-���QZ���1�mk"��	Ѳ+�#2�TT�0s+�B�Ԗ���(G��˓ �~ך�H0+����RD@C�4b�@���؁�TVh��Z�F\ߜ�Z�z��K��Uv�#��zIt��لO�M���<Q�Ӛk��j�-���-)W7�)K��`�,��c�h��5�R���݈M�t�;���KxTA�1&�ݽ��J������CƔњ��y�����3�p�}���\�X�����B0�Y����V��1g@g(U�d\���_U�B�7�a�
m'����VR�x���?G*f7�����@D���(b��]BF �}Y�إ1�T���4�7��"}�N���z�Vw Kꨲ53�Mڻ���䱙�z��|!V�({8-mU������AcJ�H�s���q�x?$����91�/����fe��,�2��"�b�ƱQʣG�a�S��I��y��l8�nf�kx�[\���|L�i�6b��)8���(�ɧ�H+p�*T5������k9\�`�i6K���']P{��n��{7��`͖�Y������gv��L!*�䩜U����F&�v���gl�����<��1��y&ݬ_�z��eYid�g�4�|/�w�(`���6��sC��W�v�����S�5��c�mU�a=��j6I��Y�6���ֶ��i���b���(���Dn'�ܘ]g�6�޲S���{;Y�*�\�
8.Ɯ%G�L)�e�S��G	N�Iۛ�Ϲ���r�Ŏ$�������&�!�bP��n���^�D�|�8��3r�����XL�� �� �{���ƽ���g�ױ2qeD�Ki���pa��j����J�(�O����n[�o�]�T�yW�9&\������(Is|5+��(^�q/��-!Eߊ�	���%4��CF�.o^�C�hʆ�?+`��͉�F�Č�?
���x���rw�$��>��3�S�;��g�r;��W����f�u�����G7OÎ�� �P��<�}�+1�Ւ-Nֵ7���_�e�~3��6�FL'L�����`N8ѩ����7��xv{I�^"��M�h͗������ws�H����MV��+�(T"n�R��3�	�x�8�}�N)����
��͋��d�9����x�Gp3�ͽE������4b�٪�Q3WMN�vp�b: