��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%������Z��B��Z����eS��D���Kg��
A�N�(�a��Q�n��U��N!8ߎ`ۼ<-:[�t1 �m��PN��߭J�]�V3E@m���nf��,rﲴ��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0���7`��&��ӽ�r�Zŏ:�j�nu�	�SO�e@z�d���b�y� g��Ø
>���c��������dL(p���>��a�;ENm�ykߏkӣ|��[������O�`ΌgE�^HKmHI��@��}���c����5�o�5,���"�Y�{��K�4�H�M�t�S&�~�Z�s=U7�5B�u�[o�g@ٲo4N�k���]
H�s��,��S��꯲`7�A�$�#V�IM��p_���V�3��t�n�XlsUK�#U{�ѵȻŖ�=�@�}��1wZ��A�`#�s�e-��f��-�Ν}슇!vP�ZaГ_�~o����h� >L��tK!�s�g@u1!T®|�~	�L!y9��*/j�����]�C'I[<8j���|�_N�X?��6���#� z�n�g
pb�3}���j��8�9w�$��0"��DI��7�k��"�I��e$�O��_�B���A�4��1�݀�ؘ�}�).�ʧkg�Ӭ	KPh�L4���� �w���"���o�0\ߘ�([^2W?:���1�v��R�9V�����h�s�Q8�,���Ř�� t�|�����O$,E���J����e�5��F����{֒���H������z/�DĒ�<8{�`�,�(�X^X�?�[9[JV���ܓP�zS÷ �H{g��saPzA���)z7�O?�Y�>;�+�ow 	���ƭ"�,�j#sm��*�l�Y�{AAlji���U���5���$
]��v₿V�ϡ �C/k:P32d�H�K(n�=X�7t���9�;�5����.�vg���ǒSG��������=	T{º�l|7����<l�u$�9h�V��ܬB��p�)6�~Eo�H�U?�b� � \/�7��i�"� 쳭;zN�_#�_��V�p�D���)�3�l@j�-���l�.͚იQ|�P��o�Rx�_�iLA��BmΆ�ߓFp6����cً��t���:T@�o&���wK���9�VG1����b_��F�(�N���	��\f��k R\h�%wUc[炄=+gg���/��M��lڐ�!ગ��/%�`*`��X�Q&�U"s�q1a)�͆��îJQ��<+N�C>$��!�Nt�������	�d���A���	U�?���!�5<�'���Z��	� �5��;1����ųO-�w��+�e�/�9?��\�؊Uc�Hl'��_�A�*i�w�ax���s��D�Va���'�s2/_�}`5=���%�m�@���Y�s�$,o�y����k,�1f;�Q{�I%S�ݳ�A�@��.x�*�H:4�e�"���w9.��i��cG;�VE�_�����V�=��L��*<�k����f��X}s�0����l ���@��"-�*���3Ĩw3Fz}���.�Ɓ6L�9U%ۢ�x���^���L��KM��e� �>��ܩ�i<n��wC�p�c���O�D���ȭ�w>Ti�JY��bh6�J��N����[���J�Y���E�lv�s	�Y���D ���`�~Ai�u�&�h豜�;Z'���`P^׫�����~ǂ���r�9t��Z��l�~wP���+ ���ڟ����oKw��ݑ���"���/yn0Բ��V�d,�FX~��ں��L`��>�l�t�dŔ�6�ܫӏ��ʸF�~I~�5��oI^5i���Jx+�q�IOR�!�������,��en�:^m��?�`��R�	�H�c0�Uފ%#z	Ѩ��ͣ'���ud+����tڇc�ҝ6Q�Ԓ;�����O����iR���(H3I��yf9F�;�d$8��e�F	�j�u���P�3� ��?����^�^����A�f�OQ2h�X�3޹t`���?�Y1����o���<�����_����'rá0���ZK���>]�e���0�0h���>'��{�6��o�m��zs��)��a�3��b:��zߡ�����$�����Kc 9e#��P�,�j�`�z�q��R�Nϐrw;�;���k���RLq��a����J_iRE�j���g�U��rzcȒ�I�z����v��)�aq-��µ�����
⦕5'�D�T����M�p��릧5dF����H1� ��+�� B3~�#�	5í�&��L�aƟ���U�vɤ�Y㲐ư��=��T�%�ۀ[�A���yl��݂�ζ}*�kv�q]uݙ��[��(ʮ���"b%>:_stb�t�@��s�Gۘ�����`����
�gcP��,�wc_v�o��8}���9u[s�����x��攨&��B �d8D�鿛��'`��D?mVˇ�+���C�a�Ch�*�q!
�]q�0XT�Hk�E��4�	
�>�J!w6���H�ڻ6����_U�l���#:=v���D�3�07��Įd�;s�i.]Rf��4/�oS	̓Ð���*���/j"_��b��a�"�LwI�jXp�!C�<Ol�/��=����xY�%L|7N�4��غD��-�}�b+c�d�(��Z4�]���������}������nM�`%�]c� o�h�V��
"������H̡w����M��P��Nŋ|T��6Va�hRx�"Za\\}���b+�2juĪM[���B��IMx)� l�l���,�VS��~�v��w5����F�o�>� <��-��f1�]/�i�h�[������o���^?�vA���6�����t�ݧ�a���� rPU����Q����
 f�����ħ��$W��ށ*���{0$7C�R�q�X���D��5�Y���;�JQc	����̉������:6����,X���Kȗ��}ֹ����G)��[/b��P3��Eg'T��Sf�;y��ЌM�WH/��&1t�d�Z2׊X�d�:�.��d@�yҴG"�N	2KJ0��!��\�2�Y�ӌ:$߈������0��c�u݄��Lɬ�YYo�g0�b������XC`�f�}��.*$�ƺ�ק��ZN{���:)]D�� ��S���`�ɛ���W�]����Tg�y�4���LvF�s��ض�)D�7�c(o���6Q6�upx��;�̔]��fqX�*�h�7�I���&�˙�o��Q����caΐ����4�"���	@O6�yΚ��lP1޸���q�>�l\?`�\�8�\~Y�-� E�VG�g֎:�pQ[�+�}!)� �	��ƙ�8�z���q`�iVz{�ײ�IaT�L�YO������� ]��퍰/���Z�]Op�tKK�gфu�Y	 �f�g�`*�}+8$2,J��(S�d��b�I����G������Ʀ��U�l�c���|�eFj[�1����ر�|���Y>�Pi�LUx�=r�WlbStx��,��w�T�����G5���O����~�s��i]\��Ѷ�S�aq��S� �v�`Z�R��O�\T���t�t�h%|U>ǒ7��-��@��-_�e:� ��[-Yā��f>�*������x�=�W���S��˝��Y��̢�1���ֺ�����]�|Fz���V�� `ǉ��4���$�S�p��Y�θ�~��W��]M�t����NM
���Y�.�G�ITQi�������Ck+���`j��!��i(�|�Nu��T]��/<u�y@�p�K3��oi��
�p�O��a��Ǧ���=��j���߂ކ:�_��Q���ο�P��>ٱ����`�\i� �2\Q섿���,�ן� �/����<���J��t{���*���j�Zq�l@����Q�_՚j�1��x���*�v�+�/�7�ڌw�Mq�j�����Yvz3����ީ��12��!�JM��ҥCg񏀪v� ��ϳ|W�̃����V���ʆq����4>w�=1j�+��B4{�У>8�C��Ohm��RTBY�
��h��:��&�Om�!��kn�W�=�0?��`�͛9��s�5	З����
B5��=X���`7i�Z��˵��q��9�����\��d�~6���)��d�`SK=�>�y��+���U�����������`�`��Ԗ���>��'Xk����dw�q�f��0Uf��i����$P)3���=au/��0bM��V�>��Kј�a9����/7�⏤B�%O�˶��K?%�:w�����lP�(���z���Ŀ�<���k��o�B�b���-�����P�1��)t�.;&d)�,�anqeV$�A��O�Z��@�V?�7���,�nW�����K�q�f�-Si,���z>���� A�7u��N���>v���u��9Y�;AK�Q�
�֩�-�f�����x��PJ�-��!���&@e�&����ޱ�́e�Y��Z4aH@&�'��9ܦ8~�������d�=\�e�q������-��ȶ�%<�7P�z��RG��Xl��C�-\BjVq���qb��Gб����%�S�-��W�bS�����&�͟/ڂ�>(2�b�j�2`����>�O�=*�hG�w��@�i�N6�:G���aH�c��>͜�6/_���&N"y�\8l�9#���?bf�^�h��ȓ�M�H�U�Щ�.I�t�z�?8mc=Hm/��A�{)K�.�?�A�L�:'K���!��R)W��rkF� *�d��Gn_/Ҭ�偻��!�I�2��>#m"p��0�\�Dޖ�{�4���� ��f�(��&'ǲ��+wB1cŵc�X��z��'�ۜ�w��{��a���@-�''r�࠲��O�b��h�'�/�G@nH�Epc0gf��'��(��pV#��y~P��ͤ�_7CUO����?É
�E`ם���0��Li�+'�F)vS�m�g텍*d��4�LQLA���w���۞_fK�t�b��)��qq�fo� ���nO�Z��Љ��q_ �FWa�����3� 62�s�ʩ�#�#'�sso���&,�3^�#����s��
l�<}�����-�� Z�~`D\��	��#Y)ʫ1Y��ۀQ�
��z������'�ue���dAsg*V����%q^��G�U����X~oŤ���)�M������S�̲���,����������z z$�����#��e�NDqkÁ�l&��#��E�,)�>I�H-�'�����+��aC���Y�;|����/����7����$6�E��<��ux�����k��㠪~z�ֆM��W(�h�ħ�e'GlTb���w������!��J'��#���x�a*�<iN��D	�}���0�n���I�Y�ЏC��@���K6.��U/��-��� ���V�vIg��꩙}M��h(h����T��I2����+N�
E[�|���kw�-2�⎏b���d��Z����LMz����
_���B�;���_q5�{��x�1ú��h'��^�V�|�c����'����"ԑd@�Ov����=�6o-{T���C�K�yH07]�Rѥ�y�p��6/�Qx�{�#�n�r������3M��&ᐦ8�2C���z�R��ȐR6�-���#����,�ٽ�f`�,̪"�v�R{�Ⱥ�%'Dʆ����܂h��/Wen(���n�D9���=;�8A `A���M�CR�WF���s�}w-j(��P/b����n�z�}N-���J����L�D���X�^�<s�|Nb�OnD��mU����H�s�]6��V9G�w�p&�A'��zCʗ�9�tm�zBp�-y%�����L��b���V��$n}�'<U2�+�L� K�P��ғ������ �]���<��~%a����{� �՚W�0�8F�)uߕ�_��65v r�kH|�< � ���{OF������#��\�p�����B�<�G�=��T,�of 8�^ҝ}������Yo�m��ݥ�A�T�h(�s4��6�˷����"C�jK��j��W���?n@��TA&�!	1���t��4�ȹ�	\�0#�QT�.Nje}�o�������?�Sl���Y�w�'x����� 1-����a�1 ���3E'� 6��G��Za�b�t�q�r�:�L�����aL��i㱧�X�������><z�A@U#��i��N6�-��,~Q���~~8N�5��8�k�@�Cp��^P�̛~vh/����>�`~V��m��D�@p�klP��MY�������� �<áh�4�%�	���7T���3=ϡ����J;*f������;��  W�o�j�j7��'2<$�&}eNR�~����N���-�k;[�G�p#����,(��/ॵC�]O 2�rZ��O�p7��啑{����!'7>�m�НC�h�t�yC}����W�M��-�+R�{�-/�MX����I�uV`y.��ZS)2�J3�A	/��H�����ݚ�C)��X���Ӝ	����Uw4V�r�	S��ؒ��:<�;q폛��7K��@^����iL3�����{<1�LA�_�~�S�)������A(�=���Z`>���vl��c�|u'1b��Q�pKe�Ki7�7Wdu��n&=smY�Gצg�*z�gv�6&��ޞ�5���m97 ԕ8�R�s�r�|�=����*[��������g�םe�ŷ�Ff���
���M���)m�$8�\.<�Z�� ,%;}�����>>Q�U8���;{���Pjt%�l(�-9�;~Y_凥��k�J B�Pm��>��\��@�J�������A"��Գ��I��iy5�{9=��crz��ⱼ�����,:��g��|,��2�(ҕS��20�*���M��B��L�&�ǥF��bn�����4q5�vG�eȔh��>�a�|9�:�C�%l�ԬH?o<�${�l��<�F�V'l�����[_m��c*>�<,ўc?��`���S��
�&}a
��˺����6n@u��.�Qֻ6k��JH�.ޮ�مDJ�$����g��yP��߹�(�<�|���ܒ�wyF�b	O���jiA��$\��w�I�f���|)�r¨�'��h�=��>�yR�@�f$����Z��V�l�×l�&TTj*qR(�j�*�Xw��^_we�s���}8��h6,,�U=�U�)y�h�?�f��z �BGvTC&ӍÝ��9Ă�l���R��@wb��#"����l�(�e��QQž?]ޚ#')"-1%K8���LDۚ{��ذ|�R]*�����2�noy쓓E%eæ�������Z���B��z6���	��7�{x`�t�6�;Lui�,�P��8G�2��\ey4M�[Q��&��c�&�o��nd�'�e�N��[/��4�H���G����ܬ����B1�u��O2��H}�0	}k;ij�Σ�g}@����%�b�B����)3Q�%���-lY(�F��+�PS�ɪ%O�>&��ѱx��רg���p�en��iX�.�T"T�vأcQ�#!Z�,0lm%Q�d��v���¡ƉmP�1X�1�1x���%,O=7wg�\^��;����K�~��k�<B��dE�k0ɮ�0y��aw���L4�Y�\v�F�k���9h��Ǐ���iA�U:�́j��I�#Lc�%��SB�(���%G�+n]z1��G���R=�X��������3���*-�qY=J�g��{�3�<?��eԁfh��Z�� �������2������rMҟ��s���?)�����Nc�E=�Y�a��1ߞ�n��������]�s�77{�!o�:�&O�4էX�Ȯ]F^)ަl�I�"���m>0l�d_a(19y��k��Q��9��юٛ�Y��x4���¼���耚�[��r��QzM�%[�f+BwE�X�� � U��ۨC)J�l��{�(xӞ<�jN8Pߎ��w�2�䝄��fs��\�L���Ja�Xd����飼��D	�Y����b��[�U����@[��$��_��V�q4���O��a�y��)�Rdkq�/J\IN����o��\~���nsD��P�V���)tB(����ڔ��jc����<$XB�7'�j�p$�R�;qB���8�<�,��s�v�����n1iߍ{-��'A �}��1f����_I7�	r�lj3WpM*�4�rya���m���݀�ׄf��f������dGS�tx"B������F���W-�������m[�1Fg=N��R���/���<b0�@��2Y�g����hɝ� Ζ:�}ixh���c�!/�^�qZ�!@�8n\Y:�V��9@��:��gS��[R:�,������ʬ�/rKWa���o��bu!8�egM��X��i���g��DOԣ���2N�����V�W�~2�R%�g�Wu
���`=�__X¼ ���Io-Y�{ 70��v�����晳̄��J{�<8�(zȱq�����&�Hy��i|����Ii!��lH�s��{#��ێo�������D����{Ӑ�����У�F,������&n�y�����^68��m!�'/��*+l�C��f3�q��P9%@���E��"~v��|��n����ʹ!�nn4]�Y���آdVm0y�����eEgr����ћ�%��D�N�Ǽ�JL<�	�����՟�K�V׆���xX� /��� P�R�	�\"��c:-����j�1���� ��g���7��N�]kӪ|rDg��ycP��#5�Ơ��j�?�<�&~4B=;��xtWe��wc�͒^n�����g��aR_]ᵋ)_��rw���4)n5�Ko4���!�&����� Qz`��g�}k��NjWu˻=>R_Wb�x.#0��X��\v�%�:v����(��	��m���!�/���l�!�:�㟲l�C��b��g>�a�Q��!
��/:�
S�]z)�0�R�t��¤�9�sT7⊠���zk1�N-)^��~����\���^��Q�I!p޶
=1 �'8 �c��7/e?RۣDr��،w��҆i�S�$�g���z4	����!xܾ�~��t�~j���+{X����Ј	��,�̬قh&c�kѾwa����|�aw����F'����P�FB^��
�"�L�H��!1����V����
O�D2�v�Z�n�e�>Y)�pO��r<_|�kw�����!v�]�r�I���ZRm�>ƈ#�{���>�^�*jHT_��ʌ�;���"ko��0��q�*0|��w��aT�u�If�/y�шM��T��U�T�0hz��nR:l41d�B
��H�l�b��4}���f�tS=)i�t�y/�|G񁋅D#�o���l�i�z>�#|7���[��Ea� LP2%c.�)�����v�����l ��? �X���ޖ�B'խ?���`�h]�a�i�k����W-�4PI��z&����,�9��0�N��Ө�4��J�WRQ�!5�A��!�C�/��t
�#��E@���=�ϵ���ny*�x�۷�]�QC�����%��F�$/��
�虣,(����Ȳ�|��Z@
�K8�s@X��bJso]��_3�i��ڛR�iǆd-�ār�~å�3�W��R�xF?�����:4Syh7ԡh������徧��A�P��S_�]�DT'`U�\;T��.؇)u����>��Jbę,�/�w���u}̃��ܨP<h���G|"I~�M��������*�"��>�wJ?�+��#�r6&��*f���uQ
R9�s	λ�rׇ~��L�i�K1K�~Q�Do(���z��Y��E$]+a-�vx��>��W��㲍�6�z������:h��Ui?|S��آ�;�9� ���*(�h2}\Svk�=5�I��>|�~�p	id.����p��ޤ�Eƫ��Vk�Q����ܶ��\���G�GȾ��.��-�YW�0l��u��-���7�_o�(a��d0�/����ח����-�H��V��/`���`<���8=��q	@�"���4�Ŵ�L2�i&@�(� F���c��PD�� ����~ޱ9��dM����!̼�s�f!�`�P�r���M��{#�]L�Ec=�/6%P�Ⱥ"���B�H��t�����mؼ#L�6���C�~d���0��i�������$_�,a��b��t�6W��қ�SБ37�6QL���,�T�ݘP�������?{bE��ա�2����@ U�7����&@�;_��_1(�
;���Q3I�I�5�Uj�6��]nz@�V�I���R[�)�^�ͽD�cL�@������3�{R���qR�%�l>U'(M��#�X������(M�[�6�ɸ�
�*�q���ף*�˼㡛��]�p{~*g��G"�}apF1Ih
fZ<�/��&tI���(>i�ϼ]xsA_|�'o��d=|��ħ���0AKE����cր���X�䅑d���}��N� p�[O	��N�%s8�^���B$Q��f�8R�S�^�T��c�����3c�S}�[��.1��F�v���/��I@����]�r";w�e�vpNEF��w���pʚ����/��3`�T`�tks/Z��<c�s�>~�}|�v�;�%'�����"�$j7����`�q_��\t�Ӟ��@��wKè�[�A���a���6:
l��,r;�Mo�I��fJ�E$lt�{Ey(D�����.�xDW��	~�EuYK� �Ly��3I��e��8"��*���@g_?	r�Η�V�'jΌ��b�H��2��ݍF�o�6�05U-�M���R��QvB�	9�������x�,�������D��b!� �;N�a�֯��	�!�4t[=R����ȕ�$Y��]s7I�7��W�qȅ���2m��fݒ;��4��
�t�S(8B;�=��5�
��?��D_h~3�(I��F��3e��C>�c��ӽW��/9G� �N,8u=�PՐ5U8CWI<����&�6�O ���K�S���@����N7��GtR��V[�u��|b]���.��k�\Nc*2=����{�t<|K�g����<����r��������yE�#�x'����z,9��#���v�Z"��7�A^a����a�ۏ�LV��~w��$'�v�L��4����u7z���뼸:��_܉����'t�Ƙ�%f����N�h��,��*���<	U��S ����<�6�`L%��
*%2������`$.�y���8;��5�Y����'���b���U&��Tj�Ae%���z��K̞*㤄Va�%����v�pVe@��B��2r ���٨<=w�N]��k%��a��G>	�������&B@Ա��*�<�ڮ���t��7����(�Vڸ����BUy���$�V�-�:����7E/ݠ�y%�������De)��O�\�6�����&\e�la����2E��� ub�|s�Y*g�����	�����YL���W�I#]��-%F W���0�p�5�_�.Q��:hȾ�uF6o-�>=�����E#{IM��zM�f)q��r���yq�u��[/>ɾY"'Y>���#�_�ۀ07���ݞ��ˈ\3)'n�`S��(_r���ǀ���� �+=#Vi�&rڋ'��jN�ĄW�!A{=J�v|^�N���(�5}	2F��YJ�o�A�F\���\ľ��E���P� S�N���������Z/9�ƖƷ�7�skU����|�=��|�/�����3f��R?搜	���XP�x�Wd��{j��V.�4L	)i�'b_�WT�#ε}�?�)M�̸�� ���ĤU!�����3���'zϡ���J�V3=�H�k��?��8F
@X�0�el��İ�$�$�i��_�����kwH׿W�7��s��4��L�B�m}W{�j���,{�& ��W�0y�������$x�N�	q�o���7�X�B6O�]L�ʶ�;
A�u�EO�u��~z�L�I����Y��ҵ�xH��v����jh�Y�9wM��s^W�huY)��_�g�ҏ��.�:�i��rA���FWjЌ�xG#�-�w��%�� 6HyC�~�9|��3Z�>�FnD�_ކ�ၩ�����Ah�Z�ԡ
��q-��Ƨ.>V����[����r�J���n����[ww�\���q�6�6��e� �2쉕��kw!��/�`!�&
�U���e�=FJ|:���j�u�ma	dx���)�s�&��_Ş7O*2��q����)h��O@�^�qo[ރ��cd���= �y�7p�T\�B��}?t[2=�S<`��"�K����G�Zs��眥�=z�[�aK,Iz��]ؾ���Z�Um]m��1��V+�{>��v=�,"x�A����������������S�J�1-3H�y��Z��I̬�DUf���}�3ۥ�N��= ]�C֘��
}���wm59p����'�R���sb�tX`b�$nT���qe�m��2SDu,Ы�����gչ��(2d���Nٷ9����?�඾m���K�;��qMދ:�D8A;�5~�����}����{>��r\@��tvh��� ��l\�Z_&PU=����+�:��4yd��`9�w_i3������{��0�|�Z`6��T��d���.�eG���)�P�qZ�{��#5�]ɅX��A������2�Y�F{ia��{
�1�n�Z{hTWt�OGs�w��Q������ $�O%�Զ�c�?��KI>s�BU�>,�N��&���_O��\�V�����C��i���Ee@�����h�5��Do%�H�)�3Q���"�x�[�c_t�|&$��r���g��.C�*����#T ��'�Lc��0ͷ�B��P����3�យu ㋈?�s>*{��\��c�z#�1�c��4�ԖY�"*'|����ɹĂ��<q����ˁ����E�W��6�� �U�/̹��I~����V�:�W�=s�� Ȗ�G�dN4����SY�+e�&-y.ܴ���,|{�ب�"U�WJ:�=nG���V��BN�!|�3�-�i~<o!1٭MYm��G�d���ȇ9D���o�o����z��	������cˁZ���jf���Z�D��ɺ�N})lq�c��~v$�	ħ�K�w� �K�^�or��`zY���&�s^1���8ؙ�T`����<*�iK�S�"�Ս��_��d/7 D�l;�v��rV�-�&��\��1,/˺	9��d}'Y�yyOe,֐#]�a��m����G+��x��E��ʎ�Z������Bʈ=�?C���n���m՝xo��%puy����P�K�<u�yt��g��	Ji�*�RI��o�+���9���GIZ��=�Ƨ���"��u�����g��ѽ�Z�"(0�6d��W2��&�������#��UG�aj�u�9*����>e�Cm���G�Z� �]�oC�i��%��zCX�e�ꈜf@�Ԁjg�w��?�7Ȼ�g$q�;BG(��b�d�����ٔ�u��5z��n"6d�Ï�[��A�^VI���}Y6_�:	ǃ^����h\�����"���0�S���n7��D�Q��eծ"��˚���-�0`�ΏNJJ�O�^��c�e�ť�Vδٿ����z-
�*��D����*@����=��~"�޸؇��琀���4	�!�$-x�\�\mֱ3���s?&�9�������B��"�"ʕv3�%����Y'�/H��ӝ���G�~v�EUq�z
(;t�aB�Vw.�t^+V���S١pC+�ɈL<�;�QI������~g �zj�jh/ܾ�GafH�D�M8���=��c������k�9;��"��� o���ޡ?��` �ũ�W��/�t2���!�ÆL���	� ��������Ry59pq��A����i��͓��Kv7����9ɖn���=�
=�8\���!�ĉ���NUH���l ��N?8`�X��_ɍ�kj�r�(}�托`�{�K>%Zz ���G��.ed��8�����G:�Ԇ���%�*FD!��_���2y�$�}��:��B�%I�:$0-�g�(MK�&N|#�x$KG�<�9ٌ�+,�Y���S�a�~��Kf�.Ҳ�bi{4���u�@�E�óF`�L#P0[6���t쌙F���}����+���uN<���ਠ-��M�:����S�_Q�$�=�7��~4p뚢_�[�=���qfQHi��p� �6���N�JJu�db���5�,|�g��Ș��!V�mYY
:�}]��VmڤV�V�U�?�uϥGJX���1�BP�� ��6h|��<�柤d��i54ҳn�i�r�T�x[O�8�o�߲�����I���(;����%T	���2z*	����S���=y?�丠I4�-~�1�2��ǰ���A���C�1AX��a�	�N�� �R���P,#W���
��l��<�%G�掣�r��V������1��V�Oo� z��p�c)\��=�u����i�t�&P��r�j�+/�A��������;�>�w�$\y��%k�׉	�䣞��q�����E^ZݳN����o�1m����c����H𹴓}هtB��}.����S_xz)5����Y�9Ș1j�r�g��x��i�\���$&�d�8#�얞+-HCqsB��vE�����s�QR��^bc7�CF��E��0�L&7y��	��U�3&�2J���:Y<V��xl,B,������M�Q+f���Ս�e l@iT�xq��l��"R�X��!���V��$=�ԫs}RBVB��, A}b�5�u�h�5�������ȼNU5�R��C��2vI�C�]ֈo�J7��{��iQ0�z-h:j���^�Q���:�4|�#-[\q�c��;�s�{�䬓(�ŷ���'���M���h#IW�y���"��D����M++�������Y]������΁A6��-��}�㎗�x ���A�祷� �X��Eߒ�5�@ۿ�n�+�<�?���r*��2+P!�y��TP#G��υ�¡��X�<�����C�/��ɉ�~ ,�.Ԑ^�s��ӥ^?*��f�S� jT�F�7Aj���#������w�a�"�cIk�9����beP"�����ey�4nC���mr�U,�8�X:���g�C
�RÃ�����V���r��r�|����4e]��}~Ǯ(����χ�	� 	2��B�J&���X�~�������'^AA�G���U'��4 )όq��}�h�(*3�fIf�si�x�E��N1����S�l��?�G*2*xi}.ԮU�Y&�~S�e��i&�+q�RO�f*ą9O�tż��b�W��ش΂#l��a��]��n��U���5R�{BJ'����*C�B�*a�)�z"VE
�i$>ঠڀ54��ѭfVS�b��G�w�G8)�QE�P�>o���(��]-n��8����&�	�|�:Mw�-�)m*H�u����#��'|���vh��*��d����Ӻ��ÅY�u��G�u�(lD�C���t*ġ��&!�v�>����]~9�t�dD6Y=��U����B�Y9-U��Q �مf�����g�Do�6�?J�ú���O
9żE��ѬT^Ğ��@�k����0��hX��;K4�/8l�zG��q�����j?�I���t��w?��i�+��i�9nhH�3Uix85z�U:����q����Ø���C���9P��-4�m�3�ߊ��vr>�@��p{_����L�X�̇����H�Н�R�"'d*����Ӑ�!��ۣ::�>U��4��ݞ��V?�̜��<D�
G@���/	��>`��`�h���N]B�f_9 ��\�Ĵ:�IsxCc8��B��cU���.1��>u����z�R8a����(,g����~�k,փY{g�e���λ����	�|ɒoj$˂�f�  =^&C�����wN*��v�ʣ�C>��>0�ɶ*9���o�:�n0:N,Ȃ�?����B=�>u;�Y������]� sQ�0.,F��n&�#obf-�=�S���K]#<]�V^��H}�����{�^���)���Ѭw�	$W��{�Y8<�m�N1>���T�%05��?�|�B�)6���MHb�N���+
_q�x?=������)�!�{5��/�&Ǣ��습���2�#�W�'9X�[0g�Q��2�b�U�މY�3�Q�:�}T�nҤv�`�(#��H���Q�O���J�V��p�E����N�õ�����9��<ܗ�0�Rl՛Yx�h���YEkE�m��TȞ�|�(���.Q�f�cj��ʧ��*���,�7?�	�PG�n"���Xe���*��Wi�_E�/�fѶZ�%2��~�oJȵ�7�o��P~��<�=ե͢$����R��B�F3c���Wm���#��\b��C�!�fC��ss�O`�2�d�:��#��f8R,'�o��J�/�wl�����PT����;YE��<m6��3k�Mʪ�X�jߋx�b����P�!����+;�;�.�u�gJ'"H���tI �lv��HO΍P���.���N-!�>�<P�C�/�c��ޥ�<��5���q"W^9�5���(�����6�a�9�wc����I�O�o	%]�Kl�h��d8{�Id�R~|,�D�6�׏���Xѕ|x%�X�;͡p��/5���|,/ݔ��Cv ��'�)?F��f�V��B�~8D��#�����;�u��C��"Lf��b�;��
�T 3���i�Q1!��]�i������@���f��7�}�+�%�VBV˼��@9	��.j=E�☎`	�e��&�؂�W�B������wKx�"�h�o��}C8�N�:AF��$��L��z"�U��#�L��X,iphJ�6�r�L�>c~�%Sr��+=���Gv�����|D�~������#�ܞ�0�W@"�B]j ��`	�o�G �l� HVOUSxZ?���D�RU��xw�s-�MUm�r��"���?��q�t��1�+u�%����Y���d�xfeEyem�ׅH�����\�P�� ��L�����>�l��#��h��LH��%\��Y�H��g����;��n�@����Cݞ`"�6��P���r��0��69�IlPAHE"U�L���C�n4����q���q��JSiǆ!BV���W��9��8%�9�.;`�Ɨ,�.��%M�� �pkj�H�,��Vq)�h`H��Ϲ��:����R�5�t����C�M��j��գ?��m�����(�b{Pm5�P	��H��h�Ǔ��e��_�<0��&�h��v�Y����y�'_��وBn-L�~��\Emʳ��"�a(F���A�[&�k����Q�Bw�>yK����"��U���&�e���Ɛ�Y�y�������r��e�Tj5��E�=�p��K|%kQN޿�x�V���Iw�
���}��i�6�~)���݋�W����8)�{x.�!A�g�2�ĭ)�ԏ�2���w����ԫ0�o�)�5x��RxL����<� T��]p�a��&p�9�:C�J���a���d�J�h�_@��+ss�e��qo�>�q��#h!z��-!���n��?}��j`������|�߸�����>�~��3s[ ���^��U�Gpn�^\�\�:v=�ŧ�y��NaT��)z�
N�wođ�j�b��ԣ��e�8s¢OR��S�O�lp����v@�(�v�b%i*���u�������4:�~��ps{^�.��a�zvN���.�þ�ǹI!�PƪV���_M*��AZ�'B�"2�L4���bn��#��o���Kܚ_�'� m�?�ɯ�Y'����F�Ԣ:�zf�M_�L�Yj�	i�bA�E�q���L��5������%����$cj�u�HI`���)uf��'������乁d�yԸzܵr�lōW#���/&�Ը��E�q!�R�BX�ܷǍ���M+�~���0���.�<��!;���勢5���ck=9���W:��t�H��¥Ȑ�2j)��
.,G��̸���:���#����{VEM_�b͜�hd�t�����������b���sKQW+���|J���&D��s%&J�-�vk>��))�cN�
��+q|y�[�{n/�V*���	s�H�q�X��r��؜�H��V*ͦ���6҉LRlRs�v�����[���WEz��t�M�S���� ��/_�[B[�`�U�jt�*�6uYwK�b�V��|�5��6��x���
�*�\�u,o�Ve/�q3�Ct޼�&k#�r�S��r���؀�j��ȯ`
1������������,בV <Bs^��c�'��q�k�rH,����Щ�8�y�����ڛ�;�`��"_����d�q<��pmfʇ9��=C�]�1��ҏ[�Ⱦ��!�jZj��>*��Ⱦ�������=�<�,�%l��lkߥ	gM�R�kO���s��4��R�9��`����[[�E���ѓ���]2�|�d�:�6G�u(@/'Y�{*9	[=\����[V8n�p��Z�{7��n�����Ჰ��Z�'M��Vu��^�	��K�S�J�E�"@/;q��5U�Sנ� ���Aے��Л?/;��w��+�g���(�s{�[mG�ھ�;�?����~,�g # �~��������0�>����[�aJ���aZ '�[�N*'�7Y��ag��7���� 0�4�K�"QtV~�����b�t���h]�W�פD�j���@I`a���:`�/(K���F�9.<������}H�zD���oj6Q6~����zX�����㫥�xX��m�YIx������!�X�+��9����B"���lޯ��B�A��8�ا/��� �5���;�S����N�L����O��`�㇇���� &�Ɯ�a�I�;���X}:w�c��� ��""s��)IƷ��Z��9�:l�Ink^@j��r��'��0{/��J%l�DZeΧ�т�X��[�_���>��C}0Ê�
I�X�TvsZH�b��R �y�n���vT�������z��;������̹�
e��pB��tʭ��52��:��^M�L�"LW�/��8^;��"uL�Ŕ�l#�Em�m3�f�s���3�/eK��3��Gv��v�|�T�r���EJ�!^!N�dL*u�@�
�&���d�s�c���(�+���3�+�rm�a�����g��Y��q���Y��cޚ�����V�f2�q,�e&�����Zm>��I�v��¢w����V�K�T"� ����؟��V(P+�����'��;����o���@l�QO�y4Ż\7zSj���j��Q�'�*2������/�{��Y����{s������;�C��8I�e`F&�~���5��о�	{�ڛQ���F"i=�sW���r�bbB2v�
����o��ׯ�"�R�Z��k�Z���փ�f�o�����0Nސ��5��PK4a���	jQ�;��3����Rq��ڈ��/��Op����0
z������m�Ϸ9��Y#U(v'����2 �m�2�������Nߟ'|���k�i��9W-�E+^NPm�
�!uQ�2�8��	�`i�$ ���܊|V�����b�
���|����2��._|&fG8�w�>(�۹7p`��"m�K%��Q0�&1�]��ƙ҉�;r��iCRpy58�r��A[�A-%�V/4]�a�ekQw04���-Jjr;���n*��a�<�V�Y�,F_Z6���Ѿ)��?�Wt���,�U���_ɵ6*��jX��s�>�ǎ�B� a�ͦ��$��7��!�O��TxcR��N��v��Z����d�C�3nF�Ӂ 2ӟ�7-Yo@	���1��A� gn2����-��6:B�����E����Q�{�{i*�v�k�Ӳ>��_ig�ͻ��kb��"9�����1J�����ݬ�P�����(��s6��g%�(H0����r����(�I��%=�⾏�%H�����:S���������}�'=v�8�)F�{�J����Q�3�T�ra�܏������o�7
S��Լa\�K��l�oռ��[�F�]c�)ȳ��G�h��������v��"yI�z/h,�,�i��RD�NcFj�6Ot�����wn�79�K�*��&�d����yzb�o0>(>�,�۱H:���m�����r���:⹝�iޔ�:)nH����Jj�Mύ����l��nb�����!{�s9�W�̂L�o �R;2��!Ǯ.	��|֔k�"�&`	_f����S��%�)�yĝ����Hͫ�@�|��Y��u��`vF�֫�W�
���F���!�L�.�5WT6��&p0_��:��+�R�+���ꑡζ�Mw��o����F&�7�6����b��w��3�0�(����[g�t�I��|1�]sR�;tN	O�(�l�CI��%�jt*��Ė�͏1�Wտ�x���K��r�ҳ�cC�O{�űϐ��@�^��FR����>9>�3���mhi;��/y�w{ͪ��wnz�>ø���\�"Z�u�efu�*�7�D��A�܆�]�aI4��N�[�����(m���4���N���B(&�GD�0���+$�?��F�\7�:Z��롊�>�=�Dz�3 eN�,�z^����MyR�1 ���|�5<�Y��X	�b2�ɤ�Ȗ��n�E	u�Kj3?�A�v��s���O��ݜ���D�Ks����4��%�gɱz�Xޗ&	�w���;����x�擇�8��^u�Y]�%�6ٽ��X��×����Wn� �,���= 6x���nP���c�%�j	��G�V�h>)qZ����R��K����#��2Z��lv�-���1���m�vXL�IS������zN!��DqA�ĲLIJE�uI3B�����wY�B�XL$2C�ƪ7�Xs��� �a��2c.y���Y������VZ%���Л�L���+lW `�x8A軻Dn�D-F���D��۠
EӢ��o�f�g@,�h�g�ϒ��p��v�[hp�,[e ��1�/�+�����B1SI>p�K����q�NOG=�2]DȦ��S�l	֪�e��f�N�J槻ׂx�N|�������0Ik�c&G���=V�����g��!÷��5�=�hF�����-��/)Z�XY蛀xi����J�m�ο���8G��4��F���S��$,�5���t��|�G)�|r��s��-o�7�җ���n���)�~������Fu1z$^3L��!�c3�&K=�h�7�d��9��\b��&�����)���{���w=�Ƹ��
�~�>D:�%{5�Ǌ *�n�9M��c��
Op����zf�O.�P�mM쿇�ۡ�L�hI�W�k��O�8rF�����*B[o���x��+�{�9p��_��\�V16�����p#Z��hY����?��G
 ���*�b�P���IY�ܾs�rm�B_�$T��^�I�Ib���>�a�~S5P����N���u ���\�W��'͡w�^U�?g�ғ�$o���	�EK����a��λ����u6�rm7ы���A��1��a@���i#�
l���~(��-��<-R��U�Ʌ`��I���1$�~�3d�qV��\ؿ ���f�~ ��e� ��A���KE9�}o�ޗ���&�Vtz�/ 8�or�W%�w�"b�[6��C�5���}��\�7��?��>-P���7�w|ɡ<�uH�M|囧^�x�p������ߛ��9|n��n�_�����v���#7t���|}�F"Cu��o�J�%�#&���|��v�b�e�ϗ����;������h��措 ϓ�G���KΠ�����l��1����;3��<����@�(3�36��g�X�+�8�^#k"�h�+�����굣d������f�hj�� �������9�N�����R�o����# ���M�318��y�8���H�p��G@�M�"K�<
���=qS7��9�%v7Tڍ�L�ac6'&��V	=���Ow2J!1��k?�k�fO2Jݴ4�EmCz�	JW�	@J�o7����%�͞j� ��	�;z�:U����ۓ�A��Q�ßԓ�3a_ı]t��'��r�bAT�m%�V@�|�ګ���&�4�r$�D�W1���[/���qv� o��.�����sΰ8���Z�G�G)F˹�(���4I�Mwx����*P׮d��HS�yU�-�5�	�d�Q�'N%�ͻ�@���i�Cχ�Ը��u	{��:�Ѭ���,��}Y/Z��,�}\�V�Tb��󶨍���g��S8מ��KP�Zm3J1�g�+r�D��H6�:��*=�TE
Y��_ֹ ���!���W��9��K>ߚ+�a�󉟋,�����8�w7�����@�#�R6�^��R:#�H�-�^��� G7��!�?�]�Q���G�����D?r�69\��p��a��d�˜��	��x*�U�+t��O3���y�na'�d�$LOnl�kƃ6"���� wi�c��������9Ov+�H&l=T�k��3<K�C�	���~��.�<�z��;�ɲ�q`�ܼy� �i�	�����
�H�4��`��~�\�A�-��a�[W��+�H	$�2T���]�J+Kk�˹�L�Ƚ����*�����F�Z�.�]���W5�M`��7#�y���(w���5?�s
чaf������b5�z"��L��1�BNVҗ�Q�+��q_�Ax��oq	^1��w�H��J�'/��j:�~>��Ϣ�K�r��g��>�e�C��
J�O�9�!ќ�0�{�sD0.�|�L��a�7R3 �+��Ҽ�m������n�
�z���U��$���G�̤�+K���̇('�>U�j�/�B�$�4\ت"�}j�qa�85g��\��8��ڰ�>���k$�#7mU���9�c
�W�)=⨌ ���Hf��I;�c>����'�O|����};��gMJ������*��q ��(9�P��Ww�p u���|z'/��?	I����<���Bd�AV�d�jQ�P�1\�a��&B�A�4�\�X�+x�$ȱhG���/k��dn��$�����F0���Yx���F���� �Do�p�������E��m��y��`pA��D�I�CB��S��
y�Rn���Oϸ�r�lߜ���R��ܒ��c��.t����&��3���i报X�<?�V��@V����JC�=�?\+p��Ĺ"��Ͽ5����<�tu�*�9z�� �}�|��w�֫�x^�t!1��$ł =�ht_�*-�["����� �8N�kNY��<�����o�U�a��H����y�\��{��8%(� �L�9"����W[�E�7L�|�_鸫�!O��u� )��|�䳇B�Ⰿbo\��_�3�� G���zD�	\�[/T����� <N��~ö�t��@y�_PԚ��sJ5�N�����G,=-�;��`,F��-���E�J��m�p\]�P��{���������t�P���w%�c��&��}� �g����A)�+���~��AI�f�j#���Y�`���~���,���]2-��䨭#�8B,�5C���Z��Zx��:�A�͢g��vz����'��Kd��;���݄�*�o�~��jm�+8e^5�w\�7��S˴	�շ���>�=���  �+����h"�XT�Z��@��?�`a���;b�e��@�q���)���Դ;�^�6n�)q�Z�u�MK?� �ߖ��/��#�1���t+ ����D��2�8����L^�(0���wS�'�;Jz?�nL6�����,��rG���I�ApW���'��E�䶠�y�t".��z�Yh�˃2=wEa�?�7���5�<RF����;,�{i��혳<��E]�00� g�.�l?�f�G_P���L�̉G�-G^ ��+�'e��i����Q���j�XjɃ6��>z��i�����JH>�t����'`�vԾ����#۞�1=_X�r�fmV��j�D��6�:�"s��n��4�P���x��FP����Z'GOsa��D×���AW�i��X�ӳ4|�mg��F�kU0h�(���a������"�3bx B�@+{�ré�vg�Q��*m��)ks��\:�zGY ��N�I:$��*�9�ˇS�e��8c�kq�����~�g���Vyɵɳ�AI.�E�������%B9��w<�Y���k��8�Ӣ�'e:i��x#y��ݶ�t;gj�?��{�^d���m��m���V��	�]�6g�ˈ��K�N���P���ԅ�乴I��.���@FC���$�h�\]уA��C�p[U�X��)mP�O���;<�E���ٴt�G,SL�@z� �T0�*�E��`���DM��f�bEpj�����Z�����#1��e�h�wXK���D��Ȭs��+��8���Y�4�Xs�%��zer3(/g+<�4A��csU�6�kb���6��A�!��=Pٻg<��m���o��ERJL��D��+\7n
��XIh���P��z�@���^l�]��N@��툧�R��V���0r���īE�Jޅ�|p�,v�1��Mj�7���/)�B@��ݨJ;��9�+A��Q/�$��/��s|t��e~=�߂�W@g�q�C�7u�Y_��V2b1��\�<3�k~�������?O��{X���i,��/�-k�n�,2Ś�(H�C�M	��x ����t5g���M�\`	�Ҹ[�V�߉���D��#D�y����^x�0T������Y��7��{�CZ�o��}�P$0f�E�w��=3�d`休�Q;�B��m�Eo �*ha�@�Q��h�h��SRu�	 eN��؍���8����$Exsd���rp��2&/��E�;O��4�xֳ%�D|�-�+�UR�o<m�Y(e��I �~�|�)Te���Ix���:�ND{����ߡ�����UV�v�)@�Fۜģ";��#�$��v}h�/O4۰���J��
QBi�U��J��"�"w��)�W��/�i$,l��ɾc�KZ�g��2R�ǽ���R�1z旹?c
?�Nv��\��[~�B�|�@VY�2%�����?�J��D��(Ye�-�������³C��'5����6 ,�W���O�bT5��L�sQ����Ժ�	-J  ��
�j��[LUH�x�1�}Ͼ�!�����xA����ǲ�q�D����rP2/9g��pf�&dg�;��ף�����p�-9!ð�S��d��8Hx��V��[���?�`���&",̶u.��\h�K�c��pk�܈?o9ڹ:���h�.FW@���+��rly|u���a�V��\|�Ǵw�|�a��Z1��p���>佩��#Wں�8Q뵟`��*��O�.�ވ3����_IǍ���H�6ɡ�����4��P.}�U�~.����FVD��kI;!u=?��3>\��w=��F�}0����8�	je��{�9x~ɝ�W ��e�1O�b�O�,�a/��+�K�()�����)��Mw(����_�&�O'�h��r�Q6{��u��|x������x��+3^�y�^�鏱d�8��Z�^�A=wrM���ւ��}
%(a/q*�<�sTj�r��-SC��Ce�����Q������h�r���L���';*2jڴ�<�go�3r���<XW�2����}��,�[�o�W-[�.���8��̘ۿ�w֋�X����	iҤ�Ԭ�U����*���&������>ޯ�>B��g��".��	C��f��g]���q����ʢa�`%�y���c���>)J��&<���`hE��'F�c:�Lݼ��H��r��y]��em{���@�;�j.^N�H	�&Բ��EOu�rD�lڔ�'=
Qۮ�_[���'ϫ�kaLr�:�4_S�D���F{�YK֝W��}�t��)N��H �Pڏx�Z�� �SV�𫕍6/�����-��_�tČ
�䭿_�0Gے�)����:�s����A�΄kO���f�¯8T/l�bvHt3��f�3�]�*��Z��q�~�������IE�(V�c�>�:B�BZ�`uC����@��th!�_���h3��Z$���8f�ճ���@�y���=����se�rP*�{fh�d5��ؽ����i[�y𪵴�r��n0�~�j��*v���+�6&�j��X�T��g\-����hCx�޾(�bt��]��@)�&����U����{Ǣo�"�n����,�+�;dj�H)����d*��˩�F�;Ii����vM9	4fW�ۣY*Ï�qD�4�K���c3[������b�ǎ��BQLD�YD.ʆ���g�������@�إ���y��>KG��Y���͗G�­����P�)�K�P*���O���~�`�QHU���t��h�J�3Ւj��QCَ7�7E�sYL9e��/����I]�A�8�[�Ty�����^xN��I���p�xh�!� 7�{���
�������+�&�6 ���]�պ�����^'����l"��o�v퓉V4aۣm�%�8jg�7Tĵj�����n�>�uu\�fJ�\�'�#,=�d�nwh_u��ދ�Qu��C}�P;l�e�h����������2���D�P�Y �v���a�;�LQ���t�Qn�J��~*�I8bX~�q�T��P�kj��./���c4�Ņ��-�r��6�{e���.Q����d�%���hX=nO9jY�_1�E���%�a���^�Z	l��P�j�3-��34�A,8+����Y�|o���yH*���ļn�5"]�h�?�p`#k4:~�C�ilL�N kݣyCp�6v}�:��T�K3B�,���7�� �Sd(7�f�H�4�bJr�EY@.��������NiT�oafc�����v��Qr<�
��)o��6��v|&�ǚ����oX�u���P�wf������R�zS�h\�2����tt��R��`$�q�2��?�?i��Ѐ��%�|{Ό�=
ݙJV��3-) �Ɓ�7�Ș�V�;ڗ�־Q.�b��]O{�D~@�ඥ?T�D���"9�0j�|F�q�<I��ۣ|4 gJ��NJ���ug?cM �(2��U���������QL��fv�F��l�Q�د�}�׭M����w�R����J)� ���^\��ӆ�WP����Ξ[A�w���+����Q�[ǩ]��dM��S�?
^~BU����z[�Ks{�شo�ng����*���*Z(��!9u�W��Bar��Ԕ�p\�5�2����\��oc����zrw.L����F��e�I��Z��S�g�9G�,P��K���7��a)�SI�Z_�ê�lJr�f�N99x���?\
�m��I@���c��\�D�iO��e�����r��`+tL82l�E�?}v�ț��e�|ܻ��@RKI���A���d���ˈ�=q��|�r�)^�qI�$��e����G��IN����s��n\(ʛ�V-���BWD�~Ò�}[��v�(��ӧ�kְ���Ш��w��O��D<�6���|�K�^���h�_�.{RAVs�Lq�M�=��1����<'f_^Z 
���e��}���a%�fft��X��L8[="�"��up<h|�=�4��~C��'���9��]e6��DU����j�Dz�7��K�I��w�{(����e����@�2�������|F���[����4�}�>���i��Pn��V��tT�ڏ���,#�Q���i� �L߾��^�vt?u��]t�������6���*��bL���<to2��Y3�X*���4��&�G��>ą�ꐇ��
%��l#]z�`�Ɍ;���h؁��|���)^�,3�{���UYz�V��rw�"c��v���oc���.v� ���r�#��=���;r���(���H�I��խ���!�s��EP̈́$ҜKڄ���儙�$7�כvi��N�D�Ƌ#7����#VcX�Xq���܌��fN��<#$�]<Ӡ��#�z�����������'5q/��C��YF3v"1�%&�P��Yg�Z�l5��/OǸ���DO��k����f���h-X�� I�;D:������^� ��?��Hx��A��K=Ž�@7k�q��x~eء��;B��r�6��Ѐ�v���U���հC�����c�+�?�	�8��D-_h
��d��-�B�:���~��,�S �.4[ A`uJ�0F���k�*^����<�r���4�v�Vx�*hL(�mu���ĝ0���k�rJ�D�*�L�K�u���yB�7� ��hܔ)�7�}nݓ�>A�N�*�6�9�fJ�����J��T��43G,�	��72��L~��B4P �5�ܽ��6iYE7Q����>�bn�����|�gx�^��mr���QƶKO�%���z��h3X����B�W� g�bH���9���pl��36�(D����a��Q�B�1%��V����7Qm@)���y&ف�,A���#��͐w�U1܆�'{�ak����V]��ϳڰ�
����E���r����bS��m���d���C���A����)蟹��DPX�V�4��Ov5�E��µ�5����n|���D#-I���~ru��=��C6ݱ�ϻW^�>���8Bv�F,օ-*��שJE�_����]��}7{��$1��������9�5�O�k^6,��I���ϝw��\f�@�ʑ�*n��~v�:*�����A��b����$�x�5^J�y�N��1�i�O?���)4񢤘y�'5$;#Jaa��ؿ���B�������x�������ҧ���/���=��k�`�J�>��;CԼ���)���NO�+�Z\�ΕkE�*����hׁ�-�� ��7V>��+����<=?�u�]���H�o �4&p��E����۠�yÒ���&�ەl��Xz߂��7��kS�%	��w��/c�^���w�*�eA.��b��F	T�+���q �*Xy6��Պ�����,�s"�&r���d����E�m�+ϡ��8�ѱ�l��_9�O���G��3$	arB��9���o�}����u1��p�`�hX�oկ���eq)>���O(�����E�'"� �8 �0� �CK�*�'�E����l:�r*j�P�	��e�0G�m�2��u �Dp�6cM#�ֈK����;�Ւb�d��is���
� �v8�
j��E�`[���T��^}O<��	~f�m�?I)�����$���䓛�ᩫD]��o����q�a�
q)�`�܅�!��sՃ/r�35<���'NQߡ��3l]��
}(��.%�KP�e��q��z~d����X�l�h�� ��W\֤GU=m�`����s��Y�7z�߽>�3�^߈C�-4�I�״�~!���׍�<:��><�� �]��d1_�k�Pͭ3'�$ ��;���m|�n{�Y�!οkF
�k�4D�U*V���D�_[D[ʟv;�����EYQ�����).�����*m�l^v��M\c�s����8���W���p�/ 5��6���/մ�K�Όײ]1c��Iѱ$\�P W��QYXr�9oW���S����do��N�f�{��?�ʠ�\��O|M��*��}��j����t�1�A8(��j�7<�2�K�u���{�jm��O��7Κ�Q޻��:�Q�j��B�����?+�佹�G���v�#3�ίܬ]�8���?����NL��P�-W�꾡Dt�� �V_Tۓ;�����%�#�x��dR%��Ҙ�j��K�&j�t�'�[����>��+�I�T���jx�}�X{zdZ���&�7DQ��DimeX�Ho���y�������M��"x�Z{�"�r�m�Q�jrK�I!�<�e�
�'H��q	���o{'9��2qc�k�ct��a+!�T���la���`2O��L��q'k�J5�@�ëdu����]��B"=������}��k/&ED���4�j�7��g9�K,�4���~���Q�`o�q�܇��G=�-����.ES�@2:�a�� �Uj{�8�5)RN�lk�U����Φ�B��7L�5lu&�Ƭ�ɱ���6sZ�ӽjYݧ��p��o��8n����4�闎��kl���
�ڳ�"��K>V�2��L��.�X��H3:[#$��g-�>�,�+�d���������=�b�)����e�S�t;�$�"4u��6����,���
4n�I�e�G�h��H[YӰ%;��e�,�T�҉��w�N?io4��ŕ�r�����
ɗ��۔*����^͐F9@a
�|�����3��F�Z�uv�6d�h�2�B��}:���j�x_���(���?�B��qĐ�$��Zҹ�W��u�K����f"�oģߓŨ괜�QN������[)ĳ8ǹ%mIF=rw�_���ti��嘼�|M=5�q�Fdp��ʏ��/�����5����\�;<j5�	Z�,�;�Ə�Ԓ/���4K�0:qDd�+�p���
S	 ?Z��-������2�`KG)BK��h�2��q�@9o
��HK.����
�m�}K�7n&D��J8����,�>q�}��ę�.9Ŋ���ҥ}�K�{mSr*�P7�N.����O[�Z��ȗ���M
j��iЉM������T��Q���w�ő��v���J� �r�cȁͣf4W��o��ַ�r���v$��J�2œ�t��r��d��lvZ]�4'����lE3�V��@99
ߢ�����uCYJ�''�kX�[������n��E�B�Wr����rz��A��8:nĒs�3<Rټe�Zֶ�>��aZғ�-ó�	Bi���-�>b$���@��.s��������뫫�ót�rd���'P���}��8l��~��;r�{b��д`@�J��Q9���c&J�1Ί����ĂQ��>��h��*���"o�j Xr�\��î�od�LAu�������2_T� �K$�ڸ�2��3[�`ܭ��dW=�aOlJ���}_C�FWB����.r���d�	q�d�=�+|b+������!�\�q7F7���Y�y�8����зc:�D)�mVO�����\t|�쿄�z�!i�H�.ta�t?�-�_���X&f}�/���Za�Pw����֊�%T&A�I�dF��S�W��ts掋ņګ�Hx\aq�~���^;JF�v��pB4�i�)?�I֗�����M��<cD��ٛ��U�s�)��M��佀����%�676�Gg���7�d�Y���ږ���Ω@���k�%���nY���z`� �\�hf(��I���F�4���c��%z tU�NPF�L�B�� �v�9�q���EG/4/��eJ���ޮM�˪���,��Ҝ�8MA{�L	R0+�QBZ�rv9!Vf��TH�τ��q�j ��QL+ӷ
�j�J	���G!Ș.u��5�Xvi%���_�#�Q+��x����"Cd�z��O2l��������U�t�nO��OΞI৅e��:�Y2F0o}��&�gP3��4ԺB�mt<�gn������o��WyX4P&�0��6���ۅ^A������Q1�}b�R]H*�Ͼq3fo�����4OA(�U�$�'�T	���&ٲ:�T��N�PȖ�����G.	QP��&SS�B�MF/T5\WF���k�K��}�6},/��a����^��̒����)��{O���)��9���m:��.�J������+����gn��`=�'d{���Q�CD�ڞlJ���>����/�	������^�!���G���ߙe*AH�_H��i׎���62ʆ����{�3�
��M�̔>��b�
�r��|	q6aX����:P�`�I#1��^�X����E?��f��@8DU���7��`M�v��2�G�Z��I����D��L$�tد�'�u,�L���Au�^�F��5�$Up_3S�Y�9�����ڧ��N���C�����~���iaR��v��M���z��M�if��1�o�����2��j�>��1�m�㮡�F���4 ��P�*����Ĥ�з��a��|L�Y�6:��NЩ��tt�w���9t\B�+ҔL�E�����L��-�����lFvz�X�4��
�C�
��*�=��yq�����x�X��p�JRő���;�["R���Q�ǣ�O���:�1� Gh�F��
�O)k�p�D������J�܊��`�e}F�ޤ2NɧҴ�\�N?�?b�A�����!�'�!,��;����J�g���v"��Db<)o�}@	�bTe�Lq4��a�AR[o�)��@R��W�o:Sʫ�<{ !p2Kǉ�S����:EM��1")�Mr�1:/���T��Ÿ����iF=}9�
Vu>�����!�H��~��*��x]��<���(���y���`����oN��=ޫkN*,2V��]��ԇJ�t�T/mF���Q�cތ�IEFגiYO��,,�!dV�������ǝ;����-�"}�/5"K�8<WRら�g�ٰ�b�f���F=�R�d����}`�y���\êJr�HC��KV��9��Ν*s⧘ tl�q�Su��\bܚ���"�E�R���{��N��X�ɏsKy��A�
�3��5�-��T�)Q�cH
��O��^(Ic���Ǥ?�k�~2�6����7�w@��<%���=��8ڄ��xՃ��{!��Mv����̔�>F��G3�2���d�jP��/MAr����}�4[xy��7����֪TF?N}����$L�cA/z*�a$@�Kgu���,c?�N�<ǰ����ß���@�v
sD���zD@�8E�#aV���M�տT� iZ2]��7��GM�&u�W��9���q�$��"/sJ:���0�j26�5�L��_���VY��y�c놢�VLF��0ʢG���m^W�R zy�x�U�����v��&.�����=���&-�����0��0�e�\?w'X�u� �������n�Ą$T���ל�>���'d~�MQ	t�wN���ez�%4[��1م=��ΣL��Nv�1�٢-U̥rν�&����>X7ƗK��ǝ���/�)�ƞ�ۧMo �Bԃ��2�ǋ6�\
?�&�	׸���2����3[���D��޼��c��5����58F. ^飖;���]as����]��JHz�Rh�
1�9��Pb"���B*j-��S�`(�Uʹ΢�;b�/�"��񈐡G�4o�����e�kS�p�EE΁�U�g1�ɞ����@�A�MZ"��#	3U����u��L��>H]O�;�� 	��C�A�
�������%x9B̌~*d�B��4��9�$�]uku�5�p����p4��/��Pgu�.F�sF�>i.�>��	�n�:4��OL�!�*��� &V�|�ݰ̡�J:G)�_	����)LA�l�(�K��k^i�Y@���41h0�6��h����*�}"Tc�)�c6C��G�53�<T��l��A#�����.��GV+��c���$`ST,�)4�מ���Fj��i�Ih���)��@b�qE���?�Y�~D�w\�4Th��,�?W2�҆Zn�q)�`Y����|��@L�r'��S��I_m�ɜ�q�}��Yv_��2�<���AZ߮��`~/R_�X��W3���z��?���',�D���QD��i�a��p>�=�5��9�t�������8��w��gF2+NVM�m�i����I`�7OΓ�[��j��p(��بg���i`Z\�n�M��R���ds���{$�OӨ��nG�~D��O�9�Fbw����*��$��Ũ�ҖT��o�� ҏ���*0~�ӣ��y�F�ze3��6���Jΰ��-l$'�v�%<u�f�4�y��0�FUC�t���P���z0�u��c�J'��P���z=��-���޶����4f�ć9Kڞg?I��yO׽��|����)�Yל���)@�i�o��+���S�����}zM\�c����	��^u�sWb`�R}��J=�l�����3m����?T���Wm�w�h���Q��N��^������9��>���X�6�Õ�꩟��?�?EP[
�bD��)�c�0���o��@+8`&���n.��6ʾ~,����u)�匘��z��q�����;b�����mET-�uHY�j�ly�s�9 hL�kEaL��
�����2��dEW&���P1N_R��.T�b����$��	�YI�,b��1�z���k��r ��Ųw+�d��{{��UF87�ނ9�a���U�/'�嚣���}�3:�ƟI��Xr��n�>�ߓ̠���:�fV��I3�	���W{�=KZ�Z�}�i<�FP� ) �+򚰅�N�D�'ܳ�^np=U=�*�(�O�O�:?#1��>͙�Jy����@ꭣVN���-�NòE��}T�{ꭰ Z�,2<�q}m�@C�QY%K����|xm ��A�0��(/��=K�L�i��M��dng�ky;�Us6]κ�x"}��ڕD%+�H�9+ *ZAu?�؇D�vˋ|HC�(_p���B�c�<9��M���W`��"IS��5�r�t�Z�ֶ����1�h��أ��L�n���9�N�%Ӟ3{���eM���ʘ�?��q�7��ޣ��p҂�c<{��1�R�U�5[��\ ��t�y;j�{X���8�,�sG�!������M(�����k�U�3��)n�Pf�ま�����{���JF������/���3�@{�])6�����I��୞�(}�8!J��dɝ�����B�R��YcӲ�L�~���ӥ`#{������bŜ.����f���1�ř�e�^�r�������
2��V���X���ҷq��O[�}�Hx�n{�:��£F�����T(l�z�Ty�P�\=~��-_����AM��[~xC��G�u;M�2��
5�JW���'5��t��ИA�u�Ea�$J��Q���C[4�I�2�p�l�%�����;Y>^Ks �C^ڧ�� �:����-@T:m�S��Q���{��9�ū~� �\t�h��R3N��w���9��WO�H�A;��^~�C��{& ĲiDa��ҳ���H�����}�6�pNp�g�]��2�)�
}J{8�ˀ���d
��@:4ML+�7�e	��p�Y�z,�2���qJ�;o�t�{��5ysIR�g�|<�Wo��k���T����;z��H�K�r��f|1xW5�7y9���!�Tf <}�8��q4'��6+vT��f��*0��m� ����_nY~�FF�S��[{f���K���]\UX�RT�ڎ�VT�<���f�?��{����ڳ�m��, P��ģL_RA'DW�CXwIC�,�[��Y�8?gi:�~q�j]��}h+`������T���E��\3�-I�"?N�J%<l�V��Y�\Uj�.(�\;���rv ����/y�*|�����,
U6�6�Q�g�P��"�l4X`�M�4��J�R��,�����|��"[��L� �͛-�� "&ob�Gץ�z�_t�{�Q��l��4�� ���H�C\8�0�g�ݷcF:��=�"�7pQY������Zs�%��층{���*Q�Q��©�����w:d���L���.��X��w��",?B�,�-@z��}E��+y���Z�oH�T{�%��B@�� r��##�?^�<��#C�sqJ_R~���Tx� �%]UU��bۏ����#rk�����Y���FW�:s�4��,�U>�w6��۹�YE�1�!+�#�Oq�hL�CB��\G�9���XF�r���z!�/��i>���ǋ@��ڞE8�?�Jɬ��7z*d{����w�Nr,Jy/QMӒޑ}t���x}OjIZ�OJ������S� rM����-���'�"��c�|	����q4q��*�X�U���~�� #���I�"� 6rW��i���ߓ���S��dґ�����R߲���U�vDmNG4�Л�jٵ%�(#���n|�(|˫�����]�J���v� ��$��ܸ⇸\����������F�Ԕ+�ik�P�H$�\�e����sS0�'��+��ִ��u��
#K�Ƽ�k�|�_�	�L���.}o�����ʓ��V�*�"��tˣ���������uQ��}>.���y��y[ƕ��ж�]U����&��d��l�UM�s�#���M��xG6z}��"H��:1bY�+	�rtO1Z��9��`5O��:�������*�0)�a�0M���T#���LmQ�N/�K�78�Ēb�v�o�x���@'�{��m���M�ɵܰ]=��.��i�����7Ѧ{J�	4j��?��F
�@ y2�t�#80>�q�\4!�#$r�}$L'_� ��a�g�"ɶ�Z��[�b�+#���-"G�$�\[Hp�٘r�@ ���S�OW:�6'�=�K����~(oUH'�ОW�����N�1��3�� &nS�awՙI�����x_f��(I�,O���o6�u��1���QC��	�xa��Qr�r>2+ӻ�m��A�`��&���s��v7���R1;W�a$m����(�0{=��!�Һ�=��:#�w!�}Z�mЧ�Ͽ��0C�{^t��;��mnCe:[�`�]v{�d���n��%����Q�7:3�ߙ|׳^Mt���u���I�b�X�v��Q��MG�:�X�H�0#�'#�B��ʁPU?r���S´�Mk�u��"�hlͺ^�f%_��kg�eI�^�����;� � �C���%0�]��3��6�J��}\�����|��ճ;��1����Uʫr2q��jbK����j����;X��J�o|�g�YFL-%ƢK��3f����A��������SP;:��z���i�U!ޒ,��%��@O����'Ѱ=�����8(Ԕٍ������.�®l^*�(��L��PHנ���=�*��� �V�?��1!�nl��l�3�������[�H�gܒ0�ݔ�N^.�2�<wAv=Ȫ~籴S^�A� �@��<�Or[�۬P�c�4Ї�Wغ�|��4���J��h<8J��G>�i����;������M�<�g�M�O�����,�
��3�(�C��Ѐ#wyEyQ��4>�09G�VER3G�iu��KZU	��_r�Ty����#���ͱ��i5A���M��kY��$HB�TGsb#��=�R�V/��E�n/E5$��.�I*��v0���fH��c�Ϩ1���������NNI^��CE[��Մi�l���l�[f���N�����G�0@�G�R�����Ⱦ 0�\��k�T��J?�<!�$3�ګUs����}9����}��ǬR�I91H䢾��[a��{��/$��U��AL��
�?��6��x���[dI����/���Y�n�G��"�:Јdފm�;gY������f����tn��H	`����h��=ܜ77�0����ޘ9������F���o�~��4�uML%��?��*���B�>��cQ��{��h�<�5�&�F{Q7��v�~0k�wIk��\Ku�>cTACY��y&G��&�[���Z����=� Y�W5��<��Eyw"��u Ǟ��������bP�q�],&���$��-�/�����!fuwy�M�e�*�75�����YrZ%�ڀ��*ڶ���#��C!����'D��
B=��)N�~>NCP��\�]RbI�w���x��S�X�2�!旅����4,��D�Pe]'�b.���r}��H<�hpCf\��F��3m�Q�U�N���@'bG�CN[��pH�s���Ê�"Y%��b �Q����������]����S���EҎ�/�j�f�T���}�r�����7��VX�9T�b����~�Rm�8�+��:���P؛�M�s���ZQ�4|4���F��EZ�*��f�l����z͏�p�4(��������y)��E/�н;���ء��y
^B~2Ve����˽6�LV����R�Fa��̱���b���W�O_z����g��� �����"�:\���[�u��BG*o��/��^�9ٷ& g�{Ay���IDjvV�Ȅ�����u�qo�:h<��&�N�"l�!w�����60�U�W���1z�L=��7��f%c�=�����nj��sC.G���-��SC��B���n<u���ױ���r=�<�I."���'�d�(+Bv����r���Ni����w���D�2�Z���l}r��G��4(���I@�]e�]�����l��R����*��ƺF�
4V��IF���I��3���k�x!Z�ɒ�����BP0��m7"�y��,i��f��
��A�l�ϟ���oz�ar�]���h�@~R��u�%�;��)�>��s{K��-s9�ށ�q�,B�n�iDD��x�|+�9�W����Ӂ5�+4oo��D��
Kd_ђ�{������h�.�k�+U��]���D�J����N���[�ܛ�����_��|2���Ʃ{�F^�e~I2�xe ��!z�����-�R��gߊ��UF�[�g>ᚕφ,�0�7V=p�hf;p�G98�ic��Z�W7�:���~c	�bz(�b�;9�F�wĿbγ�AN ��{Dߴ���Æ~x��m��d
l��cW�_���F�Qcc=��2I��Ut�0����4�?���'�Ҧl��Aͪ��Zbs^���=��Da��B$u���\X�κ����;`��)��z�;�A*>>���R[�!�� iд���:"@���Eμ{�2,��*�E���h\i�	ݦ\�
t�6?�<V.i��wK��^K����"5�H�>0���ԫRu���!��T亟���ہo��ދ��8�XW�q�3�{��yS�h���I��dH�	vS�l�� ��	5���w's(�8Hz�/��K��?����s��C������D���~N�o ���d�:CS��<�X��Ӳo�j8��=��&{E+P����4�c2�b����-�'�_�Y�Rj��,����e��p���_�vw7@�����p^�C1�s?]Y���4i"�R+Q]Zy� D'JΐN���O"&�ҽ��șǟ��<��W��p��x@s�Q ��D(F�:�+Wj�}����~E��p?B�Z��l4i&�~[y��Oʏ U��.�e��!��X��@��-�Da/@l&�V~EꈖV�.�y�~7�l9WP��8��g4W7h%N����S�<؏���SO�t�ǵ`{~�!��`<�jz��V�{�RG�
��Q|��5s*��N2rkձ�6���T>�2�uІ���ɍy����+;�ϣ�<�c'�#�h�n��f"f�C���H�%�Ø�����P��@���κyb{J�	��a`��m:nWQ������������q�'{U�Mb��]Z���f�ŋ`�
�KL1_%b��:����&��n���W�9� JU)ޭ� O�ÀkC��{��?:N _�ȃ�g�;pi^A���W�Hh��d�
 #=�"q9�=�y�I3j��~j��Ԋ��#�gۋ�$p-���<1wS��>)d~��a���3_�N1�1A��B�4Y3b�*-�n�֮S�C��e݉$T.y֜���P2�xU"�',)B �8�?�hV��KS!�bP{T�������������m��k%��b�������-���hTO)	rj:ȃK���$���������{_D�A����$�oPl��"so	M�)�2�*�95�X��.5�q�;��,u�'d�#�(��%��J\�X�N����k~4������0�u�7"P�9v|�!"Tz'�V��]b�3���jn���Ì�^�QNB�Ã_`��$��F �׉J��Y��nG��9�g�	n%�凊�wtY-���N��h�<?�Q��M&��NЈ5v�G:l��v�
�˼�X`�
ޔ�R�r!��a(�:�Ձ���:�\^�G_�kW�o�F�--Ȧ?����!S�v˦7�#U�K�YFB�Y@�Kn�ΧcS>1D9X�н{���8{[(��jb���3ZZZ�����緾d: W�%����َ��HV����i��t��D��� ������O��a�%�m��]E�.�H�;'ª5H.C���L�n�T��6�sK���\?������1�hM��0��<�y������"�vx.�\"�Z����ZJ����l>f�~(e(j�?�.J����V:�u<z��{]�~�QZ�1q���,긫n�.[>��Փ҆��M�7	��`ɚ����x/:q�f���f̉�|�(���M~�w��a���m��@�qm��|BT#�A�ӳB��(�����J�u]P�#�w�Q���1Q�d�|������k�&5(�k�TO���G�kf�B� <�X�I�]��ܬ0ȏ.���U)�S��8S<�b�2���k�k 5�/BH�+Ŕ�쇮�o_�,�*C����!`~����#fC�qL�-~w���w%꒮��������h憍��I�D��Q�/�wy�P1x���CEI��ν�6����	v��g6�ʵbo��������q*�c�nյS��"�൦^���Gn�K�N����A��	' #�eSFi��"��S���д܆��{y���a�.��p=�D7�J����7�B�1����L�&z~8�Ú?E�&�ąW�-lF�D�l7�����c�{ ~7IT�
X f8�r��0%�8Ι�g�5�i�?�2)�&Pr��ݏj������0���;��rK.�(g�������4�(Nu}t��Ȕδ����Ӣ�t�[�͐�C�x�*����%H���dbF�q�	�$EP��~G"�R�XC~��[$�2���l��s����Ü�)�&�뤀�j��g.&�r���.��I}��pVp.��ʡ�P��U-��"2�7��|����J~�=M�8�\��H�wٔ��v.:��*�r�o�W�}�Ϗ	Q����7i�Nc�|O��Aw�ICe=��P��`J��#�p��� �ٔ��0o��� b���>��	�e�����b�C������^�{��gaX
�ϓɕ�`�;��L�����r��Y�f/gm,��.S�2j`{?��´�:��iR�A�4q�p����$�M_aQ;x���u�r:?�&=�U� ������Ԅ]�e����$nG���K܀��ӿ]q^��Ƃ
�0n$�<ִ3���7HNH�9̓h`������jzm�"1.?~t����� A�*����ߖ��Ya���e �
��<��hj���΂��������ڡlC�C7�-���ƓTSY3��!t���2�\�
H��4��u���9�bmS��ˏx#DNڃ��XO�o=�o���Y��%$	P�IW�7��a:!v����ݧ`�~�DӋ��7!)�ƱÁ� �Γ�rjS�w⒇��:�m�Z�������u"]V�^�Φ����b;~�=�搵��Cu�� <ٻ����8� 	��n�:�u���>g�ݱ޲5e�x��)"�),��XPq�hb�;�� `���j�W�&��y�I��_+��3�{�l�D�G��},09>���!�\o@�	��U���dX�Gt<EW��TavJ;r�9�
{$S��D���F�����wC��=��FO$R�cm������D�&H�u#'f	�K�r���E���_H$�-�qL��y��߅���-��m�ꪺcc�{���d�G�)�,�:e���M�\;���A�����}�d���ei> �)B�p�=b��*l5�R��q�f�7���O���?�Y�̷�������[�%϶A�Z0�I�hz9z�� )/\	幊���`\?ees���z�'hF�\�fc����D��I����4�9�K������t�f���^)˰a`W��cRE��@U{� ?�c����"Q��q�c�f܅^C��i�=��t���lbs֖$[V�f6��mٚ�*�|��
���}�/���������p�}�����ln��b�3�nV�i���
hH	�~���C�vyɒۅ>��y��}�SQ�~�ĦRL���뉥as�9J��\{7���3��y	6��)c(u����?� �V�:�:��9��%?�����%��.V���qGVGv�dٻThߦ���r	v|'������ţj��P�6�}�<`dK����(U/�#����w��0�A�ű�}T��Q��O������+�I��B
7u+*���cS���in=`|)*,�z��N�cLYDa���R^���^�*�QJ�(��Uj������uq-� ��~em�#�����%�����B ���+>~�@oV�6�̾�S������F��t�VXx #���5*8D�����>i��E��pdJc�����ɗZϳ��� �2��V5`
H!d�� `r��.���!�sgǓc;�P=��XC���Xr�b������ίhTF�:	c���V�~��ڪ��.>E1��(���/z!l"���iEQ�SxqcsԒy�Qc�.3�W�x;�q �±,?�����s��\ZY��d���I'Ł�����_"^�<~2n��������zE_���Lfn^4���@E#	.�rIP���rq�C�2e
��e5P �<�:n�:O;g�'��P&�dB���5�Ż�	%��<���;�����E���~�� ��kReHQ��.H��[[����I�N����&o��G��<ݛb�*0�!���,�A3��������������;g�����FЛV�����:%�!�݁���w����J~_�ޏz�3�Q^t��$����]\]M�L*GU��Q�Q`I�%J�	,�"~3�X��s'0��A�|�q3a�� V�lHu�'��<����f��`�tk���r�W��X[5��>'�r,�qW��d</��veMU� �̎��h*g+H���&z}I����%1�V��҇<��.� )������s<K����LT�ZZ��p���p꾔e�5������X��Ks�1�Ŏ�w*�H9��m��F�g�>1�#���P�P�6 ԛ���5����]�n�2��#�I!�O��\}����l>�������,�g��RN�vc,�'�rb�-�;\l�4=��(�_�*m�kM�Vc։D�k��</�����g�݀�FY"ә2�Y1s�t�3Ct]q���
��Q�|��ݶ*<��Z�AL/GWZ^&�[��� (P+'D����k�t������ɜ^{S���=0�nq���iQ~��!�1B8�Y�
���_���;1�7�㌬"��XV�~`�@�����K���rr\	M��U�b@��Yφj?�ڸ]WC5=Y�1#/.���j�N�����;�~�h�u�j�� �J���{�A�߻n��;x�S����?!�|�����`L�� �?aKi};6Y,3����G��\]V���j�3�L2(����^��C�*������s�Hh�ɶ�3:��:{��G�NE1���6������"L�oH(KhpL"�Ҡ%l' Pv���FJ��
��Pc+��&͟�k������e������]�_���:R˘�sB���{��L�����b���y����G���ct��d�\�u�aҰt%$�R��������TǧB�@y�cUL��F��.����?'�ڈ���t��P@���u�,?�2o/���ȰHr����|�O;�ՇV X�?��{����!'��gD�i�h�E��M/RKm#�o~G�� �uG[�6N [ȥ�,��a?h��U���k:o������_�8�R��T�����%�\�wh�%{v�<A�]��ς�\-��[����M1m��m(�;! ����F ��˳�B���Ï�r���o�'����mZۨ�-5D>��k%ȥC��L51#ˇ�F)�^:���B��葕��,�%���aD�l뽸竜�s�˜�s"�U��r�L�!��j���){�"�ƔY�yS�VԐ�2J��lVŻ)�(��� �'ڇL�����CE�����`�U�lΡ9��.	��{�]ʳ�R�TXw�ś줴�Ĥ�H�&�� 3�2�IŮ����"�_0�\�'(@!~�Ȳ<�t������SyS
�M'��{���u�m=����2p�ZA���m|���7:�?'A��mm������RBܱ���ݶ����_v��T�|�9&�-���ך�����w��V耔H��O�7�[,�k[�^n����}MG�|� @���SD�,�����G�\n�(��=�Ԟ�k4�m�	��Y� Q	�KܼQ���z��s(ED��΁GĨ9y����oZ���1Us�����i�jE>���eh���}^�4�=�r ��q�GI�\G���Gt`����o�Ya��j�{�LJsO�]��D���mA,��юc�?��ay�Ǳ����J%g��./#٭������1��ʹ�}����p;����+t��O���.2g#�7z]��2G�u�w�K���CM�0. �8�l��믁j} yrAJ�����@|
{�����p�w���d�ǡV��zrpF1� �����S���ݪ��8�.�9�>�F	/G@���HF{�ǘ�QC~R��������([cp��pk8����ҟn������G gn?8�p������9�l��e񔰬3�E%D��X�ZP�C��B�O'	0y�C��uJ$�K�f-ʽ�+���S� ��+,v1(kз��O�"7�f�[�z�"��p��T����}E�l�S!G
��]o�N#�f�)��K�Os_z���F5��!���)���K������^�C��&�������k�?��(��l��M����E ެJM�o
��.�_d6��į&�Ln8��Tq6^�7��.s�j2z����n��������>`��c[���D���?Y�gQ�߬��0����.]m��q�|CM��](���e�I�����>4�+�y��*�[?\
8�[��N�+���Er�y_��읽���3��K��i��-��R��ݎ���^[��:C20L"���:�mKx�簇h��z���"���4^��[hg�!�3"8��d