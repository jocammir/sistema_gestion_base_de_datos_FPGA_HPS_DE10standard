��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��Nڭ�	�����B�#Z���?�4�j��0�ΐz�A�y�[��I4�fB���_Ɛ���-����B���M'~��k,���'zf���]A�� -̭���ҧ���D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0�������c���Āu�T��Y�2d]񜩳������Ů�e�ɤ��kyǉ���7��B�p�������	�≾���*�D��=3xn���5Zh����	6\�>Zs�}�K���i��O�|��>���BD)rQ/v�=B���R�ru��Ql�)�s}�w�sN�NNK�$Ϊ���I��V���Qzs�<@.�$�x\�ȗ�����?��S���k=��-�j��j�
}�| ��.e�e�=�P���Y^��:&�%��{s�{Բ�7�z��^�M%�u_�V�� \��{�\�RG;OS��'ޱH��5WDi���+i�'�Q��������Z!P�O�}��Ս�Jl��ڠ�Ǯۺ7�/�P<�T{ *�I���\��/��b�F���XÍ��~ƄXN%Q�%ҽ��BŦmD[��Jc���y�Ʃ�)��ڥ��]����F��!�k�,
�֢t��h�2�����B����f�N�9[�b��9I0���i ?@xɯo�@��<aW�E��8
^	�uW��G�Qr�Hjl�	��>�=Ă"��2H���*0���Ny,��U��!�:U�U�x���?��ݝ�sU�ceF p���9+�q��0e9�y�ϣ��)��U��!���Q�5n$H
��u�}�w�'K\ӿ�V]�U��IM k�s�cZK�p:qݏsŉ���#9'?�ᩎ�d�cч�A�:�P�(�V.�}Ļ��g�y�JrSV3)8W�S�&A`�=��9�
L�9#fkx���E���Q%?��z�i"(NQ����9��*��Z��$�T
e���Ca�yW*�/6Ϩ�O��`�����P#+�*��'�D��v��x���g� �Z��r��6ŝ��٣�)R5^�z�kϩ��A������<��ީF�#�ɍZ@ތ:AAa��@<e�����}c�ks.�8��,����f�%�Q�x��g�F���*hgAM�$���s�qG�oy���#�K��i\N(�J$c����x%�5�03�&B�`�_���fw��%�vp'�qx��v�i_����x%���ZT�P�L�\(�Ǫn��jJY��S��9̐�@� �x�O9�\�u���-`Z��L�>囹��Dt����#h*�ݳ���Ղ(4Y�H��Z��x��3^=��==�����a��P���@�,�UPek���pP������]E����?��4l�|DtZك����,׊�)Q�R���5A�4�ʵ�hb������qK�e�[��4�-cT�=]�M�+2[�P�f���1�_UL=q��1->�*�Ӛc�p�7�5�ѿC4�>����c��J#�,���<)� �Q��O \z,�Lg�C�Xʭf+�{���j<
z4.���eF>��f~M�f���*�А�ύ!�g��5N3H�s?��LBi�ˮ��\�k�G�&x��3g݌Jڳm������qK�Mq7#�8�sOȋ9;ǦE��7�ӈ���1��Ћ"E�ѾG`��#m	��h�H^�0 zO%�1Bo2)<Ky��gB!�-�Q�~ɿv�
��ŵS�
�_����s(Ҫ��옕l=�B"^,/��x����ʂ�"f���n���K�&������2�H'柟�~���cЀ�'�,u�>��]�c[�E���t�?��M�&�!����:'kc]Ed�,u�,���ѽ�{Ro�\� �F��&Z%���hb��":�)��(���瘶��釣e���|�%�)"v^M�2KT=H���:�x���y�v���_ҤSE�M����Z�O~�ϱ)�Ii�-s嗶�O�[`؅i�i�O�;��Ȥ����.�Hj�x���Տ�/�ڮQIH��:��o��.���;&x��K��K�J��3q�3���<� "���d��a�M�ɖ���΂���r*���x�N�b*/�˺Ȳp���~?0�A<螘L��?=�����M�$��ɥ�&��B�Jj�q; ݆pd(:g�{:�[+/]���7J��KrE��x�ܽ��-"Č��'�1��.�+[���4Y`��Z�~���ț���	�.(>
�=�KS]�z�N3�J���b��`)/;��c�d�V�Ϻ3�y�`�>܄��\�d"�w�V�!���ԂY��j?�./��}�Δ���pH�'-�G�K���YU�H��Հ^(�-bW1	fT�Q�-<U����2�l|vsUH>�O��'/v�ح\��=GRF���ܵ�S��>^n��"Z~�ڬ�ѕ�o� �F'����x�?F�ɯX��c�+�8I�[���)�M2�O5{�$h.(��r$	p�O�a�.���[�,T~Pڸ��g������V��ȪI���b96����v�:YFZ<�A�n�q�.������K>#ߤ� �����Dc�YRL6�P�L�y���0X���J^��e�X;g�Z��F2|l8�$U�1o�B�����C2X���1��*6iq�F^Rz�^uk��6 S���ݩ�Z֟z�n��Z�%��B�Ҫ /��A��o8IH��K��Q
���Q��n^O{�Cy�?y�׶"�r7��IX�������jl��q98�����<�8�R�/�6+"%JU-�)j�@����F�(�?1�c����s�(�����0��F�y�X�������M��`lK<���FtZd�}LA�=�b���{�v�w~X���;K�J��x��Y�P��u��a ST��_�$������"N/�D2��:_'t�(tz^uS$���4(>��*A�a2�ǃ�dHxJ艃_Fu	vjȎ�!��i���|�`Z�(&�����(DYnN���dZ�L����-q|����h��1�Iq����~D|/q!淨��Y��k�a�`�Rڳ�8��
C~lq�89uԳC�nI�`m5�\��_-jg����0BZ� ��THX�'W�(��ֵ��y%��p�O����A�e|��'�U�F*�̉-��T�_�&�)ECz�{��震N�:/�q%��A��Y[�*��F�A[�u��me���u�����=7��)a������Z���\Њ�԰�f?aA9n��9qM������,?�!d+�A*{9�,$�E]���pܙ�A8�9�� ������&��25������A��ޣ�H.��=�{�Y����j�hi��r<K_�"ps�(���t�(Dx�(�m�?�������~oݫ�?����?��U�.�<���RL�Rǻ���m2��^�x���0�ڄ��N�8�!&��
��=�;�|�q@N17���!�o\�t��Fv��U��?�Z�n�B��V�*d���0�,�@�BY|��d�@:��ʊ%�@��K۲��'6���y;929��}��W�?w��3��|K.>�a�%��J�������MP�0���1�Ta/�48�[��v ��![.����s���g��g�Rv�D� ���\�wA�i�P�`��78��--j)�4h��,{x}��c�����j�UƝ�%[w��F�&��N��e"6
i�շV��iv6؈���j��d�wli��ه���.x�bE��0�cU���S]�P��9N �}.�0����y\1�.��ۮFR�`U�a>�|Is�x���`	/���H��qߛ�< �j vd�+�|g�1��B����I��^h-F�/���ܼw�jH��0�P?�.j�w��?���~���Fvu�>�J�ΰ�[���f���(�&E�FF2�;d������M�&���?��j3�4�E�]���DRAM)ά�ۣj*��[r��p�K�l�9�ڕo���~n=�tZ���(��q��>��J�5���*pOe�ޭxhޜ�=ϙ����?�	�##�Zr�R��n7�a����^E�����1��n�>��d���$t��t���晽�Ai5'�oY��8��̧Ch�?���Q��w6T�	�Ѽ$��'/��'�����% �{9��R���n
��gy*�h5��=Q)rg��.�L���gLR�c�I��$���\�u�I�ey�(��>^�d��_wF�D�(W��[�fi�g�Or�&�Cc�7�X4�WK���!4�nR��rpf�L%�?�}g���=/{��bǴ'|jsӍpX�C/�Q�@���$*�����51@Drc)[-�`F�-���&J%G?��G��t�7�9}�# 0�2tK+s%b���g��	J^�����%;C��?�)6���	��3|cN���93��`�;5�-�<x�G�.���&��(
ʀ���%����w�@�L��$c�b���Wҕ���`��1�,�X�M�6�����wL@dV�1*�Ӳ���RT\�(��s�x�WǤM�����Y����*��e<���������1�%L�4y�X��c��>z��Z&����M\��&h�%�э�����;o�k3�m�P�Dc��q�����^�U3��_�!0鉄۴�����I]h+�Wjf�`��|��6��1O`y��\�q�Iݟ��3�D>��>�f�@�g�������$�_��W7s���(�g�L�i���E�8��
�en�6l�=���s${w���죰��&���r6
��y�w�KS�oB��|�.�	�A�O�v�����5j=���W�/r4h�dx�pl'��0�O�!��, �)�л��B�(��ͅ���6*:��ǣ��]Z��vO6t��m�w ��T�I�X�x�e�nV�#�@��5�S�K>D�v��0:�{5��|\n�k��6������ɘ�e�[�{½�r�|@'�A�� y\�(m�X��2ttX�Ys��-f��F�X�dW줭�,Tb��wb�+q��4 Y��%£{�Nۏ��h>�%��C�;��/�������87���g�*���5W������әڋ��BC9�T��3
�ĸ;���P��f���˟=J�vcC+���	$�
mO�Ǘ�H�A��px�,/��E1�}�׏H{�.��c>*O;�ֵ:σʂҒ���t~�M0:�~唰9�ϢY٢*q��uͬ�&�����?¨�C�>�G9�����%����ݧ9z�VV��𩜮�Kkb��(�.ο-I�\L��Zp���W�ͯW:&�^w(,�l$T!��0�]�]��|���V�w����QI�)�}c�}�	14%ا��pe��E��ΩL���^�/���U{K�2��PX嘊���ݏ�6��x耒�~\�A��n��W�L��L��(��Vy��b�����ku1���оn^9������i�+(����_��Δ&��(�kЁ�]w,�}�3�U}4��.=��p�!�@���Y��m;D
V�X{W�y�E����2|	�wc���0��Y��t_Knp�M��:d����+5�Y8b8,��o�v	���.����qG��܃)j�x2���&(fC�t����3ger��p����bW��_�ZZ0�3Ȗt�{��� �x���`t3� �,+΄��?R/MHN�]�F�y�Z��������_�;"O���6�>?�[� �_��ɐ��v��솺~s^B���l��f��A9�d��P�~�\OD���%��M�	G��'xdxXf;�w�I��V�z ���r�cD���4d��� �-UG ��ٟ�C�0�J��lN{�F�5�X������,:����J�D����3�ЃJS"2��^Rw/()FԼ�����+�S[����O�F�����WN�E�������sd�;_�-�O\���?�;�j�")˓KB�+���t�{�I���s��Rhi�+e<�h8�Go�@tW�k��ɬ�g�"�W*�G�����~�п���i��~VJ�;6�`�0�@U�b��%�AaSf7�}�͌r��~b���~�B�c�]���\��d�r�$l��)��A�4��|i`�б���?!��qP/U!^��5�[N�]�z)�� ��2�'o9�mL�����&��gf����բ�8�p"���`m��^�;���F#�Q��z�U�U�5̓�V�V
���^�rGT�/��C�bȈ0��/��<��_)sOl<�TG_gT���W�,Pn��(���?X�v�Q��Ǥ×�f�yx���,09`z����H�E)�B�q��a?��A����Xy����;�b�M��&�`r�}˼��:�SȭO�]��f.Pz�7Tqgʇ���01��e:��_���w!��w����\�[<�o_��[v���g{�t�����٨[�y_x�}��#��a�-�fgpa�mr�~����E�ݔ�b�~&���?�,x�R:Cmc��l�wAAx�&"������ ���V��MtqrE�$O�D*&�,"ہSB|���єo�``�V%�J,(th�;��h]�QX�;$x5b�+������u1�ݎ
�G1}���7k?uv�pP�T�.�y³m�0�R�~��cq�էc�ɺ��&�Ο�$�|w$R�AS�����p����W���g���� ~�[�`
�����k�z���wXA��B�.]m;�:Pe-�z�Ԗ�lvq[#aq.ǥ:�'T�0�b����r�a%���e���M����l��a��Az��ҷ�W�ӼV��
^˄�yO_�<���i��ն��j}��=D�W��h�ݧ=:�z��r)�5H��\,X�º��7���O�p��+ ����'�
��>�
�>ˑ���U�<�w)�����m	,�%="��H;�^⁬M %�`�����᭧G[�@b�>�OH}��:�4	�o����}��l�`D��Cac3='�,)�.Ҷ������
eL��t�� ��#YL��/d/��C����k��B�m���մPl>���T/tǦ|��0�)����,j�d��M��6��KV�
�lܗ7)'Ӈ��;��`�d�0�~���!𔖙�K��5�2:O�~��恞I��H�,�ީ�S!�����e�q����Y"������/��KP0L��{��E)�#~�`	�r'|��!�RMV%n�/�w�L�d�W'��H�#��K�[g�uL&��6gHX���EDHe�a-\�<���@Zu�ə��c4��O�^�<V~�_D�L}�Ca����-O�F[-�ގ!X`��T� E�P,��+�Zj��9��`�I���㨚��it؅JlD�hOV� 1J�8~^�Q̢w�G��г P�J���j�A����Ǖ4����?ԟ��J_��Usw�v:)�k�8k�ɥ}'i_q�>3ͱ�����I7SP��V��M-�,w�Bì�
&�x�F������3��@��Il�?��M
��%���gw	�ȨK�(}�p���;��h@T'VYB�*$�1zH�3��o�[\�%A>9��[r:M�� ��G���ǅ�0tr�����%��h�N��sʳ���P��O%O5+Q�B��fw����d˯}Hl5�uH���c��l��!�5��>=�A��b�5����3}�����,�3���{�Į�v��1�� �����M��Rp��}9�-���ܸ�$���Q��):;��?ה������&}?�'a�c�D�pwo�D�-��a�u��S�8S�;���;p��'���ox�B��瞫�^��*r*�Db���L�D��|�Hge�ܜ51fF|WP���V%�@�:�����ml<�������`_�zᩪ�V
���}v��q�A\�%@��?Hb�!���߻�_$��ϦyU��4!�z8�>�C�1���4zK0{�>���rI�l��
X����aץ]��^Ik`����)9�s}�.�E�\��?�c��c�r���œ�Fxl.x;�gZ����OJ�w�=#=�׫@f7���?�'�0lW2I�uy����ǩ�d�)��' �wC}穟yʬ���vB���*�]T��xʫ`Ȯ��M�s5�O�,�/�r"�����S��lkuBҊX_8=�� f_� �WL�x��y�ߑJU]H���;�*O�L�7��.?Y�H���A%���R
 T;(�[�M9U��'��hBs�>����[/1�dѾ1�9���-�<�FV���u�e�^�Mt6����<��y���O�iOQZ��<���,��)R��^��2�~�^��/^��E>f9"4��WÐΈ�T�5e�鸈���b�7_��I�4~�+rt䘄�l�dƇ!X�pM7�Btx��M8�-?.��N<t�΁��90k�-w$v��#�i���#v�_K��
�M��n�i�X5���Ρ9��I�yHN�sɟ�W��f�\����@+<+�~�(���D��)QqA��M�]�{Ԑ��83ޱ_�}ɱ�4���5B0�rԪqn�W����mO��#�,���룑0BS+M7@��<2]��H��$A�ӈ.����Y�hH�P�D=1?�x�ͥa�2��L"�wh�� �oAطI*GB�HF���*ưR������m���b�f\o�g�K� 2؍�V^!���LG2�#����q���N���/��z�}��z(}D��n~�V��
	&Q��3g�R��Pa�g�k�f��'���=�^~"o��O-8��W��#�L�-���C���M��f7�q�X- �mr�}7W�Ǡuю6}�ڳQ�R�����vZ�o,��1מE����/����%���<��x�y8�����I[�$����T�o��C0����l��]���ܠ66��T(���%2O�=�D���gA{�X���@jK��k{P�n!5�抔�K��
AH	�T��@��3vl/�����&S��������Q|��Waˁ�$��kbef�����M���l]@�&�EL�
WKTzf�y�Y>V殴�*��OT��Ըˢ~��� c�W���My�h��I�R�"jT�`�Hs�Rͩ�#PT_F���R�6�%���^�cG���]mU���o���>��~�ڠ������,M*2Hd�8����Q�!Gɡ��#��Yk*���)Y1�JK;�����F-����̶�K�Rm�x�.��'��#�� Z����ʕɿu�� >��M�^�7�=����]�
S[<��Z񮀋����x��Ċ"]�g@���1�ݶ�G�� ]O�x�eU��W���3�J1:˹%����!2�	�������.�E<�@��:+���ܛ�V����v|
W	��D�L@�[��!M���Փ�l�C�?���&�@8Oٴ)�D|A��I�ہ� ��ϖV��� �ލ.w�J����S�0r@��%������3h�<�ɑ��#E�n̄�;�~�As�A<M�U�)�{�%)�~��FH��
�#6f!�	�݅�0�v�-�z��.���c�G�%���S������W�p�ɭ�N{1���i��%|�}�.��E���HC��r-��@_FO�.���A�Z��=#j�δ�kͱ�Dt�ʑ��R�*=j�e��*��N����L����i`��6P��:�@2�Qf��&�У��`��-���m/	۩.T����p.uʧl3��:�T��k3������h�����fk�/��٬�Ȍmn�������bH����b Pbf\ *�z�m�r�)�Հ� �:	׼���h�'��S6������X�C���!��2 �E�7���}fv��c�!����� ܼ���B�Q������X[�ulh$�2�%ʙ�眔�d������$��>\adHQ���m?�}n3�[Y�=~�.����o��