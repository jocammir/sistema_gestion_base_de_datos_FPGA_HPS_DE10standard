��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��ܼ��e߈SU���AR�>+�y$kgG����)!"���S-�e�%]�gf5Դ���s<G&�,H��gX�
܎­SH��76���kEb���Z,��O�\��X��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�s^W���0A��T�B-z��=�V1j�*^���`�����'�����W�����2t�G>��,x�\\�\�� ?�ڍx�hM��H�Ə^�1����۷�u��zg�Ɽ�U2�[m���I�aA�X��N��A�7%�OD
_�,Ӕv�\䗺S����%�T~�6�ѥ~����lj�z�.V;l�	�#�9���dh�������Z@��~Ǝ)����\I�L:���)�`f���f���^
�����<~�	�2@�?���mܛ�7;\�y�g��"���J�m>حj8v��R����S+����6bAxRN>M�u��V@� �^�Jȵ�|@w�(���²��_�E�Q�S� �+�I�Y�:���'���L!�(�zr�Jɳ����~�<(F�u�}:�X���Ŋ60E3\�ӧ|�oP��O=�peRP�0d"aL�������c��<f��Ir��$��Q�؜�&�M`�a�Lx?p|s�;A�{2
�|M����ϯ<`�(}�$k���F��3�2��$h� N`�T��ĿX�T��dZ�Tmoު�In�5�r��@��ԭ�l��@E@��y7l8&�*=R�i#]yxV59�����5T��<��-�+��l9�~�'�踤�J�Q��{Te�\h��P���6lgd�s��׸�s��"��"�%U�A��ǜ�J��H�@�'�,��Y9�إ��5����.5~�@��[p�ʘ)v�-������{!�T%N�+hd�@����\�B��w���i�aV�����6�nƠN��<���&�eEI��;�}��gB9z��a�ַ��u��fQ�Hz@��';��/l9��b��t}Ue��uk�Lb�Yyr�Ώ���RiT�@�)���Dݷ�>}*�;p_��#W}-�v\�M5��x���-�nWm��m�4^��HO�[x�����>��'���3�%S@��S��ꈶ0�[�����u.�`�ͫ6\��X�=�sEE�w��4�`�H,Ӷ�l��B )�iXM���>��\��'��*��R���N��'�猍�߹�yp��IJ��fY�RzU�O΄�Ww���ܕ ��V32�k�]\+�N0b������z��]��5V_gf���z�,>&01(�/�]���͊8W�c̓42"D�!�^r�٣$9�4��;�G�Th(��t܈�wO=���{9�X�V�e@�^Y�bN��~��+cƜj%LIm������d����g]��9Q�7�& �͕Z��
^?\�x�œd&#{k�����0웢�p�`�KZ"Y@���)�� ��_v�^��*��G:�r��c��/d�ٲ	7r�M�Q������&�������2H��p~�����3��n�ҐeT~��d'�YT�Y��s�T!�oe--3/�<�Si���4饪��i���V;��@t ��ntO1pPݵ��b��Pȝ�������V�2z�77�WB!�3�ն��#v��^�_���B�q��L�2l]ȳp�+�.���{ �"<Mc��=s!ݳ�8�Z7G =����I?j�?Ł�߀�e1���󀬝jd��5��4BHJ���NTp��{� ��=�)x�6��������*�͌Cr�HSn��Y��(�S���w���-ne�$��}9�n�'�����m�ϒs����s�'���1���a���Ũ"4+��q�B��vOt�s��K�T�i�\�A8{4��eiZ�^�������5UT1M�#�S����PӒ��a�V��V�&W(E��-Ԣ�c��yOuDm��X�N�pZ v���@�_�pd�:��+:lIwqq�^�N+����� �Ts�g<韠����A�z�ٞX^�^��:�6\���@���ǿ�EY嵒y��	��rH�j�'Ű�h�TX�Ā�?VgCu}qͭk����LP�\\�k.����@��� �URp�6�A9�ٞ�K��X4�Sa���jj�1��m���1�$R���9��r>�-�C��-i�D}��\��w�(V>8��Z3�3)�sYE��̰
ģ4��'�r��͂�L�Q�w��uD��Z)��<ה��n��<�K���N�ٺ6P/ј@����U�� �:�u�m�bgwQ��������l���2�}�Y=�Foő�ĻP(E���������z���O��k`�Њ6���7um43�����B|>��+��FV=�';i5���~&�����p����ɒO�U�ɻ+�_A]���cQ�r<~����^�ɭ�叇Z��&�,��ކ)����1���?�M�t�
A�΢��-��QKD�m��ԝ�"�"�n�m�CEd;�[�����Rk(E��ܚwh�`i<��� �jGW�WY����N���4���s�z���_.�M���Q�TX	�R�$�,&ϐ�h�Y���c�P]=D���	~７�q�O�Z23G�}�Y�L������TQ�+�а�K�����е�S�p̤d;�O$�]渧��y |0L��lkU2q�.�$\'���I��z��=7|�Q�G]lK�J*���E6��V�n��<���Qr�sΦ��`��6]��S)�+�\~;� �9hRF�>�5F��d����.���-f��n?���� >�����pF�!a������`����.��1�$mNt�j��[d���U���ԦfbXq�k|v��>2��1 ZQ�@AC��6́��=<h�*��.eS� P�z�pn�.Lą��[��8gG�*��	�r��.7�ʫ�k�4�̺���l(� ��.i��AT���`�����.�ϯ`�sK֩��S]�iWl�W�X��79�aO��j 9�/���l �m*&���h�Dl�.���I�W^�V~(>I~?�p���c�������0�ь����Us�l?W�P_����ٜ�]��|-��O��$ !{0g˓Ky(�O�"��u��w��;����`�+p�@���qlp����X�V��C�z�瓱s�;��(�Q��9糍�ab��]��s��	q�Y!��1mRA����P�S��L����R^��\KB��(6���_g�rm��v	�T���U�3O[�
�h���1�����F�ӧ*�1�!ӓ&| 1�����_� g%t�@~�ߚ�yT��^z>�0�C��QxTk��Tp�ShA�ڽR�p:��r���ё��Q8Xd�}�ż->�xз��d�BЩ+��N��CE{�lP{��}A�6�B���p1���H��Q�LΟ-�`_�����
���>W�6Lz;��5y�P����*Q���p�[Zt��?P#�4�K=��C�N��\��xk"�R>��,r��	뿻���ĹJ������ z� b�z�B9��
%F�7Мu �c���ܛ��(U;vbq�f-�,��+D�M�q����l2�B��ā�T=�/E��LEd�7��z�ap�R��/gn��\���]0Ue��͋T�paP�;�\
��.�z�K�	KVy '��e�����y�̴S�|�g=�k0�8+��*-U2.mvN-X�y�K�H�E9P����)�r%�`�O�a���-�m���D��-���a�Ic&0�1�fx��Y���!�%�l޷������1�g�J
�w�����X��=�}a(� �DYpK�1��u����>��CLg�����t��D�2���&�������Bߣk�q��У �D`����昻�#irز�uʪ8n����vĲ���!��ŰJ̆����lw�	��IX�=�ėF�@H��A����iE����F]]Z�5�Q��⽇$�C�(n������f�N[��胧�$I�r��U Qœϥ�
 ^��@ڇ^)�!�] >���%?�𐪬%q���w�Q����8M�q_غ�6�ύ��2��ehCal˭����8�o�������|��<s�f�թc�˛���VP9�gq��2�Q�7�^MmkvH�Aԥ���C*���GP3=�UR����][
 ���dt��!5s���=�zi(�%d�$'���l����x)�R��,�p�?��?}�afi������V�"}(�Y`�.��u��
1������ (ضݞa���QR�4a�V���ܜ��F�XK#���$�Dk�d>�Ն�Kt�4�l-���x?�l'�O�9ݓj�M�p��#�"�{������c\nbq\5�3��X���1a4�a�SCn��e� ;�	�e�/3��]���Ńf�"0 �G`�kI��i�¬�*6�'S��6�Ux2��Ac�.�'���������M"$�kJ#GOz�r�l�����*�6(A%��� ����p/����S2*���cl�(F�t�V�@�F��i]�*����(t�>oq������ �*�k�L����T�6\Tی���|��� i:%�=̐����!xBu�o����2�ͧ��S��ۥ(���[3�t_�)
�.<���@�!h��'��dn̟���zɜ���R��[�CۢԜ��Q+=�����t�vƶ�@f袀QZ�@%��^��^c����*�Ef��ZY���n�+y:6a�����Iq;B��`3s�'�x����"�OH�
�p�k�1�XUlg��Af�����g�/�)�)�V��r�@&��ݤ-��&D�	^�6��Zs5���
��BV/����ɞN������l�CذS��|��nD9/��N�,�S�,���hE�c�)��#.i���0}�����47OOl����<ס�T����-m(�_��
��`�ikg��/8<^�����1�E5*{ U���y���Iā��Uy=�9�*
�����6Ἧ
��>"ـ饆*%���&J�vb�2S˗`(7�;���OH��q@����GE��@�z�G�ե�-���w䠿�^�����Z�/1F��]VR�DK�͉���ehpd,YK*�{�!�q�Ta��;����\�2���s�`t��!l������5�b��^.�=�w��i�8�y}�(�j���u�cZ��V������I[�{�yJg��7 �̃nZ�B@g&�p�n>�W��9�1�X������l7P���;d�b'(��O	1k��h�%+=(�%V�pN��Ee�L�ϿN�AXi�WZ�
@ ��ʢn"���N�@ʸ���u�(�oBXQ�Q���L ���y��H���<�S�m)t\��cj�đ%![��|E?G�-p$����{[mk _ݳ�3�C����z�/>A��)b�s�f��(���"�k�^$��b�-WU��3p��]�О�� �r��(�}C1����λ�0{�UQ���g���e���1gD����d��ih2�y�>w�?չM�&���N�j����E��������I�.��9��B�r��}A��� ��lx.="1�˵�ya�GEK}�q��=U�Eq+9xMH��>-BU�d|�D�ɺ�,���L��+�u�=��4���/'��S�x9�+c�Y&�kdz��Z�:PB��`;���0���8������a�5�)&-#~?Q-��Iڿ}E�W� )
\�%�еmwn%*��2�<G>9�RU�N߿D'"�t�_�ٌ�=|K�~��� F;4F�;�K<XFM&�B7�r7UСQ�n��#�i���W|�޿Z����5$/�L����LY_��'�Ŷ��t!'H(K�]�J]�UpV�Fr��nR�ƛ��3���F)�G�����n>U
�H����3�䛀�e�<lBW�]���ԭ���Y��B)M3�|K��A/��b�1���^)�3du�$W)��I>~;�r�T�͹�_r�2�{3�p1A&�B��·,>!�z��|{�V5�~PIC㪉��z⒰�Ub�d ieW���f;-�J��Y��{፥'����z��58��3O��D�b+�BVE%���Q��-��'B�Z�"7����p8�a@�g�UR���އNt��|�b�R�7`
,��Ư��[�Z�[�օt��>���bH�w]%�hl�\�{D�E]���b�7q��ŗeg;o��G�̆	�]��-�!���S�~|��'�u�zL��J��R}����C�<ĢE�}ĭ9�|��n�ׂ�*CR�xc���� f�*�t8��']�>+u�I2ҡ]���Hg�]��X�G57t�򪏁G��*Ɲ�.b�����Ú��{@X-�m�����|4���
=.

`��kn�&LF���ϊ:��t(�����������U)~$]�F[��QO0���Ź�r�U���el5=i�"�E���Tƴ�ǹ�cI'�:+8���W�[Ƨ_�z'_�Jj��F�xj"�^D-P�/aI�&,(�#��w�U�:�����	8�]`�9gw
�@�F}�5#���Bf�ZU]�`��CE,�"7��[c���Y��f?���B�HtUd�j6���-�%��D���B���ʲ����}y�����SP���p+{�b��W�vVy] � 	��M�5�&��Z������$l���6q��3qܖ�b�q�XX?s���0g����V
��[�U��Tx����)�ځhJ]�}�H�v��[)���䒽��@)�.Y�����Z����D
�\%��pͱ�Z���\�y`�y�F[*����Ƒ�T����A�&s�VU��w��O��(�̩�w�uT��|?��Q7�5г�+"�c�Օ孵5�_/%$���U��J
C��6�{2�ɱ��!6̻�-F�&u/k���:�y�6�B��L>I��R�hWk�,%'I����A鑠���=F���ʴ4Uo1��c�`J4#A.��:H��q���?F
_��׳>���q�l�+\�+���s#�0S��Vё7��F�j���xsh�q����i�TC�boF���|��[?rk0��i��F3����5B��S�w=��`�ܘ���"�oO�&�8�X��%�<%�ΖrQ�ׂ[�������nsN�'G�}�<l�x��<I3b�^),$� F9��`�̂�K}-�#�l�x(�r>��m�!3v&R�gIw��g��੓܈B���|����P�@�VZ\^%w�3!��t��'e[~�-�6�.Y��O7�T",��}�F?p,<�� �2M��/.\�8Z�� ����x̪ ��,���b�')�p��ό���/$���a�N���Q%����Fl�[�/Q��ǈ��!��	�CN��y*��G�������1x���K��Ԃ4B������>��� �X���;�c�)�Q�"Oh�,Lo��K{!k�9s�����k�[,���o��ᰪքcͫ)`[����L?\��
�QwEb~}��?]4�>�m�ϱ�6�KV���_ֵ���J|�F�3��`�`&N.F��i,�xm�e�:��h��
|K+�+Pk��)=zҢu�|c^E�\�YT��:�eѽ
��8k�������E��pB6X��oԶu`{��V�{*�o�����>L�ae3��ܧ{��y�,��2�c3T9��?6,��d��z�����XE�*��6��SN�ϐB�'����3�|�G#�^sy���i�!��¸Z�UhZH"�{@$n�r-�^�ǃ�$���t����Z<"e|��9�=��!�����p,=�b��o��������� Re�pE�p�Áf�2���J	�lo��YT�؄��1篚���C�Y"�	�rV�aЀ[�9�/�,������5^� ��X���8�M���ak��/Ȟ�ep�=���M��ݜ��5[�/�;q�8�6V��̍�����9 ݢ_{�����m�יX �����s��gVpـ-;3��$>��);G��NO�<u�OU[h��.�g��i�2����n{jA6^��U�=<5vl����Ȧ�+�H�c��z�P�>��	h�|�����W� �q5�οx���>��S(��6�{p��R"�rrv��������@�x�5��/l�J��7����K�i~���N�o�:�����jt�7��j�T\�^��
[.�OZ..��c��Џtq�HyBYd<q�Cv�03�T_pZ3�Z;���6%��O�z�6+nB�ʬ��)�����)�Q [e=K�T>���a�i�Z�d8G���+6��Y֕O�W�F���*bb��O�t�%���f��U�_��gO�H��V,P]k�Sd+����ĖdV�*�r�՞z���Af�w�)	���o�WM�b  ��b
�z���id��jj��h9���k�l�#Smt������وgq�L�hRL'�{*�����p�ωN-���t���������$�V)}��������6C������*	7��36�X���RF#'�1�?�
\�S�%�Z���K�n�Z[-i�F�>-�o���Q����>]�R�����=�&�R��+����<�ebX���K�Y�gI�O8��V<{f�m�����0|s�{sIF����P� k"&�ᩊF�dTW�ɯ�Z����99+�d��]4����A��9)w��lq�.Y!��{�E�]���0�kI�J��-U��f6l�aF�8����V���ε-��D"�}7crx�'�$x�?�����^49;�a3�X�5z�d\�=�d8�D.)3l]Cpڶ*v���fZ$�`�D���:1st����mF����B�2���,)\�������ujZ� ޷�F?NdK�}���X�v��s� 3l�쳃4�eL�q��]	��Xڊv��հc��� <��\]���!ߓ�$�28#a��!$�do- ,C��@��{��66��Ǥ���|˙Ӝ��.�\;��k�I�#6�'2/�p��I$�s|��:�X�ZL�E33_�Ǎ��i�5��s)rU5k~���!��(�]��fI �uږ�A�0��~���Kt-9U}Z���0�ǵ�h��J���ڰ±�v�ʠ�����]H[_T��$h��p]`��)b-��7옒z�Gc�)��!��_�
�K�v`f���b<MTRh��p���hu��XY���l[\Ǽ�/����Q�_��5%&�"���" �)���T]�N"��Ҹ��8�g����2���dU����y�oۍ����8Ĺ��^�Zni��;u�r+�.`d5GЄ��:�$	�2jp��B��z�����]��8zJǞ<O�"�(�8�
�{1�XC�2aDzA$W�?y��~��*��p��J�Ѥ�3h��ح/�֢g����F��]H�6�S~e`�����N��W��<fQp���g{ռL�)���_����J�p�X�)�"��Gű�3'��D���k�WE��{9m'BA*�� ��(���Ui`�Y�X��<W�u`�vߕ;fK�F�3Qɾ�>�ab�c��z �lլ�e��`�pd)��8Ȗ��b��>���f>�6k��z/���]�;�Fo��V(w�}>FN��P�%uL�V��W���'�_`�xA�D�4R�Ȉ?��`�z���x��45�k5t��g%-�PY9��H�4/�?h8����{�8���C�����e���n�k�C�^h�	 �TX=/�E�1�QS�k�:�ڔ���/;-��&Z�8A־ )}ß^_����>�F�.��U��4��'è�b��]�gJ�=|\  _��,���$y�=���kLe�P���o'�����4L(�f@NC�0�B�i#$�����lY54��!�+����B8�ᝁ܇��f[�R�R�BVqD�Cb� ��J 7:oc
���zM�e�ʘ�����&V��$���VE�mw������m��]��є�	~c\�P��?>��%�F����q��������/���{���q�r~t�u<�ŀU�\�J��U%\�P�VX��Etۂ斞p�Ԯ<�*w�#�YA�D�����1R�&��?|N�k'՗�56�`�3�,"4������%�z���e3d�(}Z��-����'�/%��2�eIX8��Ӗ����E6��!+��TwN����S�2\�qL�7���W��@��n���J����f�<���4�t׿I+����Q���I�����(b��d��C��F�Bq�K0�@�/B>�[��MKޡd�7z��
Q]X��j�zK�o!�uh۷���������ӝ��^�����s�g��@�L�(9�L���;����^/d�6l�75��.�a?�V��L�k6e@� �?����E2Q����ހ�/�&K"��!���gD؉/��(i��s���U���X��N��g,���3�3x�-��:V^��U�W�vqB�=<~��bV���|�'Ȱt��$V)�9* 8߭vPKP�ഏ�	ap��"��2�Yaψ�I��_|�E���QP9�w��G�,�����{����x���mWkil�Z2�P��⏳.���%�� j����~��	ㇶ_�o.~�d��=u�qn?Q��e�uŗ��٢�1���#�HϘ�l�����l�x?jM���7F��טa`d7���/���k凊�/���\���A#E%_��(V7�֎�}e��H���T���NK�Hݬy�4�w�p�.q��&!៞#�����{���C]�5c�w���m�9^ž o���V)2��䛤�Xc|���\MI�p��tj��5�ml�օ@i��.���G��K�� ��:G~��� �6W�Zx���n��`�O0�(?�Ioа������v*��;�ں�;l��qh1�- yX�<�7��4��b�j*�Q��^����z�<5�h����:�z$��<b<�����a@5�L�sܠ("p�����vs2B�WT�g���4D4�P�UY� K}��ւ�uu�%䉂�n��q\���&����md�i�M�����\����5� ��*��2����vtZkF���(X_�iÕ;���Tv���M�3�p���j� ���K��3$�J�$��.1!��kq��pgq ������G��gc,'#(a��=��'�F��S��|#�uo�Ք=��v�`z�;Qo�4��Xc�w��N;�-�k�u�J��yb�)w�����