��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0���p�?�gu:���@�6h�S��藑��92�C}���R�Xh�&,�U-H����QnU%~��^����t6;�V��	p�����<_hF�AT��o��@�Jz�U��%��Q �v^ĵ�M�@{����c�oNS�G)���Ml~gw6�209)�&0
���t��dE^9BUeQ4i#>M��Ċa��)�#Q���G�J��)M�	�d�"��HDP�� Gt��cD�?v4]r#ay�V��'�)\Ζ�z��W�E��K#*��O勷��B`mtoE>��V����[���~Wك���?�\���;����U+�c�%s��Nx���Q��>��6U0�	�t�㭢7�LV� �&(�V�J3}��2ʨ�s����!��%+��6ٓ���b�:��MdF��SU����7�`H���⵰���]�3�<zh �M6�ӆK�ؙ�<�T�Hx�9���[���,�����V0���d���眸�k(�_d/Q��)�
,)��y�����VIMu�2%?���n�<\�Z��&̥��S3;���R�D	t��B��+h3��`��'$���̴�&j2���(/��	%��{�I��T���R�S�;D[X��;�%>R���K�y�/Egm;G����p*�j�J��Q�2\���r�y �*��E"}X4�45W�F���|D��+����jt�+����p��q�S<�B�K43��;���Y���K��W��+=����W_�}�;'�E�-@�P�I�B�U���VI�-�vm�5��`���1�[��2Y��)�P-��6�	m=��]�#���9�O�f� H�����"�d�-L�.� v�*|�m?z��@�x��L���c-
�K�V�e,�;�J�y� Ϗ�*�Mt�����~�U Ȥl�Iܙ�1�zU�����~�dT��;�{|1&�y^�������6ߣD���v[�����Yh!���V�R{p���}.S��2�{^��j8�~�SΏ'����;$W� �����u�b7Xޛ5�K�ɿ���g�&��������}��w�E�_zy�#lof�6������~ǡӁ�^��\m�W}�l`�?H�M�|jOA(F��v��?z
|� ޡ>ҡL�
yng]�ن���R�ZD��	�n+ 0Q^�WRVq�$��L�2��ލ���0%s����)>k��}X��j�G�Cu�k�Z1y����\4�21���v��vL��f
���,ʀ��=b@�!�������E�����M�����+nKC�Q,�N
��a��5�`��//����t��<;N5����`��<��6��?2:4��H��Q��9<.�%��k����r~���_���9�$0�=�`��3X�i���ct&(�/.���A��h[�z;��#Aq �xL�T\1�f�A����v�5l�H�S�>w�Ջ\�<p@L�C�:�1��v������(�]).AV��r�PY��x.��yi�$>p���0��2 �Ӹb��W���g�Ϛ��/�lp_�֓�Rŀٽ`�=r�DB�n�j�e���g���%#�^7|W�躐-���$G�����s��J�w�F��e�����Uڸ�-�J��,V�*)-�w6��!9�]F!Q�{$�ѓK��Ȕ�8��`�K� *-�X~ǟ����$��+�ڧ]N�2oȎ���:���p+������y��{�
F�Кq{2��j{�v�I�S�'Z9\�=�T��M���j�Mh���g^
_x֋FآV�Č���Y���M��,G�f��R?^����͛эL�@�'��ÝUE�ŭd�U�&j镌� �<#(��MA��B�զ%�X�#|�ORj��,��b5��z_́t�@D��qG�l@�ب1��Dd��Q�>��q�""��U	���M��Q)�&w��g�����.�h�����M��s;���_+���� ��L �̷^��~a��7�ꣃK�ܪr�L��5���#8�T&���tE�T�B-�3��q�c���\J����A4!9Y�S>���FJN��s��yR~���p̾P��[�p\[3z�B�X�\����"������K�HT�a50��x�8��@E�����3�ۈP�����F��K��� ���=#7�(�\�@�>�uV��)�=����@���Ě^+��l�ƴe������R�r�A�-Eg(�=L1o$CAa0�zt_k���Iǫ7�����4z�H�Y�h�D�bm���Z�*�ؼD�@t�FD�TgAg��,RB�t�q�%����t-5��7�7���Fc�����}� ��8����1���{B|Kβ{�C�V���|	}JH��S������:�2� R|��u�2r�꟡ZW.���F���Z�#�u�wM���+8�]����K���ϧG��ů��b�m����~3����Y|���jlI ���	�f�~=���%n�ef�����w_�M��<^a�M޷�Ap�V��Z����<�j0 �W#���8Űb�����p2LyN�5����<a��df�-�^�9dy�P�b�ӟ�2�
��ZX#q���B�Cf{��oW*+C@��՜=~L+��������v �6�a���[y�\O�4�=�=�]����K,-�o��
.���v����9f>;椥ҩ!l���O�}�]F�E��j��8���Z���r��Ν
񁉏�=* �k����rA9���!K��R<?�]Z ~g�k�WH�r�
X�ą)C��:o֙=����C���#��8��US1)%7���χd�^W ��LK
1�W�a���d/s�K��󝔙I��3u������';�����R��w3�6�t�N�	����:�N#}�dU� ��b��ܬ�M����M��V߬�����ڣ>�5��a�:t�D#�N�G�_��t�NZ�H�!7I�
�n'�(�\	����
t��C�-��!�xt7?�b�T�W �]���h:;<��f�z8[���잿O	�rK��ݗ;$������uh�=�L.fFj`.�Y��"�[�����	��V�� ϣ8٨}�"�UK,���ms�J{. .lUN,MZ2)��[�hu�\��Ξpzf!^�jB���W�X���U������x��4�Yg)sH�(7�AeP.�Կ�*܈`;�������1]�^3�Vv���א�p�hj4�w�c0�P���<5s�wXH�w?�Ys����!|4w0�����u�A���i��?��(��lfٵ�r�8Ʈd]w��͡}��2�u���n��̨��U���̀�z�:q^��d��?�����y¨g���H�*����0�"r�v�Dr�k�F`BR�G��/��.���G3��j�\��I�9t���J ��y�(�+�ݩ�z��C?�Á�Fd��=S�w�yQ�G*�j��� p��,��	�M��*8�)�).ʃ�F�˅� ֢	H�`�?�̚�ӟᏧ�?��Q�ӓ�p�F��h��$ղ�9!��5n�gkX~�^���~�xY�s�kQSZCkXm��T���Q>ZhJf�曱�y_�Z�O����A��#����%��s�ϋ|e��5�sL���t�4(Aؐ�{u�C��X{I�R��0oPuK����d�����#�^`�;8������wWu���KO�A��'P蔖J�+�Ǐ15s�Ė�X���G�)�"m3X��u?��N���~v�mv�;�jҮ�cEY<���&���~�Q7�7!�hߩB^7��qb��-V�)�� ��~n���p�ZW�����S�����6��re7��S���P��(0����R)0���]����88���:f�B3��sn�>�x���fL�[j��(p�*�p$��&x7�uU¨�AF���5�X�t�'��Ұ��� OGy{�#-&�Z���_���T�4�����������l�w�V�kd$�>�0w̓�eQ��x��'^A�7���N��.l:N�T�LU?=F7 PT&�U�n���������E6��qB�;l�5�د؈���@����f�\�_D��)Ђ��}��䉇d@�WM�O"�-�Ʀ}�C��-[�Dg�u�:���/䱎k��Z��B��b��6�EA�N��=Î%1�(��Z�"\����(���I��3�H���晷b�HB�wq� �xw4���Mec��SgD�9\���h��	'
Q��5K�"ܨ��Ho ������/yb*~
��K �J-��]��W�B�"�k�\F}��ppC�
O�7\����^Z�-'µX)W�5�3�,q��O�f����H��;�6���Dp%�S���n6l�V��à����=,� ���1Cbǭq��(�\`����g��ia��p`�|�N�L�p|RNۿ�8ͮؑOh��Lo#u[�_rbiF��hW��P���i8<Q-BB:]����ҞH�����{��K���IԽ)g������r��}^،��׼Ξ�P6EWFø�G:�-[�G?p<�.�����7?Ln/Þ� ��}D۸-��Ѯ�F	j���H�j���+t�D��Չ-#"h1�D��ǵ�6+�׃"L��D둤H&����/�	!��G�j��Hi�9�9H�(���0���V��Xu���U�2��ٮ�����Q�F���a�rɯ�׫��P�P�7��\DF*�Qִ�R^�u�槳�����Wd�=R�a�цT���r��͚�~#>Ҹ���@Y����?.�N�~��8�W�؏�#s�ȝ��5��H�;)
��ۍ�n�F�_��.����&M��a8Yj�^q_��Њ��j��d�S�P��$�v��p�R.b���$�����&N��U��6�G�B�g����2�@qɾ��}�6�MR�<�a+����3$����w�,m͆�H��B�g|s[����%��J��t?����U���D�̪�S��G�/�4�����3�������sj��*K���/��i�&�����q�.Wͪ7��=�܂O+UY�/��>�ߺ������Z=@��PH��;����/Ѱl��jVe��F�N��STL��H�(�:�D?�-��~ig�mt�6��	�9H���j���$��a;��y�@��8�l�"=c�ε�[qж�O�֕�K��P!Rk��ȐߛrǺ�F�fWp��A��6-�_K�u��v;\���ڹ��jOQD(�Ԧ"3X�0��0
P
9�w��ȗ�$#}�n���r���6?e},1��+ӎ����{�(���)��M�K�_}�����9=9~:9]�a^~�����ȣN�yQX�=����6�D���L�p�=S꾟!��n�<����! �a��-�aQ,�S�TP:�Y|� X�9k��h�ד�+X��1rO/��@qN��IBb�_�(պBy��}�|����s<	����U;�@w�dYU��R��o�:a>�f���ă۬o� ��{ޕ[<L~}b�e`f��%M@Z�t��`�`н�$0\ן���^$u��'6rxd-A����M���`�z�]ǦWQ��h�^Y�GI4m�������1�r={���?db��_�cq�E��K!�[�-2=�B��@|]@�o`Y�VD^+��~�b�U����(Jי�q�"�����l]�V��`� �cq�s^�oнoE�R�X��:��:�V���s�{��?)����
�EIF���a=rm���M����T@Q��*)��d�V �&��Zg�D|ލ�N�/�X����׭����Z!wYD�ykR[�����s�0�{�Αo@̃hw�5����Gن�e)�S\���v��`DZ<�$��$���k_8���O~F\�:	�����|a$��y�����4!���/�C N�㣋4�3ߠ�X�9.�}NS#��Y�,�-BS��I<�kj�U��*�Y�������5�g�B�a��Yޮ��yY�x#���#&ٮ�������p�1pDpҜq��ˡ�a_�����Z��2ڠ���o�6�ֵj��M���DL7S���L��U�+Y�j�ᦪ଍�'�:I{�GF�).��V�ɳz�<�9�3SoP�'�.h����jp�!O3����ʽ>�/SgGX��l� YEf��C4��B�>\l�&�QD7OQ	D1t=�ݘ�����_\��X
.Y�Q܋Uƙ,Z���w�����
Ԏ��߁�=\�Uŉn,8k��ZPz� ��Ꜥ�#p^�����x�+a<�&�x,�h�Ȯ�^��ݹ��f��^��J*�Ef��y���S^�����U����Q4�/j����x�튾�4��8�A���������t�IX=���ۄ��Ӽ�2�SE�aB�ڏ�;+E�N�ϸ��n�s�X]N����@L�E�a���e���Wװ�6+�DHa}zb��D���:}Zz}�Co�'9�2ٞ�f�Qb.�
�*D2��w�5�jٕ�~~��ť�GI ��xJ�%���j�*4�5ǋ�Z�߫���{�����2���s�e��3�#\����ϊc�'g��$���>U?>����$�1_A',�d%�a��A0�p�kOF�k��:� �^�b���7�>�� a��u�`�����`�@�٫m�l�d�����!�����=(dYe��y��s�ZÆ����W_BF߼Fl�x0�際�~E�ԛ�A���s#����Rvςㅓ�M�/%��y'k<"���0�����b+wp �J��������}�!�]��a�T�#�W(��=']�`7���J�w��zcs`�����m_�����1`Z6�V�=��Tѯ%�P�o��;�$�4����+�"�S��8�ml��/��m�i�h�����%^FW:
���c0�q��n��-�	W��*�����|1V`���]�
���|�0�n���9ٝ)���d�ӗ��vGp0����:�9�h�o����Z������&U���xd��mQ��v0�+<�Kr��7f��6%���kW�6� ���Lͷ��G飡�_�2:rH��w�QhT��e��95\��ȑ� �kJ�1|�s�ݿ9�&��u�P��轚�wCT]�Mjr�3{D�(�mL���4���8"IM���ɾ���D���d"d�-�=-Ixm��USY�(!��/�0����ֱ���[k��߭M�:�2��ϑ��7�0���ؓz`�f5�Y���k&��B;��*��^\���e�K���?�YM��a2���0x���N!��"q���D�?��l�S ���S�0_I��!������mj�,��F��Z*	ӝ���˹��ÕC��ƍd��B�ǧ�#��]�M�k����Ӿ�9SB�y���9�V�����: Ӽ9�m��x�1����B�][�-�d�`0�u�f3�< �u�4B�G����i��i��D�	� ��k���Y�y�\_$m:�@�!�]��g-�$+�3MuhДr���/�\v��73�Y(;%7��zg����ƪc?}�'O����-��#7��]#:kX�p���h�ȕ�!�&� E�-~n,�(��R|�C�L=`W��Jj��&�UE�B����s�*�4��/2zwÁ��� �ZkK��6�{�����p��W�Lo�Z���_�5kۃc�%N^M�ݽ{A6�TQJ��ύ��wȖ
�.^���wtҪ!1�i��e
�q唺Dx��0�a�ش�*/dTݦf?i0�7���t;Es�Yj��C1��	(8D�L�%����u$�0���C<V���D&;������1u��8R�r/�mQ�P�Ɗ�R3d=�p�W��֦7��;Q՟<�̭�%IJ�m),W�Y��IA��7/��RM��c�8ۅx���ͨjeY���G����N>$ru�o)�(S��ZH) (�ϣ��׿� ��đ��·�A�5�tV*f
� �`���V���>Dy����H����4B�>38:B�S6�/�����z�����d�=�dNi���9���$�O6�9O�]������#�8�T	�t���>k��B�d��;J,���Q]F� �)�^�Jꡢ���^�J.s�v��MP�vp�8�©�	��I�A�?�:v{�H��=L�2���̋R����t]�!�/`S�P�LB,�Ln�;a�<`���tT�#\�l��}�}��%�?��8i_�N��׶�&< ��<$u�V�A�}@���D_��5FZ{Tu)��e�"`���F��OoV�Z�i�0�Z)���Ȋ.�2<��0n���N��N���!�gHq�k������F���6JO��5Y���t��q��,��r��\�G���C�t�1Z��7�'���gK��>�؁Sq `��Jx���A7T�f�m�Q��hO�.q�"�_�"k�p�	��:�&�l��{��=%^�1���9�<�bO*D`B�/eEcQ��
��6��[���eI]��	]V����S��):�Ap�F���e�/B��N���������V�R����d�z�{r���|%�&NR���Cޑ(�� �f��ԙ����}�N�&M7�[反hՊ�|����vq�TĲd�ze�b؛�1:��z�iW�/��#�/S���X@;y`W�u��JI* �4��p^x�ˤ��	�����z�YH�x�H�{D�^D�����Ȩ-OVR°��RE�5���h����>�̢��.ᜬ��z�\,�֍1V�?�HH��b�ښ����	�Q/�&�ʝPl.nmU~�M�^&���𽸧���6��r��Oz��N�(=��˪>��`:�I����.��t��0K��Muh[�s:]��|�QAI`�Zs둊�.����d{�7�V����sN�݊�d�,�!������Ho0����f16xl�[C�z�R�����	]%�68J
͘������4=�0B�[x�^�͢L�E�\t���>���������p�x./�������{�{PV�}j���}� ��ћ7����|
�����=Г�w�{�/�? ���%LgE�����|�o�q_��@�/�]����d��_. ��)v��4��I�$1�T��� ��p���p�Ǣ6ƍ����.
��X�n�羡����!�ϣdD�2�i6D؏��ħ�� �u6��j�q~ͧT��i��~�l���̮�;�#�dVTH��x�G�����. @�cBBLo������V$d���TA5����F�Wgz��o��z��Qφ=
m�,��k�OH��F;�V[v^j���'��0�(z���(=C?��7E���-�p���1rhxޭ|�5	�5����A�V�#�yd�\��I�wZ����>s^w:Ha���s�&(�tZ��*	e�b\-��3ё%���z7�Q4HfoX��?׵�}��(R��	�U�(a�t���+����rV���c��T���G��!�]ƞ6Ԩ3�h4���::0Ɔ���� _��m�i?`l+��[���(�Bm�y�Ә�r�� �R�+2{DU[։�m�a(�v�dY�*���a��.�u�C�g��-'y�Z��w�B����,đJ��3�[�$�5YL��kN�U�QK�X�����S@`:��ۨ�&Ӣ��l�$��w._�pO���m�����ʏ�T?"�'���7�(H(08m�fcW���8�h�i��<��	��3JKx�E�?��R	-<ε.��>�-����D-x�?��m��2?�\�w�)4� ��<YN��Q�қ�q:�@�p�p� ��.�����P���f%
g�j]*.5
o�����gK�H����\��n��@��R�`��X�=��m��^[ؙkw� �����E[v	�#�#$.�\�w�l��}��VdJ<�䳴{�Ũ�bm&�5�i�$9��l���:�[�z�3�tK�)��u�H��d��YfŶؿ~	R���x}ho�����l�����h�]}�-*�WQ�f70�<ZQݠ���z��.��\���6'e��=�
ډ�e�>.��PTqH�����i�$�����_�狒L_9��<4Y�Y���ʜP��A����q��<����}��PH`��g�����H�Q�zt= d��c�����M��XU�)��I9�⎑���>z���������$
�`��im �l��R�JV	U$�;�j�al=��u<|�2��L9���U�_�җ��^���8Rd�.(֓��\���n���^�M|>L�^��H��.��Ɣ�����9���`U�H�Lgl�v��z�=:�k�E�B�`�&*Π�`�,x�/Z�_�MX�@!e�Ȣ�$�q��.�P����-z�l�Z�2IE��2!�����p�8P��fƨ�iQ�;6��(��D�]5ai?�W���i�<ʪ������o�w��	�����o��*��y����ȱ���pM��uF���b$V��\�eʔC�4"��#0�R�J��*��=�.?x5��%�� H����p�=7��`$!,�$��k�A&*�:Xj�Wڹ�Asz�\}��n����E�L���.������g0pB���>xR�(ܛy��=Ѥ��e��H�%��,,uI�+�be˻/�*�|в><�X���i{��ܕ)���m���PI��h�Q�(\����#���37dup��n���զG좵G,��H����"�6�^nΆ]1=tTr��[s*h6^����Rn�4y�O��f��)��c�;+	�d�Oǉ$��Y[��\?&�Q�Ly�H=t�'=���H��+��ї�u!�,�r��S"��+�J||"����*Vq�ҦW.�5 1��SJ�%�0�J�ZU�%����K���]XW���c>톄�:��S_.dtst���� :�]U����(49�2,��s�a�F� �բ��P�p��2�F�<�ݣ�|����k�C���9���1H.�'��w��!�Z�t*�%��u7J���AS��Ֆ@���ݹefp^���x��Gb�Pߤ�V�������jF�9o�J�Y"Լ��rTJ�l)9�/h�����C�Q�� �YOJ�^o��
�I.z�m��w~�VRB9����dХ;|\�7Q�,�@���	�]d�G��[���K ��uZg\�j��n��6<���:Z��On %M���C��j�N����f?f�hkԶ����7�zĢ��z[D
R��݁�sk;�Rm{R�� ����#R��0�ǔ�A�������]n^˱bЯH�����"���J��ڕ����}$CQt��� �^�6�+N7b���VI,0�/w۾��qW��H������`^�U�4������p��o��S`=�"F�Ȩ�տL��&7��Pk]˓n�6������W$tC�?�����kTe�$��>`�����E�[�u�Č;D����i�ʏ�Q���+"W�����Z�hڰsl	�R�[q�sU��E��G�c�,S�Y�a�8ߣ˟N��UlLgh�꾊���Ge+�� ���9l<�ȁjs߻k�|'Ũ�(�	���P�4���j����?�����a�����2���Q�/�Rx��%B62[Y�����|l�2�sP���E��oVt�&䞍	D[k	�oC ɯOO��f���tҽ��m /g�NQ*U�L�6�M�1jW�e�����pu��s�FG/�M�+��� ���ܼ�|����(/|b�������y:����;���qTP}��ĝ�A��S6�f2�vӐ���H)ІV�QMO�-*��	6}ͰP�z�Nd�UE '	=/��ۧ{�V��%�����.D�QO�>حj�'cc_)E8�"6�g�>C�T�1�	v�D������9��c�i���F���N�\����xT���qT�eF����6�(<W \T`͗�*�v4�Gy�I����`�W�3Y��� 9N^����`;�{z+�'鷵��Y���=��ͭ���Iw]�e�	^�h$;�?4э���+�8�����u��1���޲r}��4�|�%�J.?��|�% K��οd�7����<��W��?�<t߮}T��R	��I�pЦ��`��C�����	�"_�C%P�{tE���M+B8Gut����A��`]�[���V��[J�ܒ�=��NS��-$< ��۟ȲJ��#5l�i���p)�-�,pz��Y����EA,<`ZK
27�F�,�;%� �]�6�_���HKG`u��a�8�U7�$�RS����S�w;����w������dc��˝�)D`���Ű��Q�;�x����j�����awu��Jr+��� �!Wn���1 ��z�"#���ҢU�_6e��蠦� $<�f���LE ��_�a���X�8"��&�����u6y�k9�y��aV����U�*@+D&+�ljv}�5o� �&�b
F��k���6���GN��?+�|���xg�㰢s�'������p{&IB=m½���r���ڸ�@��p�R�~�mc�����jPnm�Y�49|��m���XY_~�]�A�{��jNI�1���.����Ɉ��i� �M|�qM��wa9
;vU�s���8#�14)x�$W6���b{g�F�N= ���/�N�{���r�����������-��)������X	Z��Fb,��~�9;�*��|^��iOD��$�ph#��xw ��쎝vP|.��a �)���uH�qda�[�稻j8o��n>��;�.�h�@�QY+m�N��v�O'��gFe�C5�9�eTG��[d,�x�U�/�icd\0WF$n�I�ޱ �¤Y��t^��޿�2;�@Sx��[rG����󵃠`������K�eR�Ϳ�hZ��+<�Ճi�<���6��_���K}���X�(�=��yC��>�]?�0���r�FW�P
����jч員��0b�Q�V�	�؇tY�~^.~ov�3f�S �����	��h)Ɯ����b̑��QZi�3Zz����Ds/����`r���}^ZC��᪸��x���x�,DJ.�[t�i��b��|xx�
����עR�=y�z��Y���|�2��p�i�p�3��U�L���� ���v|~��@���O�6ѱ�`δ����6�(�9P.�Q룰;�~i����qO�O��
���ܜ��F����|ዏ�^l#-��m�6Ȅ%��g��~*�EV,/�8P!�r��0��E6W�u'�����?�\�lwB�w&�t����s :Ȓ.���YZ���n)�#͛�E�_	�G �$N�v=)A�#s��eb�l�k���^��Y��3���q���|����Ʊ�g4=B��Q�p�\�Ɩ�~��ȅW&�PA�B��&�iaI�Vj�G:����˪3��ʠ���Nx��H{U{��@�MB�E��Dl��۞g�[V��\��~�:		���z.�7������Dmz�l5���M�ۗ���|�<�ɝ��%�Y���v%��_	�űYɆ��O\W�+���Wg����ށ���7j�	��$��+�ݯ��ڗ�!y<������)�Ǻ��w���@bQ�5K�nQ��E��R?��@�r�"�h�Mʐ��Z�R���Z�-�,���yWv����Nm�it;�<ĀQuf�lnӃ���.�Dv�Eu��������m=X�����P���]
�eў{lͧQ��{�=�W0��B�'�W�s�s߽+By���X%?��m��O�;�F�S찴�����l��8����*�,C���y_�%�Ei�i*z���z��g�;��E���+`5�Eݴin���=��D��r4d)�R���n/�ZҼG!��7�l���������v`8���)���L��N#e� ��ұq�5z��v��v9ݧc	b_�GRo�F��h����*/�
��~��!�9ˇ�e��@�Cy����L��5�����3��j�����"���`R5�-�B@�0/�� >@�¡�%�ֵm��J������� +�c+�����4z����l�
cKxiWo܏��I��1�W��"<�9����wQx��Ԇ�ן���|�����d���u�w�k�.3v{�u�e��	����cТz�<���/qX:�d)�k{`��N������`����)7��n/5k�U4����E^���.O�	.lP�R\4
<\_/�9����dԿ���Ym�Ų1.�� <����o����Q�\C��S>4v���.����	W N�������,mL�8��gt�����g�=�Wyl8,T<�sƥ6��9fXq�UX�
�~�+����r���f���?���sYPn5����ĩ�'��C&~_͸�+e/�G�����k����0�}��
��;�e�{��$=f�#�"�*AfP�|
8B�gC.���E2��QhIK����'}I�z�<��@FX.I�j����#/�/���b9������0~j�Χ�@0��*�wh���]���SU빤��{����K�e�xWa�Ev��\C,T��1P�iT~���1�D�w
Zո.w��>nO	z��0	�7!�����Ǧ����:� �[,�_g�'��p���%�D��Q��1�J| �j0㓨fd�H$���#��K�f<Pɰ��Sߴh��+O�q���<�;,����1폝�d�}r�6��[NفGhZ�R/\�k�!�]�:҂nS|�xvx8��G&OhKh�l���侳Ȳ��wLZG��
���q���>�oc��6��rG��,���
9�9|+�z�&���I��>�\�}�}z��g�"�PD����!ґ�㢽�e+�y�:U�}!���--;����τ�G��Ŝ����J�?7m�}�d�n��>��&��AE�|%��5������qQh_�����,��n��'���gɰn������țn�\��7T-	��O�P�؜����tn�/��r����e��eͅ��o�KK�ދ0X�F�i~�b��N$����?5�B��M��1&�1'�lW���}���L9�Lr�vy��w�)��1`}���&�Ll(���g�.>;ۀ��ӂ�E�Q�B��=H�;�Y�bDE��]Dv��4w�����Qڈ0�Ȯg��Ͻũ޾��������1���N��W$C�$̗|��QLa !)�V
�=g�2��V���QH��L�:_X���"������3딩�ib���]�ؗ�C8�R�m�M�x�P�/p��v�����=n��Nٻ�@!F�&�(���dQbG������ύV�5I��҇���'�9,��j���{�UK�|���|���
F��PR��[��!Zrh9��vfDȍ�#ď�����j�"��$jA@pL�W��d��O �*D�Qhx;Nr���&�	z��֛�i���{�vQ��Z��?e�j���l.�n�K,��dg�$TyY���*q ]ޜ?،�O3�?-}h�\)�}4e��~�9ƹF��n6��<�,��g<�"�6;����V8���ys8kr���OF���y@�����0��m��}�P��k����.uR����O�bյy���tZ⁸�.�[� ��`�!R��������x��\�qZ����C�������*en܃�������8�:���F�S�����#}<����=́4m+�|�|��@:s@ۢ��ϗnYo�#so���9��J�[",�|
0H�Bğ?r	�ҼƔ=(�Q�P��M���"�`��)ބ�p$�{\��뾑q����WZ���I�G��|���^��9s._s��t���� ����8m[/yE�8VΥTe�`4�J�$ߨXlp�
8��IM�o��A5d���>CQO��lW�5à�wl�"N��K�ȹ��ZM�z���p#��]3�T���Eh�*y�'��o�Y��d�`?�׍���p�l#�@;#��4Ӂ~�n����k� �ｕ<o�U�4�f�'">�R�_��ê���~�\x�v ���>�r/j�3)#�۾v\�~Ьv�G<�bX�����g�AvmQ����:	�7q��]l�ak�S�U hnv������q�?T���$g�����N~u�e ���ބ^�:���-iG���+ �d'(.`�n�6�1�AA��C���M󠩱��ӛ��Vv�@1�+�r�4Un���J����/a��u���K|8"�E�x�5���dA�YZг�J5����铈�AX:KB�q9��O�;�J*,;����IJ�)�}�+u�����GB��o��7:�k�.�c9v4�w=+T�����J����WP%]�<���}��N��T�a���Lp9ϊw=mfr�L�6p�=�Zڠ�� G�,�{������PF2�#Z�����>�g<y<i��,��V<����Ԛe�����9�p�k'�&.sI��:�h:�*m:�d��5W�5�zRɥ��o2��R�v|�b�z���,�jy��ӗ��̟�M�e�ݕm���?���|���`�9
�j7���� �J]ĪE�s42%�R)�����ڻhLBj������nՁ��{h˸� ���I+ۼv��5������>@�"dy����(B�x6��~�M��]�"��{qX��Ns�j�#��ߡ"L���ڿn�MK,_0E;!�X��Q,+��
l�L ��m/l�QX
��~��9����'�cu�ͯ�$
�"���R���Os�jڤĢڪ�ŷ�`���c���I]����׋��%v4J��ex�/����
�XI�:�K�`Ĺv�)�R!E��W]l��=�d�X���T|e��}ǋԳ(`������ғU�nu��'7�4Bw�D��B�6�=Y��ݿr+��em���*	?2'��'p��wPv��-_8�r�H�Nc^E�-�іo��Xp�������y�D�_h���'�;��V+	=�7ȓt�ӣ�F������|�n�ޜ1e��	�3U�W��Q�Ბ�n�[ͻ�'d`.�-َ{e΢�-����_�e��`Ih�pH�$�y���P��׋%;�)��n �L#]IN`��w����g����a�%CdZky~x�n�S_׉�ӌ׿��?��DSFJ1U�J�
��-_�?����1��}#6
;C�P�#[7f/U���}_*kG�VY���k�4l,�ų�MN���\�W^��LP?�si$�X��|�?�S�hMc�s�<�����k|ː4Eu#`�.�����Jdhh𧾣�i�,5�P��Q�%��j�I�b��E��;�����+=�V`�w���Ňx���t96Ä�ӧ����&��C���r���H�Yq��� �V��w��%�"�^�z�k="M.���<۰�\ZA)�z/z��=�j�Ha�xP���%����Oz-g�Ֆe ����i�>�ԍ&�������$���zV�#p�����̓�zU�X�KMj�1IU�:+d�B�Ur��rܜ��/˹� �h��ܼ����@�no-3��L�8xz�l�+��w��[:���HR!A���u�-��o��e����uU49g���Jw+��:Ws.��KK���2�_�����(�n�h�^����Mw)�������������o�����r�}�m���.m�w����/!�(�:���]lo��9��/X��UڄEt/5-8M�oD���'�+���ׇ�6�L{c���2�D�>-ǌ�=k;]��z��#��y���!P���Mvԏ�l{�?��Nu?7	wO�c���C�/r#aO�km4�$59�^1��|Lh��ϧ]pO99�[�c2�7R�n12[�K,1��K�g®T+Z@|��J^�S`����@x�}�d���o��-�����U@�MKN��C��|�r��L=۪-��L�kJ�%���&����Ћ�;��ÄsG�"��f�{݈���`�j�����ǳ�����E���x�p�����`~�ςn�\}CAc`>,���Q�*�5�<�v֠O��v�}0���}��%(ԥ@�4Z�Ev�i���9d"���7Q��3�Y�/0+��Ɲ">+�rQ�'�y���Lߘx �3�5�0�%'T�!s�V �� �DL E��Y����<ٓƬ�PB�c$`�53RO��Iy���� 쌻d7menq�2�Ѐ����d�^-Q�������5��:��8��,cՕ��4y�勗�S���ʴ5jhK��w�b�i���y"T/F����Q64�t�����C4���KEg�e��_�� ��>+ ��ҹ;��Jw���c��SX�9�Br�T�ss��gٓ������kFC�s�XG��f�'������q�X�����2c:S�x��X
�FM��#��84'��.^ʙQ5�>w�k�������B��j������cg�:d��yh-&m6n�͵` ���ݽ��z&��}�+�m��c�/\Al#VT_,5����xt~�5ž��j�=����[.d����I��U��G�/&j�C���G$�lٖ�MW�ӝC�hC�Zv'ovb�p,��ީ!ý�/G�ykaQ�.�k�?� Hd�y���X�]�Pݧ��mn>���5�z�͗�og�����s
<7br֤1��˩�'�E�gt�|WWHr7f9�I�֊�[�o]�����F?��x�d�:���n���a,:=G�N�C����_�`_⼓�J�/��h>iT���jN2+	��n4��R�
�+��}$���.�Ƶ1���L쬓19�:��.n8'\����D�c/Χؔ��WRc$R
��2|l �=I��&��H���pO�I�X ��-(\S�gB	fxm;\�>9ae��f-�d�҂��i}���P*wf�ȻN���w��U����2-g˜����U�6@[�XDV��ݯV�|[b��?\�Y�4�#�O}���uS��0_S�����]P*��]�}~��	���#�de��gs-�6͇��A~1w,�Dp��1�+S�����"XYˎFL�o�J5+��BH����aJ��7*�إR&w���>��ڍ���mt1Y�aG��.�n��qhi��Q2 �k"��%.U7rv��$��!���L�^�T� -gH��"�)p6'FY�3�zh��LVu�+�pn��u9�7�k~)wA=ț�V�A}�����^�Pt���*8���u�J��m�Yw�n$ ��`^7�"H�G�G�5���������DE\)^bG@��"�2PR��*s�z$Z"��A��n��!�*/E�g#����++��6�hOy�l�`��ߡ�Z.������5�@�z����7|�>xaH��i@��l���Z���w�G��/�-x佀&�G,�iB9�*E���y���$�4����J]R%sj6hd�]C������.u���0�=���^Tn�W��D�0�Z����G�����q^�>��p�f��'؀��*B0*��s-��76݇����}�uTr������I�T=5}ʔA*g�����OՌ)S�o�4�� ��ܱ��ɩ�(�Ij���2����W�"�Q����I���?�Sk�����E�X��8N�)�; ӮM���U�H����6��f^�[�K�x�Kh�x�*���6�MT�:�G��aC��sgm���7�0����Y.L��BZ?�$��5l���&�������mS\�V�l�y@��1K�nFʡ����|��?2ڐbw2�.��.祉dͿ态bcB
�#��1lo�&�*����6����xQ̥"D�+����� �nQ~�>2#�n,�f�7��a<�`-������M���fN��D�����s�9��	�j��R��w�w���W���].4�������h���*��R$��A9��Z�~|I�<0S��vA�iDA�g�o�|����\U�*Pj/st���G��}�p�:�2p:�k��;�sn�]��0�p�.Z,��f�����:~�R�s�a�do5pa�~<�8�o{�~0�m�v�H�A�Uv�����k���^<�~V�B���5FU���Xx,oR�Nk	��F)����U��)��
�T�F?�r�����M��\4r��3�G�KG���z6A!�6�E��gSBh��ьϮ�6#I�AN��k���;>������h��
d��}�̲����҂�ZV=�)ڑ�_I���6oS��~�$�i�s�@���LPgL����C�?��"��DV�!�땉#�4#)	3i� ��V�<���)\E��ϗZ�)ܙǣ|��u.A}d@��e˪s�Nsm9t�u�n" �I�����7T�R��7� l�k�i#{4��+�F�9��ҫ3����U &����'V�p�����4P�[��s̭}a�,�զ����A��y���S�˪~g{dI�g楒)�@U���0Q4��0W�����ǣK��7G�K� �������5J���i���oSm��B��,�=n_�N���<�+F�F��e��ES��l���}�k�%��;p���4�N�Q�BE`S?O�G�)��Wq`v^�k;>�ٳ4�9}�[��z�Tdcp�ǰ�w�Ud(��v��R#��@C�|IG7
3�1(|8�m7�&yw�}�WBz)Ǹ�jb�Hh���os��T-�=�rD��@|�=ti����q��Df���c��܎�����r�A'j5�HDu,�A*b����eίj�"	S.�&��,� m��h��s��]e��~������*8��Z��K�գӤb B��F^� '�a���9B�o��и	�� [ef����\�i�����`be�)�����@�Is��, Am4T^�p�o��0�JѼ����?��R2w��-�W,�&k�X�����f���uß	{�j=U��;;mgC*���̊�KO����;A����V�*2��:֕�w�d�W�$JM����'�z����!<�>�0\a�o��p\��d�Ԡ_������{�i��Aѡ[���c�T��g?e�����'Uتc(`�_�a��M2�5�l�rN��<6��q�>	5
1%;� Pt�� |�)[����9+O�G m��|����
)J_�{X����U�'P:�.��z�[j߯W�+�Ú=����:K���N���?��#O�V��tL�n����:Q��_^��[���B�����n��=��IP�73��	ۇ[��)�}�L)A !CZelW��į�y@�7� �Hv �z��T����.����cp�,iQ~��+�W���X��A�q]�;�	�ʕ�0�1�`P���hclj�!e�R�����,���/�����(7`�����O*�u�c�K��-��h�{M�H��g�����i�\"�^�)1ed�s�p���'>�B�Z.�훢)�z�.Į��#pJs�7��
, A���]k��ٗ׺aB�OQW�X��$tg{5�9Fb��|F(�����i��5���;!"�U̕9jL1C�(k����W����/=5���~���'��z����z/���p�jX����]P��?'x�갪2��¦4��_Ѯz4���<�����:��Z�k!j��W��{�������P�s���abRĈu�I�9�dTڌs旫��<&DeE	y+����=��3t�}�:�m!iQa�?�\\X��������r:g+Gy�z^p1c��*C~]�Q�%%w��:KM�b�������7&��j�>�E��z��L �������b�wR@瑑ŕ����w�H���6�15d4��8b�Õ�S�u$��`�T\ATɼ�۞t�~��|?h�(������cጦ52/_xN{�un!�',�����Y4�����?����h~�7,�*(4=�q�n4�y�H��"�!c���7���X�cybin�A��9���>q���G��p�PX�<B��r��8Nk9�ۉ�)!�)��!8��⺀�˿ҝG|fE�M�����z�	ɚ-�!+�E,֗ʡ,@�S�फ�988�w���� �De�\.��K��e�;�S��f�A�~2ڶ$1\ʛ�����g[�;j���t}J��v�2��ƙ|;���I-E��݁�_®�m;���/Eb���A3�:����$ͷ�)��t�򊭆>�ێ�Ck�'�oK�8AΏ��}Ě����y3��w�u^���F�Z�m�f�R����0���No�W�V�p���h�Y��2�/RcV B;����=�,��Z��
G$���e#7U�z�é)�t�Db�4]��~m/��Û�LQ_�q��ª�zG��I).�-ڣ>�,��*����r�X��X:O��f���@�P��b4�I���%�,�5}\� ����e] �d=���x��#��(��\��(�&ۯb�PsR㹈W���s�x����O|q��Y�Ѷ�yF:��8�V	�v��5ƒ4r�>w�5<�~�Q����bʶ$7Z�CS�qub;����P�W�����n��JL�;�=���8�ɒ����f#�'`v��uw�?���/�������ѯ�6���礎K�}ΆO�W��T�мpN/��S~p9�H7$�ج��&���qCT��i�����+u�Eα�
q7�]�ː1��a��ߣ*̡gw'���3���%�+7�{k�P}�9r����L�h]��� �nkP ��w�{�˿���Xc�wY>�<Q̎�$��L[�u�����[�='5%�V��U�ݔj���IAS��L�^,���4��񴐈�R�d�y"�t�]ukGWT�Q�WX_��~�3�@�7͢ �J+�sh��%r@�Q���tݠk�s�vĚ��dB�!ߟy��R�Y��Rkk fљ�!za���8h�/Q�HJ�����e�%h�˱jki�HB29撊m:�w��M�tH����ǀ�9��̹ŵ��qt�W3����@�+Z��7�Q7��f�X:��k����)�q����_��=��:�#�����4�A1�2�kS��zz�s�'���^uecm������sz������j���,E���/|�]-p,��8�;����*B��@ׅ�l9B��ſ l��d�h�m����H�D$]�������$>�fϋ��VܝߧzAHh��ClMR,��l>���lLB)��^��s�.^q �T�C犨��'f�������3����{�W<�ޘ�X����.��3KQ�Ke�Fr�{s��Zp"���хJMJ�،���c�a]��D��>v@ܥZ��G�}&�@��|�m��u�B�Uq삹ʜl8E�@5Y��s*2-D�+
:{�:�Y$�?#�����O��l�L��"iLV	��:;P^k�p{�O�*M�0�&TC�V��z�UR�^��}��"�r�v`q�K��3Q��$�=$�b�:��\x�ȃ�pS�|��&�W��~��˒���h�F�G7�����$**�R��ۮ�;��VC�*l�ֆ�:
���W�����Jr[�;�0�~?�Ql_��]?�sf�|�O��Q���Z�i�B �CO6�0�@K�#���a�`��>Ԛ$��"�~��F8s��(��*$�x����	���㫓R�jQ��d6L�!t��}�#�	���hv�/�]�ȭ�΁�h;�ReN����\Vt�x:�.PY^�f�2G_RV��z�l�Z�-Ӵ8��ڴ!�����)�]���{�W�2��6�rH�H����z�_|ͭh`���/�DK{��`kh���BŰL��J��F���u��=�m46��{CN�tm��M0��E��"�SW?���,QҦ���a4zV=b�0�S�ĵ��et"�r��1,<�aZY"G�OS�
�+m�cT�=�]�02Sq�^'�;�:�����,�#-u����~�ή�b6#X^lkw�=��i-�����)���Z����� y$J�r�F��ҡY�.�I�B�A��[�b�M6N�T���o��F�)�=�x^"s)�B�Zk7T��Ǣ �R6��*��^����[�G���!T��fo~�;7�"eA�m3�1��qЄ*jA�>�ۅ=z&z9��(<���q��Ɔu� )�(.��<��:��"$�5ɇ��ź�,���Y:��s^?���}�d� c��r��OE����'��ˡ�[��o7��v�Kz�g��:�楨���p^�����Y0���>���V���{�x;zs�*)U|σ.��>�+\?�D��R��e�t���Un*t�͏a�=�M���q~a#X!�i��S{��]���)$A��3F�r���Z�漥X�����9e�U*�g�J�o!� ĭSb����t�J��P�����m��:�{�c� '{�R�vG2�.�xN�x�{��#{�M�sG2�k�_!�b����h@`�d�z/�T:���9��D�b[���T<�4�m�, ੾�V}��d�ž�tbCn58n� ��>ݭ��ϿEvtɇ��L�"�q]�_	%,䯪��}�1�;�^q5���#D��ݻa?�q��[#g+<H���<�S;H:�	��U/�i9�b��\3p��P �@;��Nƥ��4��S=�/��<0"�/к�q8�m=�;i��Z�a	C�ռTZ��V�h.�%"/R��P����v�N����x��m\�I$��V����Ӹ�,޽W��*ߴ�^+�9. ��F'�5Q1C�0��U4�GV�׉�q3P��ص��2q���6�%51&VH�^����]_Q�|�)�`@X��1fv�����y�y�q����kq%<O\��W:�ȱ���(��&3�艣�8X�>��c�����_R�K��
�52jT�o��3fEdбP�&�گ����=C�at�/��A��$`ǁ�b��K:G� ^��:h�ؙ�ߟ�qCQ�6D���������Z!�2��\���<���P��| %��I+o��y�6�T�*�˷w A1��MaA��T��(1|}���|�Y$ٿd߆�=t����D �����>ą��4�<���ҫ����Qt�X���i�3��8�T�3gR�m޻"�>~a~�pqF���PN��	ʚ���^q�r0�Y��@<$�!�b�f��xisO���XO����aA:X��`�0,)�RW˦e��BZ׆���p��֦��bž$��E|�q��\h�6Χc~���7�W�#o� �k ��Y�jD,�w��͚��(o�����sҡ.���x�Q���yo_4��w�;B��
��~�6�џ�:/k
&D7��)3�x���&��3�^kV��"\J��j!k?;�Ϣt�r9�P�Т-�γ�^֏�r�W6�N�p�.�[���} %*�:2�.�? ?}�gh;�BZʱ�&�^�Łv��|���R��5�mO���8��	V��UJ��{I�"c�M<��>�i�I>s��p���-�eT�OT����$Bin���E�Z^&�6{��{�Z��2B>rS�yr(#c���|"���D0�$�#;��mS�C4�ceQ�(��W丰�P`m=��߹(���HU�I��q�u��t!��d"p�17�:��|��1�;d���ϯ�AK�������o{���yx�d'����L�C��n>G0��͊*�}8fR���'c�x�F#N�b1F�0�w�z�\���1��\��i�c�ُ4�DEz�������Ш�:=�/��}�H������M}�BLz���_,e.�F��'��*�C=�яC9�P�$�lb�/�5����b���o�e/0f��Ȕ��|��}�
��\���Z�#F������E��V���!
����-����ڦ��is!M#R	#��
����-��͠�dwb�:�9��s��(��1Ӕ�0O�R�L�ܜ��x���sUUF�^��5Cg՛�d���%��r��n��ׂd��a�pH�(D_N��HeM�U�[��eL�R�ήg�^�Y�б:$�U����T���b0
��m�ip�@Ν�ri�vT+��9�Z��N�1����r�P�F�7:�# �"�J���L�sz0&�-9����3J,���ao��6��
�Bא�̴�v�̚��?�%QS�������S鿪��#8�I�cU����j� 3�������ww�s�BR3�CyyM��L�J�u5ؐNp8m��%@�HQMGU=��B��:�,�9�m)KT�N9�X	�֘ycX�H��_�cbm
�=�P6�a(��B������D�Oy"%��PZG �M['���mU�`�tpE��WUJ5�$�y�$�N�+U��þ�l^ਞ���U�!�]_Z�H=�$NO�
vh��@~S�(�����n5E�nvx:'�A�VV��R��r��H�	x��)�����@`8�������U�x��{�P�;6� �<�%?�g����[6���g�5�AP�TRX3���ٿ�2�1V(�I��Y�� A����s��z$g5w|�>d��)���"üuB�+\�[S�L�����S� 2:+��$z�ý����qhp�����i�Jf���@�����)HbF��_Fz��x����遭N����Y���?ߨ,׀�N� O��#Z�h��ү�=�#�Ƚ�G�)��:>�y�1NJ�]���R�c����nQ��sI�Y��Y����f!bc�n�:g�c�l�[kG�7��Z�B=	��r�w�3��>u�@� "�q��U\0�}���O�Q�3�]�1�( �(�;PG!D?�.Z���Y��f�r��J�i�k;�ue��JR�����᎑��w]q\rK w8�D{x�e�%��ql��r��V����u�QM�^�{iP�;gx�����=Wy��;������Z�u?��I�Y��e���5Z�v
?ZM���̷�W���&P�Uvd<�M�.#��6Z�n���s���Y��IHC�Eh=2l�"�(�J2���j��Py�nm̓;#ivv�SD�[%�z�f�D�Uڂ� ��9]�]U�3A>�C`�ZYdo���bynڎ��V��"��UJ�	B��l�A������/�"O����_� ~0� �۬�#��|3�hh����g4}6�]/�����O5�nvi��h�,�(O�5�߁���A����@�_@��Z��
I�҄�n~w78���M���e-mR-n9�����qx�e\�#VK�P�$񹣦���8#���KvkvC��I�S�G���9]V��B����O�t ��e[1g�=�:�_���q��:M��L6s��z��i��u�,�NIy	�ơ��Z��>ÐFͿ�#��^B1Wj�a�:+�Xn�,<�T�xI����;���L�&���&g���w��c�;���ظ�=�?]9��H˚�*�d����پ�<�s�Dt?"Z/�G
�!�㞃n�k|���݊.'��?���h# ��r���Т��Azz00�>]7���RI�n�*K� ?3fa}�S�n�}!h8 �0�����9�������Rl_8TO����;tմ��EEwL��a�?�:ݍ.rs<�qȺ���q����� ���"8��݇ρ��b>�CN���@n僿4C]��� ة���$��s%AO͗	ۨ�^���^[/4
��U���vQL��B��1�IR�H<;j��/z�!�4�*|޷�*t�E�\�"�rX�X >W ���^��zl�a�5"�B���L4�]C�-}��z7�OC��RNn(�cU\��c"�,��e�p.�.V2-����G71�a�d8�T5jg_��r��J�4���vt�e|��+U�e��:�G�����#Nr�h�/��B�C�ۇwg��]��D�9�L?����5�-�]<�曥G�syH�5��K�����"���Rw�	`�/BXI�F�v���*�@�"M�jĕ���o�� 9F������E����u��������A���gt��=d��?e [�z.��ql�۳�e��������Y	���� ;<fS[AFIjvmJ�N1�|��#����$���#�r[ ��M�w�y��F��V�jqf���DM�ٴ���7T���g�J�|�$G��[��{ޅ��˅U�{�Թ�<��_�s��f:�
����8	7]���v=X]�so;5C�����O���I�$�x�qK���}��h����N�ֳ�� 5�IO]	G9ʉ4'����