��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�s^W���0AP�<7b�HFC,�6��^���v��T�F�@3�e�_�Ѿ�bl�^��g0�1��檟�\�~2w���~g,A.�s2�ym��q�?����n�������Nt�T&�����C
���Q��� ��1�A��jw4mI�\�dU��Dm,8n� ��3ئ巎nE�|�s�.'Lk�H�eG2�&w�+YUF�ud`
D�"#�7��'�w<'E(�����e��[�9n`QԡO�!{���9|c)x`�
<G��I.f��N$.�����R�H�Hd�R_�M��U�Ι���$���`�����\��N�7i������f[����[�&�*L� �#�j�5��u�<�
�TT�Sa9�`8�-Ӆq���!�ݲn>�6�z�͡k31
��4���t6yBc{E?O?�Vvi ^�߳݉d�{s!���3��A$x��>Y�5��m��O��8]�/t����������*e�.�����ү%�W��79E�����zV4D�>k	uطWIA�I��g���Y���#v�KY��r���tr�z�N�>��^\l��m�$l�__��WMw%A��vU���^������I�*$K���d��!<DH  �<?��aSH'1��ld�¸�<c�b�˗���Ԕ=��36�z�Z���ڑ�|5��2���M<�/ �PḾ��Z��]}�6M߽z�ZvÕ5����D�/��=͑0Y�vt��eA����EJ�'�r܌rv\�#%.��ᡃRo�|fC׻p8t�X��X��
t<z��x�jXhS�����.��H{k���^9u"F#~X�ҧC�������ݱ�26�@��L�=�fo��%y~�6�yu�5�V,�"�.�l9\Fq �rR�R���np��a��"7�eɫZq%��10���3���hz��{N�^` Fu�uN���J����N�� 4~���gW�]yV�i7�����Cח%n��D�]ab�.����DZ�6���K��_ծ����K��]�u�	r��p�+Q�jV�(��3�8�:��AĮ6�+ei�۳�c����<�T0���Y�X2�N�����H��Q�� r����$�$�	��_�7���
31o�琖3�f�7�s�]��-wE���$�M�N7x@�I���2���Ӆ9B�h���さ-ZEg%���AbYg�v�����X�%
�I�U�-(����l�� �^�mm'*b�#�N����(�
X�p���l�D�0Y)<�T��6��1�$e���� �5o�ݟH�����oC���%E�q��Q*S.K���~]�Ie����`em?6�lf�$�����k�2+�]���W]�P��:�g�'���Oӆ{w$�U]�o���h�����
�RG���ky�����՟q-�V�v�}cs�=��ר}B2`��S��e��x[�
���|ؽ�-�߰J��w5 �v���E��s"�VV�h�I��G��
�GKS��Z���<��+"�/�Q�T ��M�st��PƯ�����r߈$�ۇ�X~ˁ����E�uB�q�b���z4�>f.�:����-dܷ����-��JwEdET�JN�-����/(ăNP�?�T
T��G��p�)�3 ϰ��Zq���I���"ˆ��R��l��,��PK�$��m����\&�o��P�/՟ ��M��tĞ{���^$��ǥy[�����R怼���QܰpViB�t�Z��\9����ٱ%
���
��s�)a�M�'���(H�:uB�j����{��2�V����h��I�v4lw��f,�����ހe�3��+1�ozp��o��a!���r��6����>�  Q��v:1V���[�y �(�����,��D��'{����d����J��!���r���Q_@���Z��i:T53Ӻ�Yh�W��4MK�#�ʤ��+e�Y)'�*��6����pxz�h'Z�스���8HjI�{�x�d�R��b O�� ��G=�VO�d�OB��pz՞^s}�48\}e|�QLAT��:��|<� 
���7!j�����'�t(^��{� �Z|��!�(�����	<]����2̌��6�,?:�S�2�GnE$e�R��RD?��<��WOQ���P?���(i��=��s&�������!��@�¶�I�f�34��Un+/���tV0p(p�;�ޭ��w	IYG���Bd�FH��v�-�Zb����{R��.ĥ��&�/��B�mI�]�ʚ;��{z��4+�|WC�씱�K7-��o��M�j���׷+/�Q���E)=#�;k}�>r�D����XF#7^E����z<Su@�#&��(�a�j�V�7����`������bRW�nj�K�㹅�9F��>�8������ÙĞ���,�39�C0�t�m��W�80}�
�G�H`�����qH��qq���= �ǓCI�z��|[�8�VPp��57��}? Hٗ���d=�Wrj��
ӓ� t��%�!�Y�Ӳ@��Ҟu����>�J�[.�37��j��AH���0.�󹅓�5��)�灋�E�W�o��G��5��1[s��K�h��0A������V*PA!;�)9� s�Ăi�V:dhh2l�<\:�x����HY��	���8�u3�ln���/Zh�Th��fxsc�@�0=��x-#j�ב���
��r~]�/м�����H�+�[�T[Lu��RQf����8�8����t?S�[�?�?%DDo���_��G#�4�����.R�P��p\��I����wthzZ�?u ʮ�&jcߢ�����t��Q���,]�B����(`|�~��
��/Dj}�~��V���n�8�(+�~$C���*��<��N��|f,���t+��5I�r����(CD�$�ø!�"�l:!UIl�V�'v�8ސ�����LZ�#H�j��dひ\��fu3�W��0a?J<r��/~5�hC�aHå���)��+nS�l(xf���|�ZʙyW2
6�����U��������;�:�Г50���=e����-Mx{#���?BG�;[�gm kG�JC&�,�8~�w��X�r��QD�7��T�]��Q��P��`@�fa[Y"��|b[Hw_�"�9�p�^�J-���e&��Gz"�ݎ�3<!�'��������f5 ֽyɩFK��η��
DčS��	k��|�L=Ӡ1/�i�a�<��3	w
�������dU$�տ���ӞF��dt����^o�ZSo� e�:���oa�xe�̫4C�#u�M����H�����ɴ�j����FP Ph�%گd�BaA<K��zi���6�ؓ+��nŇx������� G,뇚��]=�u]ă�\5> �Yo��S��oA��Ů[&������@�zk�D��� � W�[%j���҅��2���/Q�v����
^ҟ�+�Rge�;c�^2����)&F�)�2{g��;t��#��
 �D ���88������U�A'=���ɧd]���G�Ԩ�̽����z��hn�OG���T��&�%�@�`�����K�<�G$�=��W�r�n�h�{��c�0��{�9���UJ��`b0B�n���_�!��y�E�Cs ��O�״��6^�g�b�/=о����Y�_@#to�d���,��P����޽�>�9r�R
Kj�+U�盇Ti�9�Xy�����"@$qO����͂��/e�_����4�����\zqz~�D�Srpu�yc��+ǙC[���e��mxk�dr�+vk�X�@���������9X����97[t�TRԇ�m�"J�.���u� ���!����.A�]
�a�	i��)Al;a����4��t�P��+��x����kӪ&vTi[|(O1g����D���ED�[3 �,��t�)��QC�\;�Z$�P3
b�H�{?��vW[���NpT� �%���,1��S�P���.Ro���?�yqX�^����������Z���]Ӯ{1��ޡ���M�U�M-j^�[T�p�~��+���4 ��]����muT)J��*�Y��ݐ�-S^�9��F����γ|����z�abo�wc�#����fJ���Ճ�����@����<�z?��E��(<�&���Z�M��
�~]7����8�/��Y�EiJa��9����~��B���E�9Ӫ3��$
F�Z)�,=��l��Ō��������