��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0����R��@��77�c�S��L��������I�4��ȞX܇���
i������Pݒ=��#S$'�V�=%?>*��
��?����������� ��Qʭ�G�E�@<~�~qߨ���/'1A�V[�L_��II���f2��T[�n�ҚP} ���=f�X�|�9�V���WА���;����z��-¬����e��ߕ�d���۾�]�c�>&v�f ��ג��T,;�0�"�/,"�? ���^�����,��u賮�G�WEg����ab��͇�� �9+�����P�������ƈ)����n��5�����F�����G�s�.vϛ+�[�<0f�yˢ�}XG��)lp�K5��,��>�v�*X�Avs�I��sb��Զ��)'3�s�b��餆�JY���=+3��Thӈ��c5g\�XV�V��mJ��P�����.6����OB��H.H�QC3K�Y�z�0��ވ�ˤ���elU�	���_8���gX��+.j�kXh�ϥ2���gu��ϐyD�&;��c,��N����;hŖ���^tv�?��&��^����U��X7laSFA�i�t��]G�3-L��� Eg��=P7 ��f���Mq���i���⦛��jDN�1�{ ����x���<�xh~T�����=����6���=�����s�G:��(jg<��3-�P�Mp�`�m$������PLaB�S>ϱ��=wS%�aŇ���3͋f"�ri[Ng0���\CV�<�Gx�|+��oKx"�i���ї�}��}�>BH��YUb������?��T'�����'��~_���r�����p��~i�l��\�y���<�
�ԕ�m�k˱L��d�� �� �7Ð `�l ����w���f������������>H�и���A*��W}�����|���5E����o�#��ԏ.WN|���ˮ��v�\h�B�%8��m4ͽ�m��!\��K�RԂ�@. XJ~���q�o�3���x���#n,J��Aֳ͂^{�����5�5�r\C���b�f���Ub�379�������k�&�F$6��=��\(�5���r��JN�
�.������)I6��F�g%e�P�.�Ը���n}�U��yu�D�Y�!���%����R���Q�Ӧg���pR��e������jrş�{	�}E����0���Q� �k��W<`��86�������]�@�aq��G5���e����wߪ�I�Ɖ��O�Qa�A�cW	x�|(��o���9���Za���dBqzJ;O��X�q����K�1��>_�kOmѱWJo��*`��)�
���PhV}��a���j���"N�͜����6`e����c�j�t���-F{�<�AZ�@����ЭF[��\��?���O
���FC�{�+��Qh25���ݻ!�ܟY��-�an��L�A?Rܝl��Ҵ��MU%@XR5���\�_>�7��X��4���B�h��ּ_/l���/���Uo�v�����;����
�%��)� ��^�m�\��_���L���:u�@��h�ÂU��7;�`��e{T�v͛!���MЬK��� �Y|��g��ų�y(�޾�h��0���L@�ۢXp����������s����-��7Ĝ������~t��沔��n�e>Լ�L���0���`����¸3)k�"����}�^�[�y9�Q�|0VZ&)G����[�hSƘ	��#��Z'M,<H�P{�F~�ZMDv���H�i�����OPyx�.�#Py]�$�3"���|7 &N�@ӷ�����n6_>}N+�""�m��U��͇N�=7"���]I�Y����v�V�[q�itܹăQ��-�^�Ɣ�n�3T���]���*�&�~E��h{�p&����wzg2�H.M���ic.�K��4����_	����5P�N�>3��VJ� ��;�Ek�1�2o�;�6D4�Ow�g������0��M����Gc
f]2�H�����TXP/vr �)j��	a�m�k��a r���,��=`:���z�d���1��8����{��Lӫ][1q)z5y �o��$`�����}��~Z�!Yl{�]BG�oi�)6�pU�~�G��#�0��ʞV@��!-h�SY�Ѷ=8�C�v�ǜ兆�U��Z��Ap*#I����XƉ�DO�C��S�+��TrIRp���ܥbfU��è�0���S~~��!.}��
���w�Dkv�����T��C��p�j6�i8<�4"��U��!��Y���+�Q!��8ɾ�w��̱�JrȨ�k��׹���TBb{�8ϖa.�ă W�S!(Xt�l&��ոY��ړ"�=�5O��8�g��X2�j�k�YwJ�&�>za���#�0�Q�{2%sx'�2��޵��C�.���O�
;���m��hy3�Ai0sɊ���Jh�F��V.�-n�g���)[�9�F���󡙮hz@/������|�&w
b�g������
�Zܨ)����u���-��? ��4K��m���tc/����]Q@��& ą��h�}�;`yB��A�ľÞ���e�u�U����)�!�ޢd+Y��q��?�J��	?^>OA�BX�#��S%P�M���J�Wc)r�����,���K]�|���jl��xH^�X�͡���(|�L�z2�Tw�r����Y(�<�4��x"'c���A5�M�N��/�ex� ��E��X�[�^Z2y�Mz�n�
#1��[H��o��p�����o1��]U$H������O�{��fq��~��$Z�`��a��\9藗?a�"�$sx�v�q�ǩ�]���ðb~����MS�{W6�B1Z�&�)Y���?�%���PT������|��F�GV��K�o�ӓ�2Ȓ+�XY�~V��K{�T�p�����@W�:N*n(������`a���D��5�ݬ� �GY�0_�<P���(���!P2��6͇�v��&����t?6�S��E�8(�
�}kM*�!�f@؃9q"	�ZE�"^�~s��=�?�U�Р�9�#C�) �[o��)&W�[OTl(�����:8���g&'�>2�DQ2�]g���&p�S%ꨇ.Vջd)�9�P�
�u�(n��;3�_囼P��"�3g��o.gJp��uK�WD�9
�^��z�N���uj�<����F�;k��/��<ɨW͘���E$�1E�ČV���U�D����[�e��+��qn��29�>j9���7�=$?����P���O7W�����O���ѽ8l	R��hvMG֖:���A�ĕ�*-��/��;�})bUJ��50�l�	��Ϩ���s)���9=�g��4�M�~B�u��YJb�B��>wa+� �>�VFi����i2t���1�[>��X�����5��:���2[{� !a����A
,ԓ ���ǵ\+�yE�Ζs��jp�y�0�AI�A�w��?�(1`��!�%u[w��pR�Ч�v���@C�Ƅ I��1�{Rzy�F"�X�Mp \�x^U�_🛐v��G9�%Z>|a
i���z���R��rf�ɏ��Y��&�+F�>���S�z@ˏ���_�F��p�A���� ��:1N�m�J�J99��Ȯ�YD�Y9�ғh��6-�TBA������Q��E�a�`H4���5����oe�^���a�s6����D`�P��_����cA)�����L��A�x���@�{3^AS(���������\e"!1��(�˭+�s�U�+p�W��e�I�\c��6[�R���e<W����O�<�̫侞X�ګ�_(�p^��W�& Av���}v2�L�9����@�nD 6Bo����ΤV����+��G(-�z�h�mfb�1Bo�_��7��%��@e�_J�d��z�gO�M��^�e�9&�i��A������10s/�8k��t��1
B��ů���|Yj�#�H��V�(���![�~C���%oe�T}�	��_��]]�&��?���}y�zf���ʖ����~��w��F��RD,r�Cm*�*
.D%Yo�c�mk ���s}����]�WlaY.X���W�0���||)kt��Q0�K��2: s�$(˲��S��G��S���t���!��0�ɉ���FZ�[]c'��ң�K�"��=IU�(ЭP���'MK��ƙ��	����̉��y�y��r ��5��KLDf�M��ͅ��H���ǶŇ�K�̳�v'���*�S�W�δ��It�Y�`��ԥ7@�FJ��|���H��4����� �N�̻a�� .��uOk�O
�,u1���c�і���K#��p֕�x\���t��}��².���\�0�md�/셵�}�H�h��+��(�A���ۓ@^B}q-	�M7SO2�^��BUy͉�鲫֡'&Fn��H-)�Ձ-9z��i��Ё$.������bpQ�`.����ROf���w���s�o�S��L_. O`G{��b�O
�jLoP��#����	ɠF���<$ۯ�M�S%�E��R�睜1�-a\��
�Y�T��桧��<q>$���誽��9�)�v��&f���NÛ�(r1�`��%�{I=���#��h��.�%��CH.\��0v�'�����E��:��c�E��|ҥ�c�rP@����K'˽�Fe��H	���Q�����U�=�;$`S��-d�_U�i!.Fѵk�}��n���Rߋfg��,��D��jx^ �i���3� �7�r-w���f�;�K�ky�Uu�8��|�e���AI`��R�F��x]Z��)��'ı�,�Z���Fd2(��gѾb�H�DQܕv�`Z�lj9?�F��V��|�/7 ��I~�Y#?�\ e��;Ul`T`�����xp$ֻ��c����g�rU���NL�r㫗n) ��፵�t���`*��*��w���8A��I��QZ�:,�yC��36tp\8�]g1�D��h�TAp�Mc�~W5�5�4�j�:�˻Sݗ�GWֿ�
-@8�p"ڡ�Ĵ!��{�7r�N6v"N�H=Z+r+-�y��|aY��HV�M���@HI%K���c�@,9##���/�m��t7F@�-�c�D r]@5���b�˭��K.�����,������!��c	c6���)9�����j�-"�#7�6�
���>��q,�3�)n,�::�B$��' ��i&���-�-喇O��6z�Q~�#�dh_�M���3bs`���=��O��]���i����Y�.��⧃T/�u����'��1�ޡ��a��_�;���:}D�$X� k��=�x@��\�Og"��o�Bn�r�V;˫�d�B��,�P�r��I��n$]��{*������l&��n���iE�pK���&.�8���/�q�Z��;��Tt����	�[��Y�����&��h`/k6��&��l��{tڨ94������e/��� *���E���a����Q��a������x�����p�~ְ-C[ ��G���J�Z�Ӭ��Bms�?��Z��T�}��=���?��>8�gx���2uA� ��|�X�ד{Z�\���@'>V�B�$�N��r#����.@
p�/X� =Uv6��d�1D]�y��r�+'�����@m�Rb�N�@���w���k���!�uxf͇���*��[�����ţ3Ɩ������v���S[��$��7�:)�$�\��z��Β���E�1���?����G�@�:Mm������ݱ�ɠ?M�[o��V�T�0�g�������v�f��[JD�������Y�� ���tP�QP�Ɗ����\ß�72
ْ�o1ڣ����oB�����PҰ���בY!�C*���D=�˻�{���i�MA����\#��&q���I~-:�E,����؜�O��_�Y�����Gs�|$Rv_pT��R̈́,�L�h�_�o*`xS�R�M�'%�M���d��B|��2e�١ＨCRU��'�A��������ͣ$�Jj3��(L|Et�X(���>A�Sr��[v��W��}�a�U�%Ͱ�ρQ�^.+��T|2R|iU�T�"�-|G�VҔ�����MT��/ ��M;oz���P�_x6� �"� ���Fc*�7��:Q���-n~�.N侑h����'"�zK�o%� 5�����MJ8�o����,��x�ogE��f�k ^��S��W{<*ZZ��s��Ÿp�V�T37?��꺿�FĦ�\Ԫ�&��&pC��7# cgVxw9�w"��E�J�	�Q`)��\�n�����
�"  �;�H�Q�(h\N�r-��UN|SQW�ܺ�?h0j�QK�[����;��2+�>>j�:5��0���\3���t��Sm/���Z��D�!~��:����${@�Hf��I�Q�x�i��~��6x??�=��̀>��
c��r�F�P������k�Wݟ%�^����"$P���1G(_A��&2��P�Hl�E����W3���~`o��^CJд2Z�6P�7��E|Gu���a�i2mB��<�EA]�3�H-vo����;�+o �.H����+/8,>�mZJ��{=�����_���"�
���t��!1�M`ܵ�aq�{��T�v����9p������E&'E1%�5�Dv�;�:E��K?2'�Dd�7�VD�F���Q=�	��+�y}H�q9��h��1U�Y�("��w���#�-�w�#��4!��ג��O��UPց�/}�V�v/��m�,�6A%�$��\X��\6���!�I�}�,�
I#����sUe���z2����'���k���2V0��|8Fo���vKEC9}����o����ww�ci���!d���o$@S�El߃����va�P�.6S�L�k0�?xs2{�p��Y�8�x��O����F T ���,���gli�T�:f�,���!p�f�p���*y�߳e&��w<�� 
a�F6�@�,�!�!�+�������|c.B�.��>��^]�@�¡
�9ɭ�t��D�#*��
m`����w/�n@��Dg�oiJ����+F�R�d�5�@���n���˅gT5�QI'��cJJFw]M φ�i���_2����
�R�/�]�a��V�#�ah��}�H�Eut�<ӽE�Z<��V0�b��3�'~�E�Fq�ԲV��qrq)�g��<Nd�/
>��!$��F����T�۴���t&�@�Ŭ/R�e}����ق_����v&e�p1�"p��=i�GE�]����!��x*;{��&�x�^g����|���)̼�[��������gU�	=��5����Zn��_$�7Ο�ۚG��j_O�	Vt��a����C�}� gT�5e��9(qW1%�	����]��AD-B.�Kk5�U����A�`�U/���.j'f�����������G�����W�o�V�����}[J݁�Ka�Lu���D&�i{Q^q���uԍ�%��v��Q��v�	F_,��i�!~�M2��Q��h��	�@D�)�:���Z@2#���wds��O��V@�hy-TZ�Pl�X���=U�ƙ�;���_u4�٫֭��E�G�{r,	��J�@�K�j�T�Ul##��viHVN���7^澕�NyG1�a��ak4��e�]�F����r��<�Oy�%^���B�*�]����%�,��N?��][�y�������=4Y�k�	x&����Rl�}�5%��|�b}�u��zY�L�q�<�� �|��5���,�m� @{,���ف|Cpu��	7
�i#��	�G!�U�#(!�(�`K�NI�lۄ}Ù*�.���O~k��v��?�$xm�5�_����5m5
�O((�8�	�t�a-��n�d������|oD~˷�Q��c�yt�9��]���ȱ6�pEO#�CX�k��Ͱ|(��9Z*�ƝeP��&��y�Lٟ��/��vt��ƺ(�#�;�ޔ�Z;*��]L�D>��L�8%zA]?X�%�H��2t*�)�-dz���D3#xSN����s58v�S2xKo�U���SQ�ܻ����p:ϡD���P��$��n��5ET��*�<_>�ؗ`��Y=֟�ޢ�Ґ��G��9��][�n��A2�q&��~N�F����Ҕ��MI�p��p��b���f$��_=��#��8e������ҩcr6p�OʖlAD6f��h���6�E�}����IHy��!�h��)~���t�L���J�[�m9H�Fw�����\9Ng�E�dh����u'O\�p���DG�M���xj��1��֫���|�U���:�Wv��� �6��c �|d�p������x�Յ�Y����+���Pgs*c(�3қ��&�������%�������_bv��6>��8s�|�gd�,GS�8����	���@*�^�sϋtv�����3C ޷��Zo���]X���87v��d�A�T�$��K��#-��K���}��taMb��3��V��y~.0��P���X��v��f�$�,W�C��I,ތ(ŭ�j4G
l�(�@U(V>9��V�xK&=����V�dL������҄�l��|@+q�F�O�m�H��,��84�A�S��{����Ԇ���~�&8!��4
�t����Hjw�2V��QQ���1�N����d�U�b��cB�v��w��A�uehyܘ^t�H�cQ����k�����F�p���"��f�	�0W���\Ҳ��P�}Lh!Q'���}�KB��=o-�G�#eu��K�e���gͦ�G7c�Ԭ��a��82^��i����[���rwmf�v�b��^c�B�h$���&3!@]�s�d��-�� uKyjT���nbT�����Ya��8�3��{�F�<�g���qȴR�g����lZ��s��K���6 �g�ȩ���D\�O��X�5�(��OPR-F|r����D� �J��xt�>�N�V�������	��Jt8(�\�='�^����\��쀁"�w����Z5��k�jq�A)ĥCp�;�J؉6g�޺0��݋�KV�Pt9!�͡"�k��h�}Mc�ہy<ǳN6��ݧGM���W �m������*�K�K�d��XO��՘����۾Ϭ@N}8����[�e�Ҵ�������93�R�&دn=����,l�Z־�%\^ݴ�yf�!�i��R�=�v���)�d�%��{w��if/#i;�тU�r��Ǧ�.�:����({�a��c��館 x�?=o��Y:��(��A���k�A��4���}�@XUQ�m����
>�f�Z\x�%���ک��Ơ�OF[��*�+446�6w��Z�+��ZP�k'6e��<Պ�����BuQ�ш=�7��cۢO6��v��/K�ޓz�<�(�g�@U���E��,ߪ��ʿX5����`�~��J�]g�K�A�Wl7��Q��Ե�k��Pcf��wP
0T����>��^5R9V�(�̖����X��BK�ɢ�zղKl�O	d|��-F�=���J)8�ڏŊ//{�؇7�@g��&�Jt
kD1F�;|�nE�Ÿ����N��{)�w��E��(_7tqQ�K���$�H��@����ˉ��,�7������1j\v��Ԓ����7I�$,[����@��\�;ݻ�e�|��@����o�<�0:���C��U���0Ur�\240��D@q�� �t�N��N)8�!�G��J�@0׊dM�Xd�o�k��wyA<�Z�~w�q�t��0���C1��ܙ������p���C�O���K<䶔�G��_��ɇ9��<����Iր�ˇ�%	F�_1]���HI�mˬ�m��3�{h�q�vz��+�l���͵�T2��Ҍ��nQh1*U0@e��bL�
�ϥl,��	<@]n!�Zg���8[�I��b7u������ѱ�'X���;i���qjۏf~1��Kh�4���>K(
�����S�Q�e�/�q��������_'��.�@,�"�v=�s����~���3�e?��L��+��QG�D��,�P[�2G�[`��zS��_B���1p�A`���8����N@BYXFβK������_�S�Ӹ����.�w)�x��%X����G��g�>[$�d6��E�y���rNwK6'���!��!ӛ��O~B���jڒ�D�O�H�YZ܂�
ϻ/�� I�갭����S}jb~zN�"b��WG�}�<\��b�\���� ek�/Y������|9���಺s�ϖK�G,G�W��-�X����V���fBԐ�-��w��A�zkdH`���&�=z��ǵZ��-b���Ϟ�5GR��p}�΁��L-e��Nc*d
��=kk����a���,ߥ����y��.8�p��b�
Dq\G+ϓ�pO'��q�z	� J̾��4�c͊����f���y����x�b��鍉9 �CS��8z��/��:���Nٮ{l_]��Յ���hVu��!b�z%���)�6��+�3� �9��LM��0��3�5?ͩ<��Dƌ1LﻝhC%<uk�3�"0��������6���R�|���ϨA3�u�g�2`~y�^	# �G���1�5U��ĲM�E(я�a7�C����_�f�+�Rϥ��/����[��AA�@��%6,u����栚>�w{0�ս~���E��9����2T�r�W�ӈ��g���+�Z������;���g�0%�:_hhuQUF5Ex.�H��Q��1��o�����C�		P��Q9r������FF�Z���.��O�ta (AJ�(tܚX�{^�pɺf�:O��u�����p	��$v������=%!kf�O����*����m��I\��7#�����-��3%���`{��T��̻z�j��G��1�e@��ǀ�(k��u��_�+�m���6&_�g��A����W��ߵ�hl��\�m��������h��so[WS5�w=���Vҿ*S`@�$�$cb�<�'����%�s����o��_��,*Z.DB8y�� �]�++���/*h}�&Z4VT�	Ez�� C���rM}��c�ç2��PY7�W,�v���/Q�#�jȘ���RǦ��`��z��v-������x� ��"��Z4�|\󚬌��$�o�/+١���G ��j�k�3WRҝ�jb��Q����Z8G�)��5�ZIu#9�t��h`Ċ!b�j��&"Oƨ��?~��z`@�U���0[츁�')@�{b�	.œ�)�0�?��{X��;�?������d����*pPx�һ@6Rw��涳[�g��)Gb�@s�'�0��ɂ{*O~7yh�!�'c�K�V�/]�1��;:�&ߛQ�쥝��Ԫa������}�^����5�b.A�iҷ�l#l�յ�����ǀ�	��6���Q�0�+#c��~��Яgr�/$��p����
���l��.NcqޠZ���$���#�22��G�P�A�r���0Aʍ��U}�t�^Д�ƠCIy����+X��S�4 E�zE�D7�w�02�>-;'mCy_6���K�ĀA�++c6��Jሢ2ce�L��g�EU���`�$��	�X�Cb|Vz�Ų�(CG qp�Xф�����0g`�{�	�৙bm�!5ơ��Mv5L9�6Q͡8��&���42��b�������B \��Th���D/ �<(�opH���_���
$#�ΩkJ��z�-7
�#F�dj��������T�ٚ�����ұ6ȭmvT�I�W��TX�'	%�JjJ뛙�geyagd5�0���e�^z�6a :n���R3�R���K��WB�ݫW�~r�x����!�~��	_��y%e����v�&�c���5l�xˏ$��,s�_����cG+eN��3h���3��M1Y֍O1���6�]#���l��wG�&�?�2�KS���~��\�ҎŃ~R H�W R�"d_x��,��8�{�K�?IՀ�u��hF�A�eC�ʧ>b�2�륵=B[�E�����#�ſOڝ��Ad-�hne����5KX:�q�ŷ۫�*�R���;�E�|�k����Y��-�s���V	H) &��,*���X
�T�?���f)��?�E��w�d��s:�L�x�"�G4b'fdT���	/�I���g�U7�p�]�s�>���ΡI:46�*h��Y	�(/�o����׉�+��~f���GEiC4�E-�(!y�^�oq�<��N��Z���N"7�1v*�s/�KQϡ.V�e�e?q�_?�kJ]a��%��Փ��f#zQ0 v��M0����V�Ou��i�Sk_,U=�����\�ʠ�A�F������ɦ@������w�(J��>�fSd0ǓY�ar��Sa�sq\tY|.�B���v�=V�&�F +�dk�΁���F3�b�}���]hi���0AZ��ѡ�g�&D��d�����3���P�mv�S1�-��� ]o��$ A<'�w79}n[���-���_H؋'�k�oa'0Yx�{4q������`s�x�꫸`-P>��;���%6A���Ɇv�%|��+Ǒ�+݈��Ӻ6��>�B��g����Yzݘw���ϲa�����-Î��k�<3�����{'�b� �QѦ�ש��W����gG��چ)��-$�PЄH-������L�k�[4
��%%�w~��5���8ٱX�̂�����d�d� P�LR��`L�ѱӷz;̵-	�\ka^!���~�Q�T�һ�>x����������y�ܚ߈-E���n��z�������b��8��̽�vc�T�����dy��??6���"_��h���qmH�P�~::x��ч/>	x�bE�WhY�ۏ�_��x��ru�@��R3��:ʘ�e�����ۆ��l$���*��ܝ ܀�����U�a�Rh� �uB[�}%#*4Z���v@S��QKj�����<;_�eD��As�W�(c�8V-n&�+`2���Q �9#RD���}� o$d��/�P��%u�5�,�+~p^�8�Uۊ�j�(�mJ��{�?o�Nw4�O��E�m@�N5��r�;�7�?��a�6l{�t���Ȭ�Gt��}�E��&�m�$�
T���h
�8j=�TMŗ�`
kF�,�������@���d��v�֭1Z�Qr5��qo�"�����w-��e�7R�f	<ZXO��/���
=�G��*�	�Bi?}���i���nv�8����_%;S���	�$�$B�v�*�z��R���"��k�.9ad�F���D�m�_�h���J�)���q�4n@GV_k�.�ffϩ�Q��&�KM;B½Q�9�e�X���}�mh��C���A��������y�,�H5� 3jȶ��͹�l��x��o����u��ʱS8�y(�iA�ơ`ͨ;Y�����X@���'×�^�%���(q�h�7�I�=sf�6��%?�ŧ�r}��1�{[��&Q�n
���(ظ�d����c�W]ʤ&a6���R??��Lw�(u��B�_�0��-���Z��y�� l� B�>�gڰ1���Χ�:�Et^y�[Y��JMn���C����R��t�'9S��W:��yn���'ⓦG���z3#זTA��n}��t�O�*��"D��7+1�.�|��t����{*�̦��!� ��׆�Z8���_'���k�f=�T�^KaF���׏�\Hz�W�e�R��1J<zqt%��uA�v4�L�����3M�@���hO��䃽�̓�K �h�����[F5�`��R��-C/a��[����w4�δ�l4F�J8�I�P�TN�dp���+3SX𢱎
}]$�v$�����+4ݐW˰m_�$T�[�1��(�F&ί���D����.����3أH���b�������lY�A3������գ�> 2=�[��˴!�Hm8(�������+M��n�Y6������}��+,������"�2s}����G��b�9_��^�-=�H���=���4gdj/*�^H�>��2�Bq�����du�g�0�p�]D���Ԇf����!;�ƴ~5>�br�4}1��OǢ}��c���6V�RfB��[����T*jEei&z����2�V�zx��r[�r�-�G� 0��)"��z��$�������(���]J!9���e
?^�Lx!`��g�)��BeQ�M����^�N,�7�W��(�x�b���
��r��d�}��߉C.Ѐ�:[kk�o��ǰ�&���!�1�4�\F�X0/���2���������Q�>��ε�dw�Z��R�yDԠNy�Ŵ�Ћ\�������&�,
�=���;�Z*L1��uc����ym��ԀRx�P�>����>��u����찒}[��@����Ϩ�5����|P�z��#��t���M��*mc��F�N/5$�N��X����irl�ޤٛ��+�x���-Ȑ> ���X?��.�'���Q���g���Zļ�]됂&���7ӌ��'�@��=���eظ�,͒"��Đ!����B6�W��t�ŋ�Q��Z W���}�r�{1���Ŧ�
�)��f0��:�(����41h��)��7QQ�D��U1�g%bؤ�ݟ hV����t��j�;n�a�ϴ�5@C�� y�>����`?;ϭ�ś�"ֆoH\L�&��T;�6m0֒�p<����c�}�k��\�#BX稔-xx���$e�n���0� x��p�ҟ-GO���O{y�p�>D�P�O��&��)�{�F�m�G�j
/�A���d�x���+iJ��Xӷ?�S���F�B����p������NoS�����PוS�r0�*�`q�i�Q5��*�����d5=!��X~��u���]��x��8L6���,ym'[�X���U�@��uaU��O0��!,=T/e�������=0�#Y��t��}�?Y����2 ��?��o>����H��)�L���������J��G��h�wt�P��䅰��ޠ�b�����E���G�M�����ߴ�nQ+jZ"��X��1�<��4���W,��=�P�����-���o����4{��gG��z-䜶 �s�Fs`��� �]��A�o�E�������*a��0�\k����o����%�m�P�t��_�aG�H�[�pIIo���~<<����}j�e���i��H	�T�v�]�$S(w,ܽ}����rc�͛ IY;7r;�(q#��z�<��Μq�7A��]y��ϔ�(���Ei;�!|��/��`���DR�.ꋶخ�ʉP�5];Bl�FB���$�����^�32+�/�W�R�����K��Q�Ä�jU���|�1+֫�P�
�M���g�K7\l����6�ɵs���t*�rle")�f�0�����GT�R�i��߆K��v�,T
	��g�ev��Tp��B�z�m�e�{O���ф{ ��_;�s�wCѐ��؅�#8V�D�GPg�G�%�0�8��ҦN���W�$��?('�1�{Z��X�[�
�Re>�f��*��)=�͠�/��B��2���k4��O<�n��?����f�`�,Tٓ<��"������^�ÿ徖��/Y`��43i�ۄH	����X��Q����"v�q�!E��ȈJ?�7�_h�f"z�uLJ��E*�aY��R�������9C�+W2	"��D���N�7!���_���G�Xk���/�1���RC���l�1���yC�d��ֳ �w�
����c�)��Z�f>����RJ�h�S1���ޡ�R@�M��0a�@c��a�5S���6$)8x\Ɨڀ+I\u��=9��6D��+x�싱G�=�t>%+�K�9�	�T�k�ʔ��]�t�r�~�%�`�&Jx�����g���:�Lq&�T����M����Ԁ1�xOՃ��NX�尌���:8����(��xC�և�z؜��;�2��?�|��湙���94rR�k|$���-����^�==��R��S�;"	AD�2�g=�����	�C��`|[R9H�^B��)J(��T�-�v��Zx�H^�L�w�k�������q�A->
��u�}�ߧ�D��U��b��>����ہ�y�E��7,�^���e���(c�7՞L܍�V�K����Su�*�:]�
��'t�]�x��u6�6ܹ`��.�;��=�{�WKO�����ז��Y ���6z-��#1���q˅��W����u"N��a+Ve
�U�~V`{�lD�3�����y#��<�؂-d�n�Ӳ�"��_H��kEc�g%�Rd?�.ȋ��%�[LWa(]i@��3^��?��x=�WK�ƍ�$+{5�f�6�J���2Ѓ���~��{�ܭ��{�d{���;�zۗ�R��38h�՜+��DQ�:�����֍�~������$����E�;zSM�-3P^�?�_��Ց��޸�~�d�wyesrR|��d�h$�ͨd^�q'��Eѕ��;r
�hU9������q����m��8�.c�%d�
�V�'�����7�s�!�?6p4�5D�_e�͂�U����=�w�J�N��!R~�ߑ��(�
 �)(@���7�YnpMk��1U7�X�P�Go��E��"^�'�ԞO�󔯚��G���YÚag�h���`��t4��@��"���Q��>�'���Ncss��$��U%/Jg��z�,5B��e4�?�a���0�8��.[P�Ѳ
�9�K�o�WU{�7��'N�[6P`��Tfd��������ݷN ۯ5�穫�i���kr��TF�a1�t��������n�$;�� S��@���ǟ]��^tyN��cB�jǚ4 ~��r�b�&0>-��.�*�P�հ.s�Z���4L"�#�/Ƞ��S�mv�'_H�]%�K��V�H[�x?�+Ck�ij'�
sПl;��?,t;�J�Ñ!a�_�X�!`�[d]4Z���	�/��S
�!?�,U�st�T>�	H�v�$�c&��I̅GE`�&g�� �~[��^���=ήk��r6D��Q��iW,h�B�8�\V�����Y8/{C����M�o�y�;���*p0Œ/��H�ߴ�3��R��U���<�Mon��U`�����Z���K]�$E����,��X������N�Q�|n�$oN���L�A�JV?�jnޓ�u�$�W�M�;���p�Z1 ���t f�[i �𧑎3��7\QVL�G
죶y��J旆 ���2���cv�}p��g�oG�M�H\��>�j�V�<tW���/�z�k��d����4��8�΍�6�3yL�R$�A,�D���w�	�bWW�>�.���q?�n�`jZ��(���8͙F�M�Y=��>�.cB��\�~����)㼌u��!�4o��%*l��IpF?2��Uu��P)[�L t��c�(V�}љW���J���	>��'�,��e�O�d���z� �-�8T��n�9�[w`7D���e.NY���־�򎢦[�����b�~V˜��-����rL�a<�m�Zl$�nc��A[�3K�hm%�uʙ=n��(�GD�魣��Id�S@��k#��y�������k��C��82K(|wu�6�1���FS�d�{��&��	�%��Fw�A ����8�c�4�QڣYW/	�����-ֿ)lg�4�ٷ3�̐R��Q�a����MM5�g�Nv9N��:}cFY�tu+5��v��dչ�`��,:��<����EZ�i�F�(F>�	�4�Lʗ����A� ��Q=������ОGB'����Kf�!��H��cv/��$ft�.�~J�%��4�S�O���hCܤxoՋ�~*wr�EᄉЪ�u����*��^A�ӷ_k�TJcjE�&�.ҭc�k�d��<k�f�bbŹ/�F���X�����1���a`W��G��|�#[S����c#����5֓�Y��
�7��y�� 1A▟���]��q�C�CL�@��h8I)�����(.]cqCM��dM-� ���ֱsA
`a�Ų��~
�O�F6�4ș�o���!�c3O9v%H f̠�eK��$#d/@����$~w�FY��c�$ٝ�Z�'	t�,�#0ډM�=7�|/����z�*�!'��I;����,�L��ы��[q����yKj�p4'j�߇�FUxQ�. �U����#��DM2����[+�2����6��o%���11q��XɸLH��j�C�	�����Vj$�F�|���	� ˉ�C�j`�%���s�P����E+�� ����#��ƌye�ۮ� 7��}��p�V��U[V@�^i��ȢM{�v#����)�D�NȹO�H�g���?�K0Uݧ��MR�u�x�������;�Tl��U�!�ا�F�lCeZw�����^�?�ˈ;z�.�N�~��4���j��)`AN�uw�=�u$���/�`�����vt�zS�	ZN&݈C��Ic�`�FS�؂qRD�}�J�L��1S{���q��0I��UxmvfOUz�p���h����GQ��-��7�)��!"y�tG��{��L:����ZR�,�?��ڥ���ޅ������"�]Wv/ƒ�"�Dݛ]D� �?E��V�"@�L��Q��R�d�m�X�@��m��y^4��F�-1���S����7�o�`}��x���A�B��EE�S��&]C�dC ����[*ذ<���t����CR���]T�s��?�j�&`pg��ӊ6�T?���B��]�oG�rA��D�ra�������%��:Ǆ�~�#F�g�����+���m��_�T� (�E��}�¤C&���[q=�3���珥�	e,��/���w��6�������j#�� 0'���.�k�q�xA˩1��$(���(�|��<��/�AaIg{���i�vX�9�)al�9i�\�Wg�p���2�����0k��2mLm�{��g�08F����+{&-�t�"�gmg��$1��c�}h�j�oK�H���_}��a�:�i��\�Wp ��:�����4	��_C����}�fk��:���g���k�z
p��8M�e7~NJJ<�,3���+T�;��ל�
v�P�&m�^��j�4{��ip�P��*JT4�f����@�1��/`�!�U��\���"Y--�� �˲���T��%���D�� #�!"$m��v;�p����~gv�M��b4��f��\E��o�P���٥1�RҪ@	��D�_��-T�Qz8V�Y� �8y�A~��}��Qh�إa��M������2��07����L���)����2��O9�s��S�la��t���ѬrNOk�FG����r�g��R�B�!*�� peJ���@�P��PI���K�pҎn.W)�loǵ�)t��nQ�*�����PF���d9����8�fʣ}�<�91�6��Q��	/.B�s�ꞅ�9�rv�2��jУ2�8��ZLG����yq�B��M�Kzp�A��б�S��ʟm=!k\S>	�c�T��"j�V�:rrM}�irg���5�s^��g�m�K�!��b�'^��Y����0?�9�r��l�r��Ճ�.�WE���2�br	e�����S+-�������}��	�㳓�<�ˣ�TOr�(Zt쇤�����3��.�5z�Hd٣5����_�AZ���ۉb�Î�[��:�B��oaW��!�ZK�����*���vo�T}�k��5*���!��W9�A�G�,�_��B�m#ș�G�����N��gBl~5���+_�}..N�
8=,�-���&)C?E+�U�e)>��hD�G��y}l<���E��F�I�;uL�d�(�ou�N��Z���h��Q5p�"�(q[�=%������b�&�NT4�$S�7YL�N�&�1�PA���?��������U�w�!5�J:;�S�r�h�}]V�0�q�ɢ�VQ@$����#+J�z�eh%�"G��p���	&�=|ۉa�����^*.��������H��v��SI[�Q�0u��yOy�ywL�-���EU�@)��̕�<�����k<�,Bܥҗ�o��y�B��b9)<�u����H��Ut��ӱw�����c���7)�r��,�j�@-^=S��9�bW,��Wf�4��Iu��M�7��(5lte�}+,(d���2�m��k�bW�ELhb'�ܦ��X�b�����QDƛ�A�lj��[����z!�s&�&`�r5(�:i������#�c-f[n���Y��cA��t5!j�db��rƺ����5�By������{~) .(%�W%s��_��6K��q��Y����� �븰�7�I��֋u��PE(ws��Y�Y�#�����~�(\��1�	��2vT�Re坑��(���s5-
"���f)q�'���a�Z���Pm�s�*9�����q�ǂ<Mg�j���%�/�0����4���8uE� P�.�F&bfxx���;	C�����;��?Bٰg�~.�D8���Ǫ�E)KT�q�}�S�y�
ms�O�I?Fm=��(���ny� ŧ2 ���;�3�ܭ拪�]��<5�]8�[�Z�ˁ�-�=��#�H"�5@�M��&5R�Wo�%M�%f[*���u#��Y��-�G!����X_A���AəAD1�J�=w�q��3�K��o��یJz%�ԗэ�W���j�-�v���cŔR��������Fq���{N�Kk�l�������lȿ_t��bǌ�we*��ݻcd ���,�LN��)K�ZN�S;��N��=|����zj|�ρ��@ &�j^c�[�ňsC��CND�Ńj �������˺���@��_��i*B��]S�/�P(�^e�%	�ƙ��L�}j�������N�K�ׇ2��H0a�ON��/�{��1�z1/���Qf>d�YA��������hf���lȖh?�2b��Qws��_��>!��o�_6���Қ�ks�}kc/�<A��f��"�E)��t��O�Y	g��B�u��Pa�(�����mq4��j��9�*s��;�zM{�c�S#���4A�@t����w�,���Ou$7�v��3����c��e��1�n�X�.��߸���D���� �5����u�:�DјR���:ͷ4]�w�x�I.�x��l�����=��h�5���
!筠C~.��<z_��PD'��Z<Qh������
��8��;�H
!�t/�2��Y��I�� ��qA��[�x����j����DI&ؕ�����y�=eB`㦋v�=��8��(8�8Bg>�v�E��<Q��(')X�h�i��B��P(���*͠���K�L���՜ �q0փ7��YR7"ʥ4�k����v�&gNV�zy,�b�	A8��t�'��rF0�}�7��T?���'+w>�~�s��3�K��/E�R�!�;�	^�Xo��*=e�������3p�M��w8�HR`�DR�ӒX���c,�1Ŏ%3(x���O���q�oR�V}m�+�����|�>�`A�
^�y���y]o:�F�k#4�UK�X[�"uU�S�D���̶�){��> �����oy��bw�=��;?-���ޭ2$����u=`����}���Jo���gFķ�;�
���4x��e�U2*�$��~!�_1�UPV5`�շ����{���z��Ċ׫�!���^Y5g����2Zjn}��,���+��9����U	4��B%�T�;�(����O�PJf��y~ҩ�.p���V�)Ѽ����<��M�4\B㧐l+���(Ic\����,6А����tk��1���c@���`����/U>�,��:1���I �j��N��1(�W�3�9^��y�h�`S��J�zo�^z5��I�n�