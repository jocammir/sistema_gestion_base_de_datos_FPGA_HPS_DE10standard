��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�s^W���0A<��׶{�;Y	:0ơ��4D�K�6��=�j@8��s]9r��I�H~F|�x�U����M��Ct��tpT�v@��bZ�VE��TF[S�8��Lpǫʫ]� ��k����m#R��A�^7dn�����@lhS+#n�V$�j�z�.R�Y<O��� ����o}	|e�	�L��^	�T�v�+��IV=�����/"��1���띆� ���Q�)x\�������@��Ӭ�Baw��T�>���LCa�Z(\ҥ$�gG���x��>]�~D\Yl|<eሎHcn�ݸ�i�����D���id.#�jWkG����1�	V3����3�����h���|�A���o:'5N�D���R�9�\�E�@��~ (t�x9�y@9e#�W����̅��r|�o '��9t���I���;�6Hi�|����B�At�˛��'�O�/�G��}�s���x=���͈`�k֞|Y�Q����ql������G�<�He��ŏ'	I��M��[&���n���щ�h��Hj�8JatS�R�.�a�Խ�2-�&َ��i\�x-��*r>p9tq�{-�	2�H�4p"\F�"�{b�&5��n����=�-�����į� O�~4H3��@��� �%x�����>�v����� r�[5�22��}�p�#�u�J_{\U�A����֣~��K�k��N+6��%=Sfl����,�g�	Ų ���٨M�}6M�_ ��a�3�����r�h4{oۂ���K���?��硨��1@ƾ��m�����7NʏAt+�Fiܺ��A�)ai�[�y���]q�����$�*KX��ˋN�6j9ZP���˒����\\'"��gR�8�46>�^�)���I��f2�<s��t(-z>?���S���*݊�ˊgz��P��ٖ�:�Gm����@i�bXȣ��J�GzgMI����"�vmɈ�[ڙ�Ǐ���E�IE�c�z6?��GU�t;��WO%}U���։��*�i�Q$c������&X��t��͕�z�Y��B��M��)q� �!�s�Z���_�����������b؎F!�!V���,�4Τ��o���m�Hԙy��l�5�:ء#��B2]����!�O�����G=�|T8��V��x�O�f��)1��d&��~����3�F���먂2�ĥ�>LX�S����I�j��]�k�-6��gt���#����74�'~1�{�����BB!�{�3�8��,�\�u��x3�5m�6�w�t�|e�h̼�F;�PH��+}$Q�m`����r�B���ײĬ�à�x�i��R+�������Z��TO� ���[7��e�-��s3�
=:c���W��l���#��$L�s/4��+�f����������Pݺ�C�)�\h����'���SV����S�:�0E�Hؿ���_�"��V�`I�w7l4�v�;푍��"%����睼���6�6`�ai�k&S�_�>�1�'���,1uR_�ք={z�
���uL��X\(zeu[oz�|�Z�2�� �&<B�X�o�G2�{�=ز��ٴW>�b�v���p�w��!����Z|���2��3dR��As��S�v�(�������[�P[�ƵW���T!O��.��0������[�r�|���b�� �b��%%�3ځ��1}��q=�"\�J<E-�mi����^��y#?XR�a��T�=d�5���TGJaYMtv�t.1"�n\a!O�2D T����;�d�[*ML��؀-�&P�k�Q��������O��W��d��~]�Đޡ��m[x:9��f��]G��iB�LdӶc�>t-D3��f�8q��	�-ۨ��VMw�pB��T�t$�Ei��f#�;bO���#')�� L��X ��"h��5WoI�8=��7]����އN"�E���#����C�/�[I^�H��_:���^Y���+�J�4JR��0�|�[@@�t8�
��j=#D"@�V ��<��=s�U�ł�љ���9q���uG:���08�+�铔u��o%�H	8P_rр%�u+}�nE��v���8F27&.�8� ���迻��ͅ�Q{A��kTԄ�,ި\K0�;�x�
l�A�
�����9B�%.�v�5�}���E}�"�d�"��s��3���mA�x��RfnG�1w��E�#����!N�#��qֱ���R&�
����Y�3p�"eFf�/�ZN6�|}�j_�7?�$ߝ�A�Z�����t�V�p��䲓)�0���ܡ�l;��k8� Uۮ/��n��\�HP
�Y?\��$��"�e{rK�S��֊�TK�+��v�߅�m�md�Z�`�G�,�/J��g%~�|E�yK65"9݃��J��l�,ɣ��1p����}#��E+��g �e+X�NLћm�t�o��0���íZ{���N��*u^���Hܾq���x>�Jˀ����^�*��-}\;���O9�-�Н���2��	h)���U���#�NѨ~Y{5^u�p�ɤB�-�܊�?�p��Q^�GdQ$j�����Gp��t�(�z�G�}�eKS�' R��f�1���j�{'�l�%�S��W}�p4�)�0oJ��D�ݦJ(�I�}�2M��H�e���#�s���r·��<�y.�[f�G�	������ wb�����:��P�B�'&���Q��~X�T'tZ�����##�<e��u�o���&��qҍD*��fEE�͋!�!��O� ?c�`��g��8{mE#�Q�^�Fi��|S͇����p�Χ��&�r�W̪��(�{�&� �DIQ� АD7���AK��T�\��hi���@R�����f+�,eIM�{����,���.hb"�`|:-P����O�.�n���c��- �F�0���BW��K�d��\W&�]���	I��i$c0�D��E�oQ����25�k�l_�bB����?c��m���-�9%�և�1��b�WFN����7�(u��#���3�M�T�qU�3�#�p��<��u���p�^�Q�����'��b4�x�x�~\�P��F]mnF�ķ�0�s݅�_�����]¾��J�t=D��ֽ\m?���7�Νm�П�6�C��U_:������܂�hvR����m/Ki�_TU��!v,R ��J_0�r�>�����l5+v��ݳ�t $��_���'�*�T��<-��ߥ�$�������<��9VfV�;k�~�J�U�G.�2W+�FY>�� F�|d�`�M7�4�B�G��5hԻ��@��j���Fr��Y\��>���9�� l�O����1�����m@��	H�eZN�x���x;Z���O�
��s�2X�~]S*�6S-&8xV�)I.��֕�m����`^�*��<�D�yT&+��-�
h(Ҹ��CD��g�d��c	Ҙ�ٚ��������G_����O	���]��D�6�'��*_o�$��f/��#��*R��t6����C��������k�B�l�F�U���LcxI�L+\�۷�����w�惤Ш~�����=Ew3<�qy�X�ya�얏$����(�R���Q�gd�>Do�<�/Y��PNzTNNPw�U�����z����[�IS/�i�����EE�q1:��f~z.���z�9Ρ������a����r���˶2OI4zd���|�{iQHi#�#�1fx���q$���m3�x���L�[�*�er��H�s?��=Q'���!p��Fw�����q�U)>�ʖGK9r-v3��"����bSb�;��X�C�Ĉ5��Z�O���U�5d�m����|A��1Q�GF���!V`B��B�z�R|��B"��0%�*~S��&�yk��14�l���PPŞ��{ӫ�7T��?�c��k�������촕 c�*�*�R��T�0���lV�R#s�ݹ~�Y?�a����D���s�d���A��\�~E�L�;Mq��f睮|�x<�6�Ū�����f��!����ពJQb�S�ˁ1(��V�1��ɖ�d�H����1���Z<iLϞ+����_t��/�o��Ul���P�� IXI��j\�Pr����O�9#bK~��Bk_�����ãq'٩�O:�@��,37-Gb.�Վ�]}�2SH}��M���ѭ���μ-Ϣ-���^S-��%'��
�k�䝗k����8�a��s�1Yi�����聿�x5�D-��sw�Ş��^9CN�"�K�����K���u�i˧���1��M���O�[�������<�g�E^���,��)�Δ�[����{g�S�D�[:�r!��р�j9��[�z��Hp83��(>��ˡ���э����S
.g����X3S��k�,���Ie��$?�o �&��E	����d����ў'N�[�t��h�v�xsU��9%+B�T�?����qD�tt�����i4�W$�(�No�(T�l�D]gbK;R����K�3Y�g�4؉!Mڮ,���i6��Lfw�%�p?!X(k���οz�[)��Y֍�K�B�&��=�W�n��������{+[*4�l��Q��	wD�)��$��P���/ՍO�W?�YR�����3<����qH�!����#��������z8��k���؝'s�MS��Ր]���XS�"�U�9a���V����O�؃L󭧗e�Xh�34���}&Q4���$����j��������98|�ar�{
j�~�:q��d�Юb|q*�j]	�it������N�@.XCq�"��m@nW�y��͟V�q�Z%F������'`P��C��d:@(�JQ���^a��U�l�O_���)�o�T���f���1����\Ο䐺K胖��Q�%�����Ibc�qn�|L�I�)u���Cx���2�1$�4,���b�D������\%ν�1�itgi"͖�M3�
Kċ�p>�8�@�vUz��#� ,���+}�S���FY;\�B����=��'fv\ߎ
���a��JEN�[=B ��+�_�4^��-�{3�3 �����p���i�J�П��SU�I�d��qB�~��irJ&7�{c�=b�|2���1A	�����F��f�b��TK��y�Nr��Y���Ed�8.E�E���c�r'k�]��2W9�%5����}	H���ބ�%��@6�AO ܟ�۟���{EIO�7)�E���Ҙx�rU�m
8���M ������[��<n/9Lma2R�w��v��M?r�5�|x�I�<1O�;۞���*^��*Ȅ�"� �5�Un�K?���ƳD��MV��W�NE�QI�^y
�����_�J�--Ri+��u��K֤��X����������BT	8�t4�^�DD�̠�s5��]j����}��m=�<�O��!��R��e6�UP mp.��DX���SjW?n�<ZB��s�
W� ,޼zt d����!�1�r���`j$ˢ���p+1@M������t����<N�Xy�ToX�(dڣ��[	����f���x\��ؙ��>0�����s���P J�$��不���
�%3�5�����W@�m�3� e9bp~�F��`k�L��ɆhX�	��^��9�Ч?�ڱ��M�r��Vi}y�N]A4/�#�	
d:�`�@?>=�zl?Y��5�Ϟs?��&���)�a��$�˜�x,�A�j,"��t~/K�0eH��� rv�)���Z�[��44]�m�������{ޫ�`Rѥ��"��qcS�ǰ�`�iN�u�T~qx3��c�lvF��QW��X�v�(������W]�罪�1�G'(��\2��z�TD��^wD�ܤ��5��=��o^������H����L��[漽P�(�%�gUdQ�-�u$�^b9ħ�]"f����bp�
\u�#��lW'i�܅o� ���pd��%qm�T�o��)���`�!��B��LL�<�(�L
�3�~?�	�����G��e%��P��V�����~�Ռrү��g��YC��OIAo�4ð�&�t�y�n@�y:S��4�2r,���Q��S���dm�T�Nq��_�K<���Hz��/�-��yq�v�ݙ��EƵc�u��>4�	;�0�Pn�m2C���4f�PLbj8��kY��dT�B�t�N6�:��+�zN6�29���������'�C|)ƚ��Y �v��׻d	�m��@��{n�G�)�����mg�1��_�Ȱ�)��7ȞĖ_�!Z���wb�SB�����J=Qd�x�7���<!���fF'�T�l�/��r�<W���I�g��g�0�q��U���Q��'A���Z��\U�E�ziX2j��	�:��OQ7[Rt{|��>I��9lW��\j��[�r5�����G:��i@~"�k�[tڦ�?�m�`X7���a�����χv5�Q6���/��pw��x��5EÃ�l�2|X�yH�d����W�\S������>Y��\�}�Γ�eM�_;���;�~�O\���=P��ڛ�Q�V˽�*���\	���(<�{��c^�(\�K'��p{�W;���]7�]ܺgB��ٻ�^=h�/�-�������ӆ������hڙk�L�.$@�ꝉ��>nh}��mI�%�#W�$ã����`hb�`)��YCRГ��U�AۚY;���c���^��A�'��H�X(RѤ�ѳ-_.��󕇽���zH�\����NE�&��G��Of�Empʉ0\r���	X�_%�m����w���b\��p1�ř%<�K��1���1��H���d��[����E����z\2+�S���/U��s�á�\)
�ّ�w�-9�x�\��1KTBr�-��D���g��~�X^x�G�
��5�f��`�y�h�p���#�P�V9Б����"�m�h~��]�s2Mx�(�7xM6]#S�N�j�+q �(�a�Q��|��?g%�~k	�B�e�O���ʡ�S6���ʲҭ�w���!�n�\u�G�� ŗ{h�<��5�+ܖ��Է�)X�:���G��_����V����CPL�.�o�����Ñ�\�~���P���dx-E�E��	X��،�F�H��CP=Gp��5�Y��?&4?�P�%�{?�C�И}XL���?���5���i��B����?pw�0��u��ט����E}���3�N�>z8�ď���uȎ5u�l��M[��wp�>��w!tmu]ihQ��"�����Ο4��-�lJ�fڰƂ�<#�$JA�q��0_�j�[M*�v^Q�I��j�~�a�E�E)��j�������rE��x�D���8"^NKf�Im��a�Ol�?�y�\�s#mZ7�#|ֻ�i&�#�9�����T�J-�u�-DY2h��L�&-@W�ꡐ�3B���/�,3���*{�<Ц@�[ ��aCC �_���q
O�{w�5��10����:��������b��$T�����5|S���+�<��C$�-M��Z���R=�N_UU���@�r��B����*�3h�b�i���N#6�P���ٽ�mOb���]`~�x]�ӯK5�z��[�����e��/ � +CI�Q�p���3�������V1A��x��J�'�\�<r�wS��@+�H�$�l��/_�k���)3ι'�q� (,�D'��^m��� q �3v�h8i:�d">�vYgȼ��!�w�E{z����v7uw�O���B�qcjq�k!���R.$��_�`9��t��\B��B��2qyv]�jf�$d>J�--}v��!���,��R%�5�g��Oϖp6�y&��!��i���N�-�K����E^Η=���Mtg��!삖����%����,JR� :�_��]�~W��IiH�a�д
��(�[z}��;V�㻳|�C�խ�SF�VM�[����lݙvG�,�"�l��լ+����v�@1z�,l~�s�G2J|F�M�G��tA�D:+��7M�1�yL��f�S"�,��T�Z�)�x�ە��;���> �����<����c/59��""͚8؎M�=�^��_�F��H��M��G�(�99��)(>�?LV`7���1��[+᪻��T;`�U�k'=�bݮ3ɩ���8�43\P�B-;��s��v��:K���cDk�[V�`���ܩ�O7�-E�V�l+R,_�k�+�wT�r63G���40��JX�BrnK�A����
�/��o�>����k,`C3�W������l�|˞���A��P�;o����e���[����%��^�F�r����w��F�'�y�BP���C�e��3Z���7�1O�Y��6�U�����f�^ӗ[�,b�1�eEC\����d�69Yx&O�K�}��%ܵ62�����Ð��a8����}�򛎠����U?������@�QG3I|q���g�x$��I$˯x����^	���R�uECT�u�?��$��/��J�8r�? (m���&��φҡc��>4�\I��@����~E���1��S�`[�JJ��	�N����O�Fq��g�~y}��L�|OtA�;;a�Sj�qa�HOrxD������j]��>���0��%��6�6�}l�oۉZ����C'�~�t7�|�h)��;�'e�A�����$��\ JY���5� �����ݐ�*��n�e#�d1Zb4f�>�l�$������{��0Y��9:-�q%�pX�k���:��
$����>#յGO�c����-�d�C��&��_�E�����e�~�C�_��5:PxU	h����E��Z-�� ��Ύ+#a�T��:h���ߖ:��w�V������l��o]�����NƦ�L��o�S�dE"�E��P�F����Nƨ���ێ+�B��p�6����\��T�e�+KXe�p��N�@�.LnC2ɹ����W%�Tm4X�dگ��ϱJSw��9<A��~N�0�8\��!q����Q�dW�U���\�wc�$3�t������c"p�Y����n؜R��ð!���\X����#@��a��\��R���4Y�d��Q���b<g��V�G�X���3�d�Ɲ/�|��
�O^�so�&���4����:sL����J�&�i[�e+����:lIl�j�v?aD&2�R�#��؀&sZ�
%&�CV���DKk�J��j�_x�������vbӐ�S���ܝ5����1�fZ���?'ߺ�K=�<��M���Ǽ�\p޺ �y�_�c��)V�j�[	�����#�C�KR��t��^:��'{�hRkQsƮ ^z�[��"�����i�j�͕�νC$�E/�9!�*�4Fo�*Lu~�������M2zl%'8����G��G2�>�Q����?�]�F|~�`�O:���ނ���b�ocV��]k��k��h���HH�ƹ�����Q��XƇ�HG.���*�=�5����Ph>MB�@��ٔpl2?�#LI ΢~�9D��a�_)��M�N�?�a���ko�0��Y�u�>�?љ�E����s�LE�@��^���zϩflX�&��(`VN�I6���
�~�\Y�֍��I���Z��+>�f�,�
�'"��V�e5|u���H������Ȭ/@G= -��"ܜ���c��L]��YD��|G �J��x8D��`h A����|�w�H%�)j�T"$��������r�����x��ـ���g�y�t�2
��m�{sS��,�d�@��`����) ������5:�a�&�bKZ�2��� �*�1����?�$~Z��B6��t���TIm�M���&����$������e��Ĝ` ��K�o�b-���9>�z6�QX&�Zuc�{���n�i��r�������AY�m��ȁ�� Us*��J��VFT�ET,��9�_ ��^����fSO��\+����}�+"���
&qڲ��ǀ����.�g���#z����g��(�Vٱ��|C�WA)$�l�¯N�zSC��������A�Ӹ����J��^���Y�ſ�z���v�Ŷ�pM�N�S-��#Vi��"ys#R�u��t'Ж���-�ԧ�!b��#�|�V���Ņ�,���ؙ���,h����M�1�C⯬
_uf0�"�n���Udǣ��:�F5/�=���q/޼����o2@,��'x)Ģ�|V�p�Izc۹Tp��I�Ce��wz0J�6�<E)�mH
k�T�	P�����Aq�z�gP�S�;�)����]G5�I����q�}L�r^��"�fѯ2s���W���ӏ4M����sM�;7}
�x�MRy�A"��U��/}�g-��y�V�b�a��q���<N�X�Z�'�h$��*+�"��np�	����4�fzB:�֢�cۍ�Jyw���c���Eh���	>��������wwN�z�ȸ��-ځo���������}�Y8��$��ؿ�?-�f5��+i�͙v��Vc����G��p�0�n���
^�O�W�~9h!p/ԕ=L�#^�U%{gxA2�1+B�������A2	�����R��:�eM}P̺�٦�������2�S�68��6�>��*!�j���p��S�C���k#��9�D��/���%�㪇�d�8��O`Q氰\+���Gn>�'���[�[P�S����U�ڙ)��}�Ⱦ���p=ܚ�/s�T��!JF���M����#.w֕��A��	��s1���u$�@!S��py�<eew� \zs5^'#�����������qG����\w࿠XpA/>&򠪂�cw?Ǉ�j�+�W~�� ��!PlE8;�ǩ80o��U/�i���)!��>	kzA�Q���3s��L�x�=ZX�f���] }�3@�ײ���-�H����m��+.*�Ic��K䣩���=M�Ө�0:�ϡ�/|R��+Ȍ伹]?�j��mG��U���,c�SQy@'�(��T�����Qw�i�4�
X.�Զ/F�m�s8B��gT��Y��B:���(�naw�[�I��#����H�c�j\�����]�͕�Y�/X?�ܽ��B�+�x?P)L�GH�	v�LJ��X��P(�~�o��L����k.�*��5�]��h�(âC���T0�y�㏷8�l.�T-�v׫��=$�� k�����e-�p�g���d����-4��5b	'��� �x����p����qS׆��D�0����H�X��	�?ӝZ�m����еU�m�y����"�ӆU��g5��L��=�Ի�A��ͽ�N.�.�cLвT����`j�F��.^�j�_�?\�Y�f;H�v�s�K�ʓ}�+��R��35D��I� �,<T��[��������L��|��w�H#9��:���U����P���ۥb�����I`��y:%2� �X��V���&�Q���G��A�lbfW��	=�Rr�����z3&C����T�T�Zf+�n����~S4�:�L��)�8����/%��N�s��0�-M�=�(������9���jV�rx���|��s��\D��jp%`�?��<�������ZB^�Fx�V/��4Xæ�g�(i�w_�s��Q�nx�ܼ�#�R�P	J�hji��!*L�����mE1g��	c���S���Oޤ(�C3�Ix��h;18@��-����:���vU*7c��-������u;䶳{��&fr�l�@3��74�#��!#[�g��4c����mD{���A|��ǍG#�
�;F�9f(=�Pm�mv7��o��-�y6y~L�Q�s'�������dQ5�$-�[�9���Ҩ�SO��)/����E3�t,AB�!�0�2����'[H)��_)�INw���hD[^�U^��>�
hj#�7�.���Bs�����Ó�݀�/D���~5Wd�L�a-b�oZ�-ܥ���]���B,4���*|"�d�Dnj �f�^!vk�_ �~L�|>�����Mڸ��,�I��V�G0�S���K��K���Ǐڊ#�2X��k���+P�����}�����6���֤���Q�X&r�p4Z����=�2���Q��r��>�d,a��ᘮ��Q��zCL�v��%�r[zu�gpPn�4�<��;·f�3�阦���'F��iAʳ��?[��ȁ��%�(1��+�\�t>u���p7O��^���;.�]뻌�?땵(�o'W�>$\N���E`,���B��b��b_P,b�LQ���D�4�m���]z�M�K"�9�qiJ��I+���})��4�/�ޑ�(��Ql$�5�((@Z����ٿ�3Q<��TԚ\.<����J�T
}�e���͜(b�_T	�=� ��ӥf�j^�R��?��\%' L��8T��à,�'oaYr�W~�+��-+q�:������;ih�~�qtD{đh�:�WO.���@��5�������܉�L�st�{�(�#�)�
Os�;��Ćz��+1�x�"~~���Ah-�6@瞊�� ��Mj�] S7��+���h����å�Ť]��Sl!,,���Cy��Xڿ#�W�/2�	Y��=�a�����v�v{���AUH��o��b!�#Z��,-q)���|��UM@NU������u4\B.ct<�����Kj�\�Q�P���_+��{������IP�C�N��Vw	�H�Չ����~ I��ڹ���C��p�3���X@w�y�6o��3xӃa�V���Kͭ>N�ý�.X���x
X��ծ9�Q�h�95�<�VN��r������N~�4U
���+�&�f�����J����7*
�Jh����_�m*9SE����^�� �2�-<�\Y��ٜ$9$}�*h��]Z_ku��3Z��X�^/Z�����wx>�e�6�W.��)�,Hw�-|Qn��{��]V����,���ەfC���,�;z%}�1ea2��f���b�����U"U"rK̓U",Q�h�	fg�Y�L�g����b�a���ȒB]�ԅ�$��k�|����}��_SV?H|�ls.���+?�m�{wC�'`aR��9�ϫ�ț����,��m�۸\2D��u���r+4oa.����fn��Q���� \��a��#�Х�:��5�;�	��	w�r���gE5*�o����ä�	���`-��
[��䈿UQ�|hA��K��n�g��N�_��X#J�He����Ã;��=_�C_�| �1�|趓M&�qMY������������I`�;74��Jb�)Zz��NF嶯	�E��F6 1ɖWS��w߽[�th4���<���a��<�#�5
�'V��렫�ǽ��fr�,7�M�H�������$�����G�1����ߜ��ul�4	�NX`�]Q$�'�9����&�~�)ʕ���"6��`��qY��!�%21
^������n����ۮ��-�<TEr�3�m�bu2��b��ALIZ;������A ��pWU(�n�.	[/���Y���(�����X��l�nT_29ѠSÚ_jy�Oިq���jFhv��E�=z\8HU�����/�ao\�i���<s�'���-l4yE�i���Z�sH�E�y��b��Sf��T�n��#	5ۣ�弁�+-Cdy]���_1V��&E4r���KovBF������s�<��a�C�yE����'-�A�I.�kWۖ��m6�[�|j'��5\��&�6���4������	��5;��]�&;�H���bI?��e<$#ڀiv�U�$�N�r��aC�I�he��s��m�J�����hpc�7r����!��S�wN��y�ʟ����w6eP��l���f�Vp���r��#N]Ao-S�5��jQ-d��0�Y�P����_:�hc6F�ubJo(U�|�pv�^&4��G,��'ZU�����uE�����2&Ź�+ۍ�v�i��o��v�k��2*>ku���_eQy����p�眳�\�Ɛ�_f�[�S蝡�͂�vC�{�}L<jJn��^9���ąoJ�:|^�t0�KCr��e���3)w6l
�/*����ު_\o,��|E�,̳���_�6 ;�\��I�!
�}[�C5  ��,4�<�C�#�i�B�Ȗ>���6m8��\I;0��� OC61��P��I�~ڞ�]7��A!�	�p��98Rə��>]7����������3����������*�U�};� jY�G�N$�_%u��]B�[�b���/�ͯ��'YC�:P�ww�ܳ��ldm� x;*��9.~�a�gp��gY�w[�i@�8\�l ����/~�a�FψU�pB8x:0Wޔ��%�r����S�=a$h��:��R?��T�x�K;8+�T����{���֘��\�*�����w�z�R����W0��T]�,fR�z�x���(��0�Vg�N%��XKwQ�	�o�d���f��	�)R�Lm��� ��!j*ڛН���)o������T�z���De%��t0u���ɑ`�6���8�\��O�̚9[xKq߷ C�	�,w�<��� P�����pNSx�l>���HaLP����=Q��v�&����$��k��<.�w��R�	�x^2ٓ���r�ذ��"�N�G)>�^'��Q	߯�є���.
��9gT��745L\[�PwW���Y��G���i-,�	�!��K�8�j��(��� ����wͷ���Ͳ��X�6��ۦWn�d� ��CH"�O;J*��"�y-~�K���$@4��k��Ck�!�h��FԎh± ;��a_�\~��`;�ي>���n�'P�K��ʴ���	#sFm�V�x�ό�,�DK\�uu���3�Va�0l�n2&FbEa����%ѵw�!f�:9�d~�� 0Gӓ��E8�Ν��͞���v� Se�bG	j�	e��h��	
ޢz�H��i�^U/L/[g����"&���F��d��A�_��-�=�1YBL��@|��h��.�g�6syA	�jo~��A15XǨWm