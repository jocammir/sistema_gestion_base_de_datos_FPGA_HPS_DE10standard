��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0����_���3e���ӌ,nD��	� ���Cgv��s�żEN#�f�Q�l���G��ŷ�a�]u&�C�m�9�*KF�Q���@e�����c�V��ݙ�2�m	��h��|k_��E5���ꂙN�ˎ�Ђ��r� �5�DpIC*Br�ʮ⳾̝m��0�5����\�F1�O�H6���V�kO��k��S位��\�C3u}x���`���D�3�bU�	u^o�N�[U֓�<ЎUO��\KǊ��@��H}��ݩ_�l�6f�E�R1���̽������� ]Q⾩�]ɱ8����_�uk�כ}��r`h(�# #����o�:�;�e�����_�Q�u��=�]6������ ���.��=��'�,��f��m�o��%��������v�cb���WZr(�� �V��'Z��ȅ��%�Z2/�`BW*��Zs3����j�M ���S�����N+&����.ς�m����n�P ��'�I{�~@)��7�3(�;fP$H���"��4���M����^>:�Ʈ;�؃~�Q&d��ߜ($�j�O�_��b���ҭ�`��_kԟ�qĖ�7�ncr�5�5>������xU��~Eۤ�>�Q"��o�d !L��϶�$�s��&b�G�w�n)���EƷ�0w�K�iQWe�5�80�?'�������sz�\��d�
���;9v$^��������Cw��p�C�>�aӰ�;ʲ� z�ZܲsG�1ʞ�Bʬ���zo�}�QX������^"G��!%l�Or��Q�y�7�jk��(�>�ì������,�BH"H4��'�m;/g�s:�x���]����O�q���W���|�r�G<��Y:���דF����Id��NÈ�d�����!� <�͗d��>}ݢ�~	ذ����G�wHV1#�c	����-	���r�;!z�+]F;d�
��wN�7�53���s���%^j��q��X?@sJ���s`�B;�dǆ� ���İ�VE^��I��՚���y�l��@��p��ݮ=Rv.�����z�J��e�"~%������xz�^���*zq�s�ʟi��h�@C����+���v��"�e�m �����Y�OfaL�1�;����,��ڦ�\�a3\�k~�EVe���H 
��P��ʀ�n��[K���iY��� �GI�5�S�/�B��d�O��[��W�'Wk��cf���W�b@��~��f��Z0�D58�P\;��������H �۔����5�'-�\�m&;z��Q�|`i���b�`i��x^�;��=*gNF�6aQ��f!<K�쀔3���)���zw�ĭq���c�^��1��]i��~�4��ZJ5%�C�+�U��d��?K��Ң~�jΗ,�cm]�l��=Qn����z�r�.�����Mq�k{�VN��kgp�I��s���	<n��y�垀�
M��1";��vai��2��N�;/k�٭R��Xq�����wů5^���Uh��\ �vby�19��<��^�"��i��A���Jq�!��+[�����<(¹w����d`8m�X�-e uB}` �"0=|�'�fy#�xpd�9��\��Sg&��`�P�6�<e仞\��N����T&�LJ�=bl_W�b����?��Ob������%�d�2=����#�J꫓���C�)q4/�x)���T�e��<F}=�3��=fFxvDIu�&[1�J0��]Y��2I�E���@�,����E�����������|t1ظ�(1H���W�T�w�.��z ��|fC��P<<�G�c�&�.�l ����${���@��.2.W������O�Pl��E����N�&\�+|x�6|��B˶9�jn����%�;\��r��P�5ͅ��W��t4�
dj<J<cl��%#�Y�\���z5����;˨�n���$���F��r�)]j)���� �����$���9 f�
 T�(1��9M��Fy�)4�6��E�'��7 V�\	�"�P�W��b��O���	��D���h��y�`V�&�;.XR�2���v%Z����f��QMH���(��~�m���ۘ��N&p�=�ɽ�sb+�ӵ��+����Q�Ƅ@�V�[�R�be'�uP���П�r�36�'��3^��U���X%I@��u�������--��w9����PM_�(�y1�u�d��E��B c�s-���w��9�T��ÞIº8�C�s&N �lut�"a|�������+52�Rm�WT����:����>n��.bf�7��Poj��erK�~eP� ���^z?�N��jw�T��k;JG�5�@ ���I��I~}�~Ԏ߬ƃu���ecT.K����^⥿a���΃�1��շv�Du���V�a�]�l(%r�W����R�`�\K'��Y���HS^�Jg������?^I��OI��Kx$P4�cǭ��h��r�(���T\:)mˁà�yGm�M�\��
�é{�4:��b��Uפ\Tt�4��bh�����X��`�G�qT����O�2$�)9Yo���a5]ĲLM�����9-lp��f4��X޲���|$���߂�4쉎��������y�>���|����V|y������["mΊpo�VAc���K{@#���{3��1�M���Õ���l�����À3�����i�x�l�V�VF�o[�"�I�C6�-,�La��oD1�L%��K��yfx`�'�j�`�z[�1@Wi��6���~F���_8ݧ��zC�_5�.*P鑫<�X20��>��F�eD3{�T]t�����0�j�xA�[/�MZ�`H.��;v9+-g�f��Q^�wN�w�=fT�>�Fh�^$����p=�-���������<9z�<*]m�����.�S0%��oO`���{����"�Ծ��q��¢�dzs�n��xhO:���QHϺ	��-��(��v��<0Y�1,d��Z>P�YJ\[e-��f�A B��/��y�3�#��ma�F�P�C�
8�.�!&7I�����@�@aͲ�*�����dvjA<	I�o���Oq����7b\�	P��ĻpB��7�"4�(ş��<�m����_[��Ź�~�r�NɆқ�9<\��ͅ�n$e�����`��~1ٚ�ɉ�O��܃� �x�1~�g���8磚��6_���okᮮ���E�� �g��	S���t����k����	��-��PC^t@2�Rq6.Zv@eߴ��PGY�����BS&1C�7G���d���f�ɕM�R��]3_B��*�ND�l͖Ͱ��s[��w��W 	����G8�FJ���7E���usQ��jJ����Xu�RH�s'<�X��'�jle�#��PR����vN9�Z9�N�� X�"9�e((�g������Z���w�����v�߱��"�db���i�m.����p�	hO��~T
�'w���ľ�ͻ��AL���D�J��sH�R���濴��R���\�0t��dz;��O���>�)�hC�{��.�
��=���PK+��L�2�I�ȍ�w<��	�B.����O���L�-=�[�]��Fs[��*@!P����D�r+�@�|�)�R�rnAt�ŷ���t-eE1�f�3��Гv�IQ���{)�]r�!��Pg���dR[�Ś1X�,辭���v�|��מ|;8��v�K¢�@6�O�a���f����)ڋ���4���w�g�;��4���P ��e�[�"�r ��E����ע(���VnA}f+�&}��&*�X���qo�Ɍ�3}^�'��d�����.?ܓ?�W�%��>�����4w`hc�@<�`DO�G�aH����'�������t�A��K�/�X��UQ�1���T�S�&�eIT�	lDK�����54_m�54�{�(��QZy��, _ L����{HC�6BC�7�I�m^@�u	��S�d�={�#��"�{r�/�+7���1j�d�O�~�A��Wyu	�N��jK��{�yy�N�N��2a<)!$�syOo�v�j��`{���{܆'�����n�h�^�!����XkƜ��$�%7�b�����������ީL)������3.}�2�Ȯk�h��b���:���Cp�`�E-`��)�{�l��&���翃$f��lxJ����o���6 �u��o^2���<�8,�nus���D)���#
�9�܆D���vxm�Ӷ��O�����X��AV�zv����aPfjf�<����h&J�L�$�
�y�,��(�1��!��m�2��޻�q��P5_��+�����B>����/j=!Z�*g�(+����Җ�_��*�p�t����n�ގ-��}��׾T��UH+*sH���\q��4̶+� {�g�i�S�?�6Ŋ��Q��-rj�VQ�B�����k 
�K����lVĨ7]��h��x��ƙ��n|ߵCk+��Ns�uhf�,����)�{�ܬ�؏a�u�i&NTp9�8FK�7'��t��R_��;1�>ewaqjF80�>,5���������4���}_���K�Q���~��ѡ-^�T>=���-�o�>^G�NШ��ڌ����­a�B�5�����{��%կ�0����yJ�w��W������kxL2��rOK�0�/'h�v{���*/��i����&ݻ�f�r�x�pE�5�prq;�<dU�!���U�<	�h"qX���_�I�o���y;�ǡ�;q�~���	���WZ�d<H�n��:̮
~B��nr�,�0Mf��P��C��+9�7����
�=�4X��Hb�m���	N�	=z~Ŕ#�
T���
�p�E����Sz��$i ���2�i p�����k��!��|�nx�ĉ6r[�'�*N4��xu��A�E�A�
�����!�h
 ��(:EV4�~�`���B�9�sw)�d;�h������un>��2]W��ݱ�G��\N�� ����Ä� �y��@�;��f�#wjy�(#��r(o�	���o�h�3�fܓ����?^v�vCv��nT$o�O���˓  *u��=y���~�9��_
��!�	-(ly&��f�.C(�(|�/c��xh�{�v/�碂�����`�c�����	)t)m �'��j��������>s��u�t՜�?���Tawd&���StJ�ƃt����L�iҵ��I[�@� �:	��t�������:O�>S��2���v������2ѐ�?����Љܽ��?�}�ߙ����5_���&mk����6�6��gɀ�<�z��Jpl/.���A��VV�?&�s��ֲl��Ld:��z�啪������4�~���U���2���]�-�z	�͘�T�c�^M>�P��NW�����M��-�c2QV�w}�/=M����7v�m����]��w��&��"c罹������p�l�X�'>H/���Δ�\ƒ~�R�{kXZ��=�S�eitu̵�S`��K�HF"��^��� �.0UX�+�'*��r���ںA���F�\��}�a�GA(�e*�����}��'�'��-j�?�li���h�F5���JX�e��\��3��qL@�@'��E�s�<���0���O��O�V��n�a�����*͗�Zzu���5��f()Ε뤳I^@�V�V��L'̫/=�7N�?���`�OV�mP?���^�|f�I��3��hl3��,1� �TF@^��xd$�Gv�1��9�X������i�Y@���0�@�����β��圝��Pڣ�Q�*�����\ZK��{b����e7d����'�B�1O�Dv%�82����J���j	����4���<��,����"
��*G�+u4��"Sѱˬt���p&.�<���&t�-U"ڒ��f���B���M���<^&X��N*���´�G�V�X�nhA/�����JP0D��(E%��P|X����NۡE��J����j��|����!�N�F��aw�s	��y�&(g�d��$E�k��C�lڔB���~���GH�i��~0�"c"e���f�98�Te���Gr��X�I�go�7<16&�+z��@znL�a���BJ��ZѺ�;Ŝ�=w���S֏ޜ皳�p�t�և��������EY1�q�3~�
�x�k��)�j�;p݀��$)WK4�?o|�C��n>��jʵkKB�T�͊��6=�DI�M����$�pl�����â\Z��&���K��V��KŲ��
ňXNWye^����K��!�Q����w�$f��UL:R�������]5w\K������`zyvV%�����m�������A��UA�C���Fɸ�ߚM���z'��?�AG�<3Z�a��a{���^��:�:Mm���$������i����+�h�nz�M;z���`1��O�����o���s��.�ן��ny�-��x*�0,Za��C�I�L�T �٭��@`e�U��\�����,��ik��X"�11X����s䰘��U�PJ�������4�����dBS	K`��JM܅Ҏ�� Tŝɞ�07
�T���vs�����g��(����Z7��M���xRm�/�tc��)7�k�u�>PŪ��@��(�+�p@1�S�e�s�u��gL[R���*:q�iT�u�<J�?�c�y�쁿ʔ(��zњ)|��R���W���B�uI�t����륍9������1gDt�9~�֧��qǵhbU}_G"����l�U�	,�٘J&�M�~cI �9�/�L��Z�{�վ,~;�Q��l�������䛚����Z`�-��Z��?��W�J�+�dB�r�hg�}�˟k��450d3�/�O� Ye��_�$���������3�jޛ������b{�1���go�B
<���0G�G�[&�bߺ���>�a�=51�k��˳0&g��]�� "t��i���3M���BmW8_�A�AQ�L���q{�&W\]�2�3MJ�<#u��l�����ѕu2.��	�\-��V��ǚ�{��_���qg�ي�w�4���w� �����N��QJO�e���0��r�I��v�d0�4�JKm�X^�)��(]�5w��EHc{Si��2�����2���yo���� D�b�^��XTt�*�㠑�/!a`A	�f�8��`c�a}�g��ks�NlAO^2���t�Sq�����$����ݦp�j�!o=�����k�REITT^  �Oqg!�� N��_0�ĮV9\!ux����m�UA[��&9�o_ %�M]d���^��bv47�G)t��,PǮ7�#01��]�_��y�()]ɡ�0~}V����Dq���������xo��Hm�����~BPTm,��g�xt9Td���`��?�|7���MFO�-_0�A��b�����-h�U�޳�$V��^Uh����w�U\����zF���9��t/D�3��X	\;�J�]��@��~��a�(������fa�)��ףp�(
�f-��L�vЄ��W�>��	�'8Ӵ2�[/�Ҍ����8�Y��鸉���%7�!���n���ݥ1��5;���V�0��_�3�OW����RA@1�|L�8l:��2Σ�?�}����Lo�П�b�dv��<9�YQ�Ȍ)�cS�>�d�eH��QyXI��7J�����NW��7-���F���+�I8�qG-�Hϯb��6��KJ�p��1Fᑝ���=�8�	A��\��dICC�t���Ҙ�وL?�o���&c�{�.��W�������U\��������ͭ��T�(n�A�D��#�F���܉j�.�4� �A_�a��?<�_��<V�臭�g��0�ޮdV�Ii����`qT>�{	kB�-�����{xˆ��)�@���;=�oKG'Q)�`S��%�()Q��Oz#����C��:�q�t�X�Qq{��(~���ȧ!Sw���`e�C�¿��	)�R}�I��~�u�>�T�f3�YAߨn�7�����ћk�D��Ż�ۣ����"�G� �
���6V�v!�sj�N�r F�]c��o��+Dj����l:[N]�X�Q	y�`�i�Rs�Nr�Wn� �I9�+��Y{b������z$*�@
 '����VZ���@���X�����N�9�0
�n���MS�s��_��o����f��%��DϤV�H�����T���r���Z���R,�=��[�]�ΧP�hL�F��W
���ˁ �"��E�L0ӍMi/�#��>K?KsʣQG���n���o�*����_B�È:<�;Q:tK��Z����ʞ�(@ֿ��a���*�a
��)��F��~~�b"%������]�_%�И�DQG��E
�F���I�j}�-ͷ4��~�{�-h��</��&�U�K_��[��Fե fE ���L�!�+�\s�������D����ў�u<���)��,f`��+Z,��T��e>*�n7�.�;��g�}�N��G|\Xd7럖���)�ނ��>����d�����G��w�u-pa@|���J�@��<�1�N��� ��?���rp�Q��i��ӸP�Ο 0��~�?��7&Y����~a5ix�;��P2�XXg3]+y�~�(����|޾M_�����6Þ4�q���~�%������f�m.KLx�%����16�&zҮPO�7Hju@���y��9\�)
�Zn\�}#�of��g��dR���	���b�)3n>S��K������^vY�P�r1�j=}��(�=@�H�{V��l�ꤋB�� d�d��R%0(Ar����<�t'����ܺ��~��|.����&G�ͰW�(��"�N���x��T�庮M#������j͡�mc�+�<�[o��(�NVL|�p[���ǥ���+���M�f\%@�RV�y!�^���r�����]���	��_�#FX�T�a�7���F�J��� Aʨ��C`γ6��ݽ�hfU������5�j.ǻ�d��F�T��p^�k����3x$�IڢC	��TK݈�i
z��Y�%1�s��a��7K��q�Z%̴��m�I��&�,�|�88�%�]��vFܕ��;Z���[@x(�<�è�
��Gh�Ns��OBQ� J�r ��Y��2�I��#SM���r�� V_4�m'4����_����V�)�(L�����|��R���	��˜�2��1�(ߊAw��,m	