��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��ᕫ��H��gq�f}���+����c��0�7�*�y�HXH�+��Y�Ar�#�<�k���bu�-��.���O�;����b���7pE+�������v@��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T幭xX��8�hG��kr��'�n�IK�v3�[B���fP�e�q���7V�&����J��v�(� ��n^�ӄ�`� S��JK��W�|�	�bL�Ԡu�%��x��@:���Vì���t��d�Jr��%����9LZXY����Q؀���62Ƿ��Rx��mF�h�<�U�<?�]R����~1l&�T$��_�6ѴJ���{���kN�_���G@)+6�ԐN���'*>�c��J�2�
a�e}��%���A�\BU!���Lu��hp�%��Mۆ��T��h�mG}��_�����ep�����2��a&�ĸsK����ڴ�]CV���V�n�	��_
���S���U�c����.�s�^���T�B��ǒ	fjto>�v���6;����ċ��g����`��̀p��z���&�Cy&��^`tl9�_�<�T垘����Oc�Q�߾-�1�u/����H�[Ig9m���H��>M�F/L�0{��ܑ�G"2� E�1��N���k�_�#퓹��a$�΂&~�Ij�1���.}dt�AfAeT�4��*Jñ���e�q4��D�I�`�ϨΩ�:N�g�����u
,�^���o�rq �����h}��/���6�C���0�aw4d���n3Ranq5��S"�$tЫ�K��*�`��+Xc�ԫ�C�Ƽ"�0X�kP�N���"]B�<����f���I$���R*��e)ڋo��sj���8��.1^l�����e�=�F�щ(l�^���m΋���9Ĝ�!���8ﮪ�̋������X*nm�9��'}k{����2�߈� ���~K��:H������M�����>�ȋ��D��f�	�յT��=������{�`��	t��！��f@�y����K��?w"0���rՁ6��"�2�`�m�V�����$桧��w�5�Ł���2b��`��	(�U<D��+���8V*�K5\)_�ʑ!�p�����Y�,�o�ӯgۋ4�}���Jk�v�6C�&�k�#�_Â�n?�S�E�͊�UQ�z�j4^�Ǡ#pm�ԕKv ť5���f9�@�t�w���Cf�T�/(�Y��> g������)�S6tX��f�<�6َ�K�c���7�s.���#��A���!o�Ϥ�:�Z����U�����{��Q�~��qh���Kq�p���jR��Z�d���%���%]��T`PN�t	��^YBT6��DM2� $�b����iS�G'\k�7�c�z���)%Q!��������J�`������H̤Z�����B�#���J������]�:ĖGݱ.'S��J��95���{+�5��/�	�J�t��$㱦���*W�?��~
;h�z�)�dm-���3�h4�%�5j��v<��Ӟ�|TR5H�9K��!J���^�������x��v��Xr��B{z�)W\��T�Kv�eC�g�beM/�b#����f�)�B�P�V�)x���{6%���2��KI�9:֓�w)w����d���A�aS_.��^W��=�|��~���:� b¨��V}9q׳\�f3a5~>����'eNd|&8�~�QOQ� .A�]�L�Zd�W���� RMUX��4��P|��|������u�d���,��Tun�jh���T�C����b�l�U�N��!_Q'��,���Aӵb�Oym��'>ז�;�x����-��g����mEA�v�++P�-em�I�ȕd���F��64�xa�x hBc��a^I������>�X���-�}�'�o�pa���AM��1J�4������ �%Ɵfm�]2�]��j,�1.90��3[�&` /�����_����Gq��8��� �3��~��Jz�]c��*1��6k��z#�͔4��J�����.�"�O�חR�uF����!�^��M�~ᯮ�}��]���h���L�v�h�]��2��C]�2�;��EK(B|^�J�kt��_mPn��2��aKp֊��~G���V����k��
�(�|�/C��`��=K�̊�\w�:�%at�%cNSB�����%���}Z��>��{�(8)�+q_��&ę�pJA�,ǥ��L	�v�P7��S�����b��1
�e'}�lИ��>���m��^|; H����+H���?-��Q��'L?�y�o���]K�kL<�j�?����Hh\�zc�<�b6�&r��{�U�K'ZO������X��P_-;d��Z*|�����͞8>���x�<��x
���['R^�NI�TSu����4G{U9T�����	�O��=v_e��؟�ꔚ�
؁�.+p��b@>1ZF��;q�ߒ��
z�B�,�ỿ��p��S�b��;/@B���9oL�:�X��I��$�\�|ǰ�K��K�GoP���a��#��	����Pu}!5eb�[���ѻ������O��8"� e?����_�\�i�|e�%�qw?(dS�OYv,�#cǇ�h�� q�x늃|A<�-Hg6!ɜ,dk�j*��$������%6�@s	LD�ݯ*�2.\F(&}�����\5AzAk��D��N%��褰�����\�Y�D�)Wv�mT^cų��r��y$�^P���̢A��Őn&V�]�-Ǒ�FO�p3�1�vU��4�a��}��Lo!05��3�߉���bt�	���<<i6�� o������r,���׮y��K,z��q<u�7C���_d��@Ĕ|~z�H�{x�F�:���WQ�Qe���x�1li���\^W<��0�)m[(Yr+���;?��d�V��3��č��MR�]tC���;Z|F�.49;!ױ2<��.�7-wqƁ�ϱ������)�S&U�/����_�~b��������G��?|�]��G]�5�]�y����O��z��{��l�%��_�+[a _�oF����Z��7킣��/<�9����'�z�e��:��"�) �6��Y�0`?�-{!�l3��g��}:�x�H�ߢ�fq�d�g�_�`}�����~��jI��,{�y���;����qPA#�R�S9ؑ+��3�6P��G��L�I�EypɭB���
g��m��?9`�FC8���>�99d�>��ی�#ǳڝ�g��/�1
z�JA4��tx��!��ea'��kyJ�b[�ˎ�9o�Z�;�yB1���R�+�^�{u�ݹ�n�G�"F�*P���^�`�(�Ģ����� ș�oT�+k*3�[�^�D�%˘;(��N9&����Odܦi��(���c.��c�s����n#�4�%�۴�a�A~����ގ칒Gh 򇿔��5�ϵ;Z��W�q�Y����&���A@a�����@�g�@;�{	���C�P��� ��zAsn�a"07xf�Qb(�%��6}p����!0[��y_�9_j�`�;��w�,iRօ�(gHU��'	'�D��V�H~t���Yg����j�n�@�?{P�U��'L�m}r�c9ҿ��a������z\��t��>���u�����!� |�����eI���͈�I� �w����tb�1��6��&�|��p�2ryr�m�vyG3q�9u��s����c=�IӤ�龘JhU()a�vC&R�{�%��`p#?{b�T�鈼�?L����K^u����K�t%���6:��]��H1�椄�1�3�{	�-�^�fH���Y����g���?���H���$��=����ON[/���Ԉ{(�r�
��q�	'���2Iʩ�l�0Xrm3I�~��K��hH��k�d��zs�@�Hc�fJ�j_Pġ�a\�$�������j�kFmɵI�����j�L��|9��~:d�A;������-m�E���/	��ץ��tTW^E�T���i�:�c'����� ���x�/"7)(~
p:i�ݨ�*��g�R	����7��#�H�e��E�P�E�9��|�ռ҈=)���\���L�#��]�{��Zw:��h��Vw7�;z�n5Y<�&�ᒈ�m��N(��	4:^r0(M�i��Y�y�_�p�ˬ^�����S�(�2�m
<,T3p��_us����4��!�LzX�l��ֆg@�Zh�F--7 �]�UxLz����s�&��	�?�8̉�����c9b��u�����fn��op]y)��K�:����/�f��DX�a��#HǼ\�=+�l�+�T{�ׄ��F4�hM�d�����9�x�/Rq�Tڏ�������O"�r��Z&U��.m�Vϖ�~�V�i��.{N�Z��B�����|7�6ʇ��l�B!ϸy�{/U�$(�;0Og�A�~�:�Y����Ld��Q�~#}�<<���n��&R=N�����r���m*)�glrW#WR�w��L���*Q�mR��`�W�.�%Z8�]��hᐹ�<&�w��7�P���]�%�}c���؏Ir��f�S*82�s���b���������9F�*���_ms��ҝڟ� ��k�jG�|�7:j�=�]�H�E���N��z���.�@.�U\oR?�	���'�����+�P�U��?����N[�uYHzG����IF'iD�$$jB-ɗ�����r�����qGjK�[dE7\��H<���0�[~���+�N6��:���uR_�d����ɥYM��P�SEt8�O��U��%�,��-�[�ω�UlC�� ��/���\�4y��m��E��="��3��O�d���|����c@��\7�_�_YTˈ��9�n�x|�����IJ����N���-%QZ�+ �@���<�T!.�l�D):�YTx��D'o���:���D{m�*ܿh�l�2)�\�v�I��?<)�m4�!*�u�j{���J����f�Cx�24����L����T�©;�8���yr�I�%��e
�($VPF)g���T���p��̅@2��\'O���cg��q�u4$��oɃ��hIw������O��14�͸�n�c죑��J�nq%7c鰔 �ZG�<�h  I����\����B��z�Q����3�90�	Y�)�nZ�K^�b��n1E��5+)I��N#`@@=J]h��"�fY�B��U�$.������S�N��!�AE$f����`���M�^���vP[�^�*��h�ՖI;��5���:��<
��Br����$+a5�4{?���s ޫ�#�$@1���k�6��L����~�*X �3\*�k���d�i{�n���R�M���x�d,3����vʚ#�Z��g�	�,8�O��U�_}{���e�y'��/Ҥ��ղ��~]�H@
h춸0��i��ma��Y���?��}Nݏ3m�9�ߙ��)����x�����E��,34%TN�#�B4�8����;~O' �	nå�40}�O���S���ϚS�\�h�(�'�O�V�aٓB����wZK����J�z¢�L��:!ouP��`�q*� �-'E����í鉀
 �HX����x��mY��s����8�	�y~2�Z7�WC����E|�C��W�(��|��T��>���lD�� ��@Z�|d��!���,%�LBb�./��2&�qG�-+ϸIe�m�n@����i�i%�@�8MKف�cB:�`�-���)�S�ڲ�d�	���'%M��@��	�L�⿊��3,�T����S^,x��)w�q�<���<\O���i��J�Z�^n��BMvjr>��ӫt��Ρ�E�A�b6fg�QI���/�+���N�g��|��sBWlD����^��oG�n<ۚ�&Ю=�g*%g�e<}K˚N�3�d�Ju)��b$
D���lwJc��RrTI��p$���A�k�8�}�zd?�ÄV�*�G3g����hKn;h ��X��7٨��]�x��dzl�n#ɮQ;9�� ����IPpW��p�Jġʼ�'�`/Flj�9�ۗ*^d�;��j��_vI P�onu&��Y6`Pq�Y�Ka_$-��Q
�^���<�BcU�.����a"�8L蔳��~+��]e�Ю�iG����3�|t���*B�t	���&�Km)��g3��� �O
S�1�.M�ۼ=����'8Ǒvb^��2���К�Y�^t�����b�hnsS�V$|�.~�*�m�;�uh}'�p��ñ2m}��Vso����E�"zx��Ì�L�}�y?��s,`����m�$��t�q��/�3�~��J�pP먹&;���\�%<<�1��i��(����G`���|ET����Q��$J��S��sW�XʠJ���!z�sr�b�>'͈IU�AƮ�>����K_��AZ�-�c�c�!ެ�W�(������
Ql;@����ъ͜[�o%n�B�Q�9f�;/��@+A�~�G�~��֥8��]B���>kv�n��[�d��7}�4^��HJع�� a���S�[��d}����Nʻ[� �����M���r=� J'
�"��9w�/�Ƙ��8ئޫp�Y����P!_6�q���9��a�ܺ1��/����my��� 9�o����}��Z�NJ[);�~1bp�Y;b'�Ƃ\5,��,���ي�P�Vl��C�,t�'1rIì1��1�Ȗ�`�=�sX���nU��C�|��<���n�?��U3�Џ����"�n�-�VL�
D.�6�O�a&j�ʔ�!q���Wֵ�`�_9KW���`euܪ�;��Y�3i%\�ȤpJ���`�RiK_(�}�c~0�&nQt�iU)=���&�[�#���l�ϛ��f�M����9��[�*C)L�I�z�Q��{W�Z�|�ġA*x�.�����#)�E1���h�C�0�ǁ9�x$� Ab!�ͨ4�u� ��OXӃ�4�T����Ċ+T���.Ӿ\=��J����x��-��ݟ�/�����l[]�ӛp7�F�$��"�N��Q���yPU@8�L�4#����"��[����*�{uv��?���y1���=/,�e���B:�\$"�[��7[�g��;�Sv�x�L���Ѝ׷�?}_�s1 �V�	��k��@/aD�}kJ�8=	f+R�0�I�;�&*Ow�5��ݸp��oJ ���H��u4Ǐ���ߋ�'9�_ѵ6��I��/ƴY���-��x��]�1�^F�<}Hc#���'���-5���Q��&�W?2��O��v�S��F	�&�������l�/������#vG�40"2(��c>��hy]a�2��5�ք�(��	$��Q)!yF��%-�OI k}d(�.m����YR�l%����զL�7�A�"-�^0V���/����`�n� ��]����``9_UҼ���+��ϐ�p����i"��oB���	(����/�
ݱ�z��c��8W��ꪇ��vءO��{��l��?ITP��{�a]����S��{EY�E�'.����y�vA�Ջ���@�R'^���A��jC�uA|�֍A�J�Ȑ���~�φm	�0{�D��c1⯩��^��/�K�q��F�̬�^������$���Q���c����Q�0��6V�q����b�ߜ�\�z��K/됬���l���"J�`�pN����d=�;�〥n��s�(T�0<�-��n�ω����hV��m+�DW�P�.	����.�i�^0)���}�m��D��B�	I�,0\���պ��M����@���Fs>���XH�~y�8r�f��P�S�iSL���Ѡ0��%�}7~͜_��G����ėA�v%���1h�y(�A��71�D[��ioDF���4��O��@_q��cj�ͤ�5��vx���uDϘ7^�4��>�R
\�س�B�6����r���4E�R���z0��*��Q|��ɖ�H��ϥYf�DLm�;�U��Ӗ����l��R�\J�<�ȑ�AA"ħo
�u��f�ʃ/���Vаn�B�',˧Z���+8�q]\k�����4�3o��ô�0�;������#yl<����#����}@�*����r�*xeT��ψ&��o��㙰�f�ʸn�����5�-��N�0.ɋo5���9���%�Y_��O�:�s�ف�g��5����UL�A��M���W�$bI����13���k|�8I�8�t�}�@W\9~�GE��+��[��m<��{{��)����t���R@g%:����^LPi!�T^���B+��j���E�.��Y?Y'� ���9�;FI��0��a0�:���y���5}U*��m��22�QM�P��[�s����8��F���;nY��Z��a�.f�r׷�8�V̋ؤ.�j86"0W��H�v6� ��;�W�M����k�nKȞ�	.;��,�aTS6f�{ʶ~�iT�-4�����!L��q}��g�n�;+�k_�#z��{T}a�lV���;^W��ǝ��硏8���oR�w@b*md�>��w�nj�E���q���!,T_���*�<P�g�nJ���PlM�l�R��Nt���w7r�\E� �Ji��HM`x:u1*���ڙ�o;t��
��[&\�M��C��'�5J�n*�pb8�.,m���E�Swo�������T��!�U����2U'cV��cW��ؤ���n!r1s�8T�����$꣞�!��� �ԩ/Ë��1[,���\�	iNh�y��X��P�h�R��~7���n��a�;M�t?n�����o@���$[��L�`b^>O˥9E<��A�r\{��:f�5�>�0:ĩ�"%?.�k1�<*~��
�{fȗ]�:N���!I`+2�t�O�T�����ͳY��1B=_C���(˒�uuMܿ�%�� ���f�������M`ə��i+O`R��de�(G��'��4��d�(������x�*T��T�wDi<����::�o�a��F�nU��挼�p��s=�� ��N2��-����{*E)Nი�z!v.x@�O˥�`�|[0�{���(�+�e�^��޳%n��L��]i�~e2�@��mZ��+�?�bt�W�>-(�u����b:'s>��b�D��~���ܓħ�"3��^{��B%���
W�Ҹ��/
�.��ǁ}�7}�5}�j����~��8S�|Ԡ.��;e���|2�v�L��v>���=�ah���i�n���MPsM�;��>}3Υe���O�ʔw|XL!��Ⱦ�w�|S*_�ZZZ4;�x;�y��3-�
�c6��^wB�e�0��D�A�l�ͳY_����`��� 2�̕��5�C�z�;�tv��-�ݒl�Ie���|�1u��7zK��\�U�w��g��pK�ba=`�Y&hP�V��&��4q���#���}w9=5�:�{�-o� ����^)6'9�}��~ M�m��`�܇g2��f62s|�"��	2�y�旈�u]�jɬH0�8�J]�T3P�=T�"c܀v~�:�0��kF�J� �T2Pt4�8�Y2)^}o7*fS&��b�����F�Է�+�9S:5�<�~�-h���k�}����>�I(ٰbc��Z�8{�\;3��K��ko~.� ��p?;�� ���l���i��E���"ox���eq�Bwd�/6yg��6�Ғ��H6���⬁UE	BĢR�T��+v>��<���;N�6a3
������JLsaJ�4�HS٭Ǌ@7#>�)��Rpa�zw�FKK���pI�*p���F�={N�z��]���;g�W7|+��R�P=���O��Z�'���*^�H�$�]O��Ť
$�dsoF�������ߟ���R^�12�eQ�S eij�MF�2B�������^��'�`Y�AI�q.$l��5��)
݇���>@��Tړ <���,n�U����O�v�{�m�U��"Xx'�O�ƽ���5�O߷:]�6�q���6���2�k��{}l�~�y�}̡��)��P~�f�2HG!Er�e?iJG~��ר���HM:d�'�X'�%4�Q#�~�H��l
.��W!](Kת2ף�J�͂kX������b�~��<��fv���&�¶
��E�(�	1y$��n:ʬK��U�-�U!�����@i�ky��4"������a�#�u�����E���2٦´������S�#�k�?�����;�S1�����T�E��Ci�ʫ�Lt�(i�5�\*4��U��<&�p����ȱ ���v���7Ć�,1J�H[�[I,�]sLA*s<�0��E%dXWz���D����0W��ڍ�.��C*:�\I��R����	��Y�Z�!�����A� �x����.8��z���>�"c$Z-�(7\PW���ԕﱉ���HC�������)3��{.K������#n�+Z!����m�V�&��/P�^��eɇ������ċn�S�Z'pn�P��5Tt0R��F�pH̀|�-��̵7KkH8J���⣡,X7}厷��Rm������k���s�&�QLl��-XM�=O��X El�χC�J�̞��pn�4��*N����{�N���.�c�Z���+��H�7����
.h��/M�<s �u+�CH�f��?R�0�R��p�f]���&K�vt[ُ Is�9e-y�z���@��nI�����nP2�RO����L��Ú��="r۝[
��/l�̍�~���`FSڵd<���ʪ=q����v8|�5t���69w��K�3=��4�	L���Wv�It��&�����_�Y�ٱ`�~M���ƒ�>��#;��U���ט0P�v-�A!��(�}
��"*�:H��U�tPo��0���C�"l��J�u���������d�m:ɬ�9v���8����������q`������H�*!O������l?r��m�Y���:]��P��5$�f����,qe��F�����xvo)�si�?����/��y�R�f@��J�nJ�%E�<�����A�k羁�d=��~ y]M��_��4��H��圆��S����O"�S�Ͽ���-��B�]��ek��`£��d N;fˡ���l
S��F�bN�b�z���Ij
� 7�|��T[;�a��LɂJ���ȻX&��Yc�/!�UV�`�"��Q����}���Ō���F�@k�t�SH�i�!�M���G�Ѝ��n*�&���CDQeNa�h}9��Ԫ�7	�^R����#i���~q�=�8���QI��ŚF1l���~�Y�'���奰����g���Ch]�$�F�y9���/�\l��B���rRՠ����ڌ{��^��Z'J[��g2�<~A�A 
 <ua�إ�?����OU������A�dlru6�������ü��Z�ũ��,"%=V��jiY憶wg��诌�{$+�ϱ5��6r�ýy.3s�X˓�#��P��ڈp�e��A��g��AU�5DaVd.��زĵ㵅�<f,����H��J�:����|qg ���x=�><�R��32b�j��+]��6�f-s�~�I�Qκ�sL����:8�S�����Bbn�wd��#�D{��f[%A�щ�*/�HА���	�z�g�l.4W~=b"X�k��'�3��t�*��U��_�6)��G�:~CV�"h4��;Ym�8[�/b:p�8��`To�ʒ]�=�~miw�Ţ�0� ,�Ƿ�y9�J����	2.���]ruO�u�aYH}6nv���۫���`�78e��(�_S�wWx�ˎ�:ԝE�
�����@cʈ�JY],t��k�g���I�����z-��t��蹑B�GA:�_����Ce3u��v����3}a�DyFM��l��B;��W	�&�V�ܼ Tf���X�0���q�5��	Ӄ�7|]�Vl��r>�G%�{T�~�i&`��x]�(s�C���C���K�
o�%);�`$�{ׯC | I�x�!�Qv��&#����>k4��\��Oq��2�'�ʛ�Ti\�8B�.�����u�,�W'ͯ�L��!C��7\��M4ѵ�l��������V�cY��ئ�?��{��E�}���@dޅv�R���}/(*�����!����L�q���G|f��H����.�Poç�$�K�6$��!�ƾLu�ntX�c��jMS�/�Ù{;����.�M�����#��4�m�//z�-���ƌ&]a�jw���tݏn�l���I��1�y���>�/nJ�`dމ?�=O�V$�A��[�	�vQg�"�-X��̚ے��Xo�A�
E�ۨ�Xu��k����u�bm��,+�D��&�[I��e",MӡBp�i�"[C.S�Ōr���2�I�s��M�L�B�\� ,���O�۵c�Z��W��u
�YKPk}8�M�	���}�דܛ@u���TG�r����t��h��m�3>�R2�z�)�~�l�JJк���z^֭���^�R�"���d�O�|�s���3�.t�@�J��2B�u=�I�T���0?�|7F�1���+]zΒ�����n�Wz��ŚR�
V��'�
�K���V�
�>y�:O���7q�~?��k���R�:u����lC���4�}�%~�͘�@K�\��T �_K?��܆-�-�
cM�I b.͉i*�I t��P�ϱ�|4��<h��:����QĽ��Uq��e�%8��@7���2��{O���텵u������"�1Pun�͌������ʴEI�@��v�RF&'$��-qwj�q�ݭ��`H����͋Q_��[b�ym!�UZ�F����Ad�VAfC���>Ɛ_o$(r,����������ӯ�-��a*Ox��%�}���"L�yɾ� �-��f�&Q��p�dK��K� I�b�G��j��x��v3IҚ��������7�>uS�	2���4YE����u�я��:�rb[��\_��=m�.�#�sj��X�.⩼��W�����ب��VO쩳�ı�H�=��wm�peTZ(��+ڲ�����	uk��Ӟ�4[�V�^��*z�`W:겿1mG� �%n�����5ɾ�"v�K�T�q"�c���Wqw+��N�3� ��C�E)�X�r����4��b�S'BWK1��V^Aq �������B2hUG$��D������:0#�HЋ���R���P����K�%.x�0\� ��׺��[�3=�ra��2���5<�� ��@�fAœ��܇k�A$y�tu*h�X�:AR�A=��H��*�����ı������̴�]@]֭Bd��^� �p|E�[�Us-����T�}�ĦLMG��`T~�.y����$S�R�L�f�sƞrf�{PE�sٿd�Lǰ䙿�fLS��[�d*���2u/Fx��At[1'c���z&�\�#�7W� �#Y:�-�}�$P(8����t����a#�4#Yml���_�>C�
����,�T�nP���u���z��������cY�iq�ϳ�68�B��1�)�r)��1@*x"��S�+1�j��e�;
�Q�RE����O5Ƞ�מC3�������9vl����Zd֜q��\�Q/Q&���e�a�X:Yw��x��+��n��p�n��˾�2�i�F�c�E�p+@ر(�8�q�P�H���R�Zi^�
���� �0/d��l��m�5��:AގX�.�V
�����`���|N�*>�M�5J�|����xIap��� ʱ�hπO<���U���N���K�j�-���p�}2m�/��d=�u���SkU+��pCcG�=����� ���b�֮ U��skK��Ҹ�/	�->;�Yԝv�`�X�ǃ?�Wr�#Z�0��L�;��P�~dfU'�Jp�G��[VOx:���=.z rO�׸�A߻�m����RtLY��%Y��R1E3q缯`�2�f~s+��P���5G��u���
�a��1t�����T�2��`2�gf�1P�矼��s����6Y��a8P{�4���S7�y\YF}+��Pvn��;�k�2[�u�ʏy|�t�NQ�˒�;���O�i�~�1'l)��Gn\���H2�s�LF�FwL��B\�V9��J0�Glt�3���?]�w�#�����̅�Cw4c��G�p&������Q��۽'�d���y�\��U?��
u�Z��w�Jݶ���{Ӂs��t�����G��m �6fP4�\[��A#D<�Xߔq�`ѯ���U�[��U�`L�vY�ǭ��_����y[�p�Iz�K���8)�(u�[�2�u�Od������(D-I�����e��g�^���J��X���^Ҭ���u���&�����G2bc6�
��4��y+��˥4u(?-8HE�5��˜�#���E�4L�n�x�o�-NT@A��/���aK���G�i e�M�u[���v�R!��NO�:�oCc5�e̹͑eh(���)�c��շ���B��"�o-���o���Cfa@�Е�U�i�j�XwI��W<��p���0�V��#%����(�F	2��(�?p�2aS9l�w��V1z2],=����A���B浕_�Mi$�	U}���_���7|'���R�#��&�*1��;P�0�Ӧ��L%!�rk��,�3*Q�����҅�O+|�=Nxe�a�x�2�6��5���UViH��mt��g��}.>����˷i�)��`�+B�"H��p�)c�g���ig'�73F�/��k1�]uT�.=n��`��=��"�4e^�,�P6�.��"�f��	���]��?x'��c�s|y�ҒdR|��<������6)W
xRD��Ǝ�7�aȔ0�s��� �B�3���(��'�ćv(��v�{�E'�*m�.d��A��^�/y|�s�ik����Br|�D~���m��X��ЋuO�T�ʁ�$3�A�2��s�ё���rg�)ZP���Ὼ�N�J'۪�W�O��w����Ƥ�T��\]d��I�P�(����E��<�=n7M�ĵ&<D�_�*UL����>�qa����Pq��jbRP�LL�q�A_��sz�E������ά�s2��kMYJ~�}[��D�
��YS��f���'�H
�,�7�iXf �	.��kg�0�V�a�ilY)}z��V�и��` �����r,�S��y��g\z>&��AB����1$ǎ
ȸgvju_2�~�W4Br�φ��i�:�]��.��9A�=N����u~[h|��Y�b��wFE��4-��������p�c4�b�XcE�D@��LO�hO�����/�@k�ڑ͇#>y�,��!��K����Q���r�Jt�ťZ�!S���a�O��ⳂLS1�����=�ȅ2�M(<�8%�f���{�"X�)^{[K���f����4|B����h�b�_ �_�P�f����h��4NGm3<�i&�(P ��*DQ�c�o��d�i�q�y%�;�K��?�9) *g4�Xэ��d4D�N
%��L.��3{�E�7�c^H|̻�-��!��Ʋ2=��x�É����/�B3��2�I[<=^3V�:`�&��k�� j"<�o!�A�؋�y�3���;Z5s��;�J*��Z\��l�ĺ�o;-���mr��Mp�|X!��1�q��&������&IշS�O���r�1Y�}7���,.1z����㜑dp(?E���V�0	
"�j�2t�ʇ���'gv��t��`�ב7}t���?ێ����[^��������x�H*�Ixa��w����pC��׌�*���[�}�
�]E��r�f��a�J-A%��h�S�lM����MmQx�  ��Y%̼{s�Yƞ��Kv'�����/�w��k�%�x��
/rYW��,���ϛ� �h節���>��ҕ�Sx��_ikN�AZ7�;�/8|�]��ϱ�e%�*HX^��[�@�3��M�����^�À}�G�۶MI�\���X�F/%�w��Vx�i�dͷ��l�m�ˊ�ǢV����k�~�Aȫ�rb�Z�O�jy�pǔ�j�1n�d��Y�e*���J�	,�
Y������K��+���=��U�%ݤg^��6r(e�
\}�Cq�v����]��!T�'������l�$�K̀}܂.0��'\,	.A�*1��i�ד3���f5��s;:�z���n8\���.�c6{l
����pr�x0�/S��C1i_B�Ȟ����:6K۽cL:ӱx�����]��3/JZ����rSJ�b��1ar��e);l�㷁�SZ"�W�N%ql=�x3{l�l![b+��7���	o>�����c����6�<�
�ˁ��7���x�������g��E��'� }#�K=�\�Z@r�tp�hX���1�F~�y�	��=O���p�[�<�wu���p	��7a�o�x�r�*&�|ګ�����x&%�/A�+;�o�	h�Yf��R�W'�u<j3o�G�jVz����V�Z������9����A���c��K��6���P��u�O�����7<�.};�a޷�L�a'qŀ�Q4̵���/ �D�' a�t�.���4�lD�W�OPu�h�-�b�w^�����k�@w�Cn�V��^����.����j�Q�m�����Cb�+�K5%�����$mLq�9��8�jWb�FEd\-�\���<z�x`*�k��e�A;R����ȭׯg�F����1����SU�0s$,G��Y_�J�^zņ������Ȣ��D�4�vc��a#�b[�B��aB���u���%h!�h:~!Nw�ʍO�0?�bD �֑�c邊����$b#T�p��5��Ff�(� �DbK���m��7�:���f�.�� f\B��+�~��L�T-�^�m]��,�'=�\)-x[��)G�bxO��*��|~�Y&m��dj7�j�q�-
��N~��I�3�����ԁ5h���9�r~<��x��ل�s0[�x"G������σ]gq_Ov^&3���ۯ���p���2L~q�+#s0�c~�>/�(^���"�f��V��>�ܵ`۴�4r�!c\
�U��\�oyU]G��_a^v��\���V~l���c���xc���JNS�����v�fI�eW�0��Q �&y^&8Tm��i��L�,)���JpV�w�������kIL���O��CG�����0z���뻑���p���	���*
$��p�Y������ݛ�pZ��Y0��N��}��0� ]�2�l	�]S�3�ޤ@uP�r��a�皹X�n��ծ�=�ލS�ny�U;�Fyk�:��S�Bݗ�G �|�����oH������FF���[q��>J�LPh����t��4Z�O
v
���������x\���#O���bh<�f�����7�fʗ0���\��l�����}^�����܏`�`��~%��y_��`��?4�w���Λ�Wv����'0s�cHF��>�!���%:qzb�v�k�BKc��ꙎF�&� U�X���e+^i��,�f�و�B�h�L �O:�\����Z�Q�R�||t�'�ȩ����R���b���F�2T����%�����4���Ԁ@�9����%��-�?�����%Q��jn�?�R��1I�u�
S���ɬ�O��������|Us_ղWr���؎��yk��� �N$�`��f�Ȋi�-rn�,T���_�p�>���Y��n�[Bmԯ�#%�ح�A.=�'�X��؍h-E=bCs�`H�+�ҐWD�q���^����\$zN�?����:O�9�䔅�' "�g�J�Kየ��9�&�PM	Ԏ�JMQ�*�UI��!*��8K>`~_�����)�Akk�3�U2���K��Z �r����S��i��~P^%���bD�},�L����X�UW��w�F�G�@e_�9�4�b	�f�n�?��;TqQ" S���kJ���F�1Xf���U޲� ���hJmp�q��h#`)��àJ?�5�I��c`�q�������V��{k�,�Zg1��in����U�0�u�*�[9��<�' �)��=_�x��|��?��%ҵ�l��/w
��{�WM���l�/�N�v��
�t3�v���nOK�vZ[ӷ�%��և�b�߂���߽.�t�h%��H�G�I8z���+�Ve��;]Ԛ�O�"\4���6S3c����[Htҽl]��9�H��f96�Z8���|�/��ߛ��P�D�Hཝ*?O
�q>gW���PL��wR�E;��z�쿅N`��_�Qs�+�Ia�i77mrT����iWw� lN��g��z��Z�{3����6�8ωE���Q����B�E�t>Ua�;ꠟ�cjՈ�����A�0_��$��G1r�^^��-ω]��GJ�6�L�7�S�3�fpҗ�$؞�;�@8��C��\c.� 5����R�\^�^�G�(��E~=OЙ�WjY?��c*�mX�f/� Cs;T'��b��)�9��]��庼�mއ�����k=� &^ӏ���y�3tKפ��^nP�W�G���W�Ã�->��5�aQ��l���1�r��*�i�ed��9� m��R-�9{9A��x"�j�e��pD~��8.�O�<q����O�>c���H]���n�������H>��}�k!�����v�_~�L��|(�/"�y��rg駞i�X�x�u�W��FFͫ�-Y�V����U=�n:7������z�A�=B�)�G!_� %ؠL���~JL#3�C$�?=���.�(����r�D�RJ��I�]���wCk�kw=�f��Ǒ���щ��>��IX�ޟj�HȉF�~�Ru J����Vyc��󙓢��qB l�3������B|�h����8��9�/y.L�\f�no������?�#��^�*//k�1��ٌ��#�K/��<���x���B=�8��qժ���ު~O1��8���^ )��Go�V���<8����������9&("������o�eYө������b��y��e�s�}5=A�>G�/p�5��WؘMm;ǍA����j�IZ��"�Y�����fhՀ�����ꁁ���G%ᗫ݆{_'�t��]P]�h ����d��KU{됊bM6�'�����E�}������kUI��Et�$��+ck��ʶbp��z��
�cv^	�S���;Eť��O\��&"�x�G�q��E�/�He�!Y��%c_������E�$�Fdk3���2h`�h������\f���T�p�L����[���f�D��E�п��	��by�oB�f �Y�$�0(�-�u��}ɾtC�?�z�=�3d0t�0����2�]M�#��̱���~\��A)������G
=���F>Vg R���1��y��5Lw�ffv �*�;���_��8Q	�,@��N�L���?e,�����.�E�*�=�S7K�FFz�%~0q��`�_�@��@9�D�m%�j�_.}���_:o�Ě0��pvw��=K�]*-�y�'�Ls}�q�kz��,g5ŝpX�Y\����w5=u<����$đ����xײ�E���Wm��T��f̝�`� r��֘;;�������ۛ�ʻ��{��^g�F65��C�%��V&I�&���l"0�u�ؖ~蒪��'��e�>3Z�:m��xx�_��3�"Bo���/����$�f��i��2�!U��{�Uޥ��4��	&���rD�\L�l����:?��z!0��2�;Z#�w��_�� ��c{�̿�"��M+�L��RƬ�oe�Y2�#X`�s�t�iOZ#[\,���L9���n��`a�;�\�n^f�,-q� �=]���(�i�J�(��^�$�j6�����laB�>�I�v���������O�3@I#�Y[��ê%UA�b���%�6bH�֣ *�ЖW�H@�\��w��%#�mh�쭗@ߍ�CK]f����h}o����kU�OJ�(Ί�6J[�C������#�I�~�m�U����A��$9kq��ϓt$7���x(Ӏ���6�(�-6I��YĠa8R�N�蚓��O篇�	FZQBi2��\;��(�Dx�/~��Yug%9�*PYg˽�lO�V�z�v�Q��]��h��^J_��-z�8�}&V0`��C��p�lE�Ӗ�;�a��c��3X綉'��3���l���>(8�R��1�Jj^��5nJ���%���ht���ބJ�g ��^UiJ>`^UX��y�I~`��J��&(گ/��E�%���}��e���ֆX������Hפd�-�^�4�e��E�YV�-���Ƶ?-	L�T��HB�N��(1\���8
�o?�w0�2 �&vK�Zczz�����AGX��Ղ_ybDf��j���i��a���76�Û�9o2��%;)��(1����Z;^$(�RI����}��X��0̂yVp��ZSף���.'��?�|����q���3DH�o����h(�������G)k��0JC�8Jϟ����Ȋ/i�c�"<�x����Z��)
��kH���eu����o��ԙ
i�0����o����O�q�%k,�''��]O�W�$,�>{��!ß�ۓ�Lc���D��O�m�+�Jt�?�NEjd��
�.�U��{ye����L�D�i|+����Y�QWcf������&	�)	5��õ�!�g-tՎB�Y�p��z�������o��8�k<cҌ�����.��{>�G.�{�xd*�GC�����c30�jb0��	�1q��]��U[�P�����OL �藕�~ݭj�˔s��s_S�Qs��}p��-p8�A�J�@����=8����?D؊�9 �S�{�N�4o����i
���o���ݩ��D0���H_�е�����_�zn
�Jz�cY��V�8����uRЛ�	b1�~�����ί*�ۆ�,G��HZw���^�9� ��p��ђ��@=��������Q��`�,4�n�.�	��B�����Ѐ��#�D̿)Yu�{$�L.{GzhE��/KU!zJ%U�sa0�[Ι���ݑd�U�h4�	�|��Է�v���ȓ:�YJ?�RA�-ߪb<g���?N-,��� 8������aNV٪���'%y`"�����MVf֠S�6p�D�4u��k��Q�,N���7PYcU됂���(��q��c�ʄ*t�5�9�@^������Uc?W�*��2ɇ�����N�.�6Zӽ�p"mbKP���.7P��v*��q��8�ES>���4Ca���2ީ�KцL�Ju�h0ŷ�G��x/$���}�f��毕r|�nD��z�
�pbӀL�K����&AJ��l@ :mj�g�_ci���b3@!Ҧ_��*/�AXq���j�ޒa���;y7d�d�C�-S��,���	%�j�ܧ0�?#;���	���<�v���g����o:|��y�,s9�`��	b;��\l�!*]4$�$w;��嬫!|I�}�se��ቹD)^bF��1���p��(r���(�LO�O�T�pZK5���J�9��Ǐ���Qt��[������rwU�hg{���E^x>�҄�P>��6G���Ӱ��N�VYsj>���yJ��H�������o�o�U��+<�I ��3Q�tV]�s�
��Z��/��zώ�$���5/V����+G�f�؛\���HY�w�oQ�
.�]��Q������s������==��ߘ5�Lu�x�%G��sAbID�<�c����-V��2l�*��N�J�&�\�����9���E��=}�v����iRY`%�������1��t��`��o���D��a����3h�\��T�/��N��E��̂5���dkӍ���V+F ?F�Ep����T�� M�xP�!o�ld�ˌ0�(q���j	O�����ۀȣ/�%�PiｽB��/h���D�#��و�体� ד8CX;��vK��ša�n��hj2����(�����x�x��g�y��7�z�Ǹ�}i?����ʛ�s�dn��3��m�u���^�U�Ը;ĕ��Y#���\}�Z��x�� �B�A��~��0Wn�~��U�.��r9S���F�� �-��S�0��6n�=�����a&-�����m2Η)�8:�U�����}��b��U	���vqdJ���K�U=P ?0F&��;ٳ�������f9S��r���6�Zm� #�5��J�p�Z�|]�ΔśL���b�q��a��$auy{��aT"9)ٜ媞Ț�:��+�n�&����R��"A�: �6g�	��Ӑ-���vM���=[.H^�B���K.�u��I.8ȶ�c0Z�4�&t�!���ӂ�{3�Q���R�3���7:�-$hqţ [c�tO����d%nG����ZH1G2a4�S�ʭ�Eid�q�+ �f�w�D�������%X�}VTL�w�$ɽ��io��ݧ��l�!�u�D�4��|����5��2�5�*^��!,����˫���>#�R��.%�Q�5E��`�*�-?6�f����LB(�6x�Y�U\�R�$����������ܪ�R� �-��N��́X���8I/ؔk�+��Lٯ��E����gܰ�@���}ǿ�G.=�3�Q}-��� 2�_�B���2�Q�y��2���|��*8|1Ӎ��|���9��r��)L:�����>
�(,h��0s��|f�e�7D\��	�T�9�G��ڔ�<Kx���Wcg�%��g��bS'.���%�Z8��
3������C�l�?<�	�ٸ��pX��k/.�I�]�0Z�%�\ ��W�����J��g����d?:A桥��
n�0�*��ǻ�Řy�� XS���ƞ#~�ፍ���k���m����%�2p~��7A�'�)��	Y�l����M����6ڎ��OmWN��ꛐ3�$�v��W�OP������ӄ&X
_� 'W��g|5��q�.#�u�=R�I���=nJ^ceE#����-����S����ܓ�!����]u.H�<��tV�j�5FW�C���&7��Y�{�W�.O2Ě�h�,�=-�$�▸�e������Q-�K��/'���f� $e���8�O���|��mb��X�	9�����˧�M�[�H�注�c�����>ݶ���ݕ�Ǉ���}����P+��=���`ӢܲU��w�0�~��'���i�NBz���񋽔�Ƴ)9o���cj����o~�N  3���	����m�8���	^A~�=�����l�e�e&��9�*YsSb�z�V�{�S���)Cq5�g�Ф�Ų )̀�}הIF�Q�뻤�ތm���O��s�rtA��Ƹ�;��/V�CK>�d��WV�9.�Lj����a�_�(b�R�0*�]L��u�Y������!���d���v̎�c��0}�|N��y�*֚��C�y��A|%�o�#�6"�,Lj�Tʤ�ő:l]�
��!��L������(�ֺ�}	����8��=��i���쉫r����W���Wv媍(�}��P
� �O_��%O�з&�yQu�7���G��+7�p��v��q�A��RJ�EP.�	�+�&�Fk �@W�����:&��~�?���Zc	�+/�ǝ) �YK�%~�Zz��t@F�8a���,��yX�q�q�E>1��+����k=��HI ���������z������7� �`*N�珳d�;�g�HL��M�>��%(��≏���4#���ό�`���ndJH�\6�i>�jb�!��Ij9�:�Uίm��ȗT
X&��w!I�V}'ډ����_3�)1�;
i*����<�B�0����[H���7r�A��aa��N�$H:>ieug^O7�����i��a$��N�
{Aq&��RY�E@��cw����F���x��Y�A_[�@uī���&���g�)���KlѮr���9�Z�Ā�as�y�|,�2��#�J#����*��8��VU�{P�@����pN��ԑ��;���c�^��][x�4����Ъ����r�P=r���}�jܡ�;��i���rGq