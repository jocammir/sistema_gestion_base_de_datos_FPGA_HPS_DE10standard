��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0���C	�i��E����A�Ĉ%ɲ������O����D�v<]�vM^���r_��'�j5Eh<R���;�y��G���2reSo� h� �����=Q�96� �1��G��ek
�<���^�� ���t�0��B�F­Ǌ68LX<��An:��`��e�����m�4Ų.�Q�od�5��b�8�$�mz2�-���_H_������H H��kd��CE��3,?�w^��0.����`���4Xk��wFz��@���P�������g�3pRNq�ˊ��Fz6R�?#�cc���Uk�A��Oے)�V�Ib��_���x�p5P�I�A��_�A�8��i\�W�%?�.18���/K�\��u�Wx]}��5�h
!�&l��ػ�����}�N/g�TED�Y�b�龑F��;�FV�ϷZI���)�rv��Q��}���/���k&��H7�u�be��1�;~Z�i�Q�Y�8��4�U�Q�c�?�W B�;�$5G{ԝ�H���R���Fl=�?��I��_:�F��H�  ,�<|�ޕ�̾��B��M%a��yH3"����l�9"N���o�@	����F��E��d؉�sDN����j=��
}�]Ҿ+i�)8�Г�A|z�ۗLtL,�<M��U]� g&8Y}y�������0-/ �[gX�A(O\|�+�d^�%N1��

�X*���3�����F�7#3�a�-!rI?-m��믜p��3s�"y�I��M�>D�w�8�٩��ͱdTYLG���i
D�ѫ����W��*/f�R_���pf?{3f����5%Ć��Q�>tBL��>����
H�W���E�>�!�g�B0F,@�#j���Q����n��dx�q���vٶB����_�I��}��_����6����-�:SŞڕ��{�":��׫�aa�y~�<F�;k�L�!O�c�dV�P6�6���e<  k��kr���"�k�̔;��\ǆKE�]t+~S'�F*����~��:ʗ,���t���Z�,�iV�a���	M}�ԀSK>i������c�1���s� .vD������ݗ.��Eso9����<��3�����;��x����ï=UnFJp�3�����4.�1no7d誇�R�t�9�]53��K:��h��b���婞���XN?�b2����%v��"֌+�S,���,Sl���8�~kp���CǊ���9��^>>M�a� =8��s��XA3=��|�>v:<b��D[T�I�8�%JP���T�o�nV �Ap?�]Y�[}�����F��[[�IZk���<�Y�%՘����e\e��`���n� C��p	D��>C�6k��<\���C�Ht>�������Vf���_x�j4���+]�}j�N'�ei�3���{���\M���8Ϟ�1��D��"���G���N!"���q��R�@��:WI�3#m��FhsS��A����]˒F;$�kj�N���٫�F���~}kS�6x�]�j,?��~ou�f^��4��vYð�1y/V�uAw���>��$�h�`�-x/E�w��=�(�rsg�������a���� qYgq�}��K��A��+,��Ze$w+�W�����x}���?����5���jF�7�d�uC����v��=�dL�����\˷��)���8l�o<c�OJB�6�YOMj��zq��"d#6v�Y�֡� �sT�-k��I�mO�v|��ŭ��U�?�`�v�Y�n��Yk&�e_YӸ�cp����-
T�(����Ojd�m��'X��}�:;=�g�Ync���y?�:�Cc���nr<���k3 @���&>vu�X���G�%]����	*��ګ~�ښŐ.�|����F�ۖ�rwxMy�����	8��2�?�է�g��s����6w�e�C�p�݇�1��C<���	����'�q ���s�D�	�f����>����� �"&P$7y=�����|Kc6�ǨHe�*��y����	v�x<��SA�Sywes���db����@��I+��.��֞�舻uh���;�"z_�i�d��xşw#����l&����T��ė7n����y�!JL����M���do��$�W�ݑ�d����H��{�R�	�(�n�|f �J��2^R���X�5b��Ȳ�J �Bq�q��{͛ �0 5� Ĥ��s����8�ꤖ\�"�}ݶ08�쫢F�������<_ %f�@N ���>�}w�u�x��8�}��[���P���޳���C��XS�o���0gg��I��&���]���������t��5�sE�N�y��|m��bD@����D_Ƈ
�-���\�Ժ��w���^h�+˛�Y�A�1\�s-;���o#�H
������(�"=�P�2�$	������Q�d&�;[��04xr0<D��ٵ��������-(���R� ��V���:��sE5���^��_�:�S�ujU�)��yJ��W�m]o�amj~d�ہq�k}�H�����J�>W(NxIg�Y��h��hδ�9���ddp����C�&��B��O��D�"&�r�_r���j�ب��L�F�J�̈��V2hq�G��G'.�e>n>�z�'[�WOf�QlC{��ɵB$���f@^�>���76�JE��"�l��]�;GV�!�i$s��R�px>S�]
菟�]M1n	[�<A;�a��Gn�s�?��U�w���S��R���["M�*N��[�>}QU&_�H����n�lJ����K��ky�� �)�h��lIt�"ͿF0�X��Fq�@~�	%,��w*���;�
�p�M�
Q� �A�8�-
�Mnxћ
ߞw��P!�b?�	�#Ap���4�g��Sr+>۩��`F�ʞgsk��E�i�����N"�������"�X��u^*:�|hȟ�i='�`y���=��hW�.����$�;�`��ݧ�{�;�oI�d%��QO��uޝ!ZU��&�%�h?�+�a�ν{�᪱���o��`Q�򨌒RҊ�)h��k�?G$<S�h+|.�\=d�2w]�ٮ��$d`d:��i  %��Z��YT�B�VaM�>i9y�#����2mQJ�����2i4{�(o����U�:�f��4�D�Qb���c�NE���[�w�0���Oc;ۤɿ�&�9�򛌶Pe�y<��{����u�V�k�DQɓ�T�����؂J�Z.�@6��\���O�Ҫ;ǿ�m�ڨi���]fN���?���p���E�R 	�n�4X�!	<�^��؂�냉�v�[�8[�1����������T�TN�(��K�g�V����]ַ��w���8S8$���֓�p0S&��bU��EU�s�vi,K_M1��8�Y�@�����*�w0�\^Fv)���ɓ�H�]�Z�h�X����rd�)�g5o�O�v,�%�3>o���y�������g��0��T�MS���䂃��W��U�D�����m�l!���}�eIt#g�4��j��H�;�/��h�%j~�Fy��B��[��h���aG�2������T�� E[�]�$'vkB�]��_q��}F��Ӎ���Ղ����
�n<�=}5�,����k,�#ql�ڭ�e��[�� ��KLo$g�D7J�~�� �D���, �&��h[�/R���0�r����O���F%1��]��;]F�l�Oi���s���2�����m:�_�)�/�Ϝ��/}�-�O��Β� U3kN��h�0!��5���̦
�	X�u�Gl]m�o��"t1��͢�3qx%���S����o�-6������̡���+��}�{��.\Rhk�ARr�1sD˱S욟֥�m�p|��ymĄ
w;S���&M���k��/I3��/����U�.,��_%���4�����_��s[Hǲl�.���O��;X�Ĺ�;��]�kޚ}����� ��_��5����U
�
��TA���%�U�w}���"�����q�
���[!r�]3�s<�A���δ���hb9&�1툷IuٸwS*���pT0ir`�{/�ؘK�Lnل�F2�%W����0��ue�Ω��Q^�ɫ�	���|o*Hlg��uFy��]D��Ʊ�j�E�zU�wt�ru�ת��s̼�\	q�� �`��M:{2;r����Crń��5JOg�*���#�O?�{1�Ҕ8\�<(�J<�	0sq��/-I�J�[.����L�f��j��W�Pm7$>w ���{�B
�1��)�ݻRi;}Þ#���.l83��̃
#��?��jn� 7��"׵�Nx��J�Xc,���&C2����� ��dM���gf���-�K��X�S"��JM_��0��ŋ���г�y���c��yk���7��S�h������Z�.�x�Ξ��o�H]�;U(^��3�Ϯ�y�
Sg���ܶ�O ��2��u�@i�Q�2��WEE\���8��B�DS�bJ<BDl����#�Dk��
�G��L��>�H���`� �J3�29T�� V�P�`i�*嶸p���4��Z�z�\{��S�Y�ƙ2ULB>�Q[��M��T�v�|t6S�V�׈gP	�,��aY��Ȇ�ԩXK$y'�E��N�1�h���ࢶ�}�tsC�6V���Q�;�Z�-���l�9��[��4���Ln�_�ӏ�[̃Ñ)�����B��a�H1�� ��L2�H>]���n>�j�ek�~一���󕐔�N$*�Β�
0���Ę (�&Y*y�yק�{�^be�������I�Ƈde�w�C)o�¨!�U9Z7�ɰxS�X�($��:f�r|����%37�<ڈ�F��a}��`��s� ��j��&V$����\:7�P�ϝM�}��a��JV3��frL5;֟:-"+ K:�
ʺ0�)�j��A-b�VΛ��
c��P�x�s�y��-~��Xg���������&
���*��Y�3#D��}�P>|��N޿�R���s��?
|�F��M�{�	 k/�ME,������e�d���&\B�g�Q3�^u�L�%���\��˪bɄ�7���o������!Ĝ&$iNt��r	⟠Ƈ[_�ğ�a�I{�Skp<����Q�oN\B?a���ݩ��f�.Q��JY1��f����Pɗ>������H,�ݘ��T�����ȕ���hdĭ��'�xNE��NC��h�4�_���	�g�n#��9<�fU��QT��'m�LMM�&��px��Ј���:]oG��x�S�޵�b���1ok������8t.N�%q����I�����}N�P��ajSϝ��ap}7���;�h���n=�C�t�����w��_��#�B�{�A7�%���kc�2\�"'�G�����9�F�C7��/��Ra6�
L
�M��rH�r�d�����6J��,E�XJ�p��˲X]�@7�N6;�AL��^�����4L R�G��ȼ��0�/��V�<�_	Ti��t	o�t����m[���}vp�a��wE��d x���X����p��j���s+!C\٘ݼ�%��qt�'.Zf���|j9�LE��kx��u����q��Y��zd�w�I�h�{7�,�/\�0V2�JNj;z�K�cR��M�#��ۏ�l��;��2��RwV��'��h�q�m�����re���a�^��S��㟜���ߎ�<qN�XN���eD��dp���$�6���#� '� �%$n-в~Z:��H� <c���ٍ�)�{�gH��g`�Ɂ
s���Ie�m��a4A���e�"���g�}N��ĳb�i�@��,�(�O�
��5h982RsA{�S�j{�����,l��f�DBR�9��P����Mj��G� ��	� 1����iIYb�H�U�8'·�j����mU*���m�
R6�]e�H�՚��Y�~#Kc@__p��H,S5T�=�K
���N�%�{�*$����G�D�_��S�5�ز�B�8�����i]hV�^2��;Z��nO��&�HD��	'�����+��Ɇ)�c��\�n ��}��>���ȧ�ڶ�X{���q(*�!�cl^$-N&4�; �2�c��U���x��.2���%��Ag�ӎ������mA��\�����]�J.BPEv��[��A��W�_�Ðڨ�Y�R�g�{�+�蟂���>?|��z�"{�A�Jus��&}u���W�����9������1����NV�0[Z�^��R�.L����P����(�m�,�9VWu.�4O�~���(��\H�]����)�7as7!u�����kT���urmv���aC�~~�c�)�෉���_�`cg��?��1��Sڴ�f���²ҏߏ#۸<̤����:a.}�W�J�Sũa�/��/`3�Y���k����f��.g	]Z��+�j `�=@�E��|�H�nP/���\�F�xC8۫�x�KG��lS3	
��;H��Pс���ތ%�8��j"�mܦYU
.��F@5���� ~�$�S?�Q�:Q�>KL�ĥ�ͫ@ҏO%c'.�d�.]O�[Ħ@��o-Q�FI��ݵ�{��Y�4!9 e�Z�&�2ؾ�BwD"Q��v�6��;�,�Q�Ŝ�F�;Q���߲H1�`��bb�<E��D-���c���+��7d�<��86�8s}�S�����]z��]̥U�q�"�r�^���~*b�.E��t��������i����σ�1�*B�t<�݊jw#t�i<�u�f���F��a�C�+��3�(�c���*&Aa��-n��^P�
���C�QD��E57H�i�<�::�~78 2jZ� �j�S���m!��h�z�(oHU��X@�^����nx��\SO�.;z����iJEߙ�؛'"�%���gq-,>��d���`K�s��Ӎ>��K �����)1�ꍟ���F��T��`!�Ҋr%f�TA�21�k9e�$�r�gi����k��<�=�@�Qv����OΞ�xൠP}��\��F�d$��2���u���=��s�4�_���|�������q2Y�HyG$�\Ol�eRpQ&�`��6�ks_��9`C�r���t�^�P��Ѽ�]�ߚp9�>� ��w��6ZE���(( �<Yu�.)���u���.+�=W��HȚ����()^��BP`�qx�^}�U����ɵ�TS��h]	��lax��AeD|2K[�L	�g\� ��p���U�Ӕ��#�R���Y�ggFf<;�P��L����Ձ�)�ɛ�'�]����@�_K��(&&
��8i ����XՁ�t�w�)����s���`�N��+7u�L�ޡD����s!D��$2;�����5P��vT��Z�D������_���oP��	�?��k�y L���*�?�ܱ!�0HC�\!�Oܟ��dM��Õb<��Pz���IިI��X�K����'r���h�c6�����|��R9�	�T���8{�M��
M��.����g�_���m�4H�	/b�t�n؃��X:.er���M�_*�z�aM�L"P�S����)w�m �%׮��6!z� �r�5��I��v���Tqo~D`��$hO�a�������i�D��c��KH��8�-�#�>�=�2%�#]�H��%���'�/G�@�2,i���1���_�|��YOc��&��L�� �Gd}�y��p�W%�p8�� �jz0:�D��e>q~��v�W�蔧�߹�ʭ�0�����ѠF���ȏH�|�mNP���O�8���L��͊�;��Vʝ�'ju\Dd8��뱴� Y]�ܳo؄�+�O%O���%���K¹�b��uV!�]��f# ȫ��\oU�#)#ѥ2v@�4�p+��"�5��] A�w��w.���Յ�t i��3�`�OW�(f����IY�OR��k��oe����r��t'79F<�Tۮ�˹�=�͵�����A� P��(O�*r�^u�6��g�+�/�2��no��D�RH�f��f,)?0�W�l�����2�fy�qU<"@\\�V�B���׸ך=���˾Y��@��<�E�~m�:8cV:d��H}��P�(���"�G>kJ�@��{�%��p��Y� ��u�"��KY�{oa���w:��ݟ�3�ب���j�������2�����w���ba��W���	N�r�iّ��>|�w_�>���0A�5], j6��6tD��A����>o6�k�-�r޷[6��̍O?V��b�ݡxYv��D-dG�H+E�F&�]�����:RF]����cA�;Ԗ��>�&?a�<1�[!}y>z���'X�1�n͔�ڦ"*�}Γ�JL���s��謻�Ӱ�k^�C���)z�Ҿ�����~1/�;O�Į��<�Z|��n�xKha�	)=���,��F�|��݅xg+뚱"�zN'�`C��=��릲~1�o\ =d{��QF�9���;�1��p�dWǄ�ό��L�*�A`k�O4���Da��̆��������{��϶xr�� Ch��u��(;��>���=�lY����ڮz� �AVG��"~��������0��ģ�]rj��2��\��ʄD��H�j�!G�9[Cpd7�d���Aיּf�Eo���˳	������CH0̓B���q�-�d��II�T=ŋ��� I�ṔKS>
���1bu\���%h��Wl��u	�:b��֫O�����/jw�� =�dC���|��q�>�9%�K�1Fm%���?w/�)o�D4PmX̒qdZ�I'��q�쫛a���d3#����Yqشo��8�)��l�N�<���K�)�����y��/��m�� N��N�����\λ��b�r�H�@�L�v�GA�U���atr��)VAW���#���<���fE�s{ m g[L��1����nK0�gs��3c/TF+¶�	�Bh-�Pؙ[s/k$\�H��guݲJ��H���Zr~ �Ǵ[J��^�Ƹ����0��=�Q��DJ�8O=�2�2غxw�Be'K���Ԑ�_@��9����X�y�"�%���� oZ��l��k�K���΂������2��q����9�6��]9��Z{/F�;C�ɢ7"����X�����7Y�Zg ;�i��Q$�m�Jpw����%���VJu����il�c�ߨ
��up���u,��3T�V�=���*f̏�d�q���,�]��׀����tt�䄵
+b��7��_��6e�=A����Ů֣�#�X�<��z�li	��}���pP�F��������|z������ N܍���W���e�o+��k������vc{�g����9�𒕑�Y�bgo@��s�H����R�v����脅�׃|�/�t��;��i_ƕ�5Ta��f'��A{�}���}��R�D�?]��?T�0�nS�	�čn*�b]_����mT�@�uZ4���ƕ��e���ۄvFQ.P�T�{)��?���Jl1��i�CҏL�a@�.��R4 p�9d(��6I7�U�5�I�}]g����̐�V�KR�`�_y`�w_qm���+ �|ElM=.��?�D3�߅�	��>�
�V�o�Y��믞����[]���\�Q@T�'ZY�pu�8i�F-[f\�	0��1wW���"���'��z䒣�x����(���S�� 
�)��Ǻ��F�4
w�E]�����MXYvw]��E+=�{t�TD�@��W�d�e��-3"��qj��}
�͑�b����e�ae�l"��'�羋�D��r��+�OK{�`lK5W��,�XE��ET��x��]L��~��c%_�fv!m�ď�_��9SK|Ǚ�W\�[�HE���s�p�'Qy���-(�;�VXEt
7��;C>��]���a�OЌ#���;�ًN�@��fZGX����qk�&]0�x��|��J|�-���@X���M�2�A�O�d���r���HB�-x��������<(p�Ξ	�<E�tf�lA������Ǆ�h�s���r�]R����vR����Kw�����럢[�8(�-��Yy  ����i��Ҫ�o��%��)�%�#>�U[H�43�~�0 �v��~�wI~� ,]
��d}�z�{�y�v��Wn�-]��3lv0��ͬټ�@W�G%.�e?ň��|k��k0��]�u	}���3�tugT5�cx���e��2��=+��k?�Ў�כ��\�a�c�bR��u���L�ὸ���ow�5m��-����?8��C�e>۶Nޑ�R�9:b(*��uk��7�'|i�L#�w�L���pq�ט[:����S���:J�a��S�>���YF9�{$�A4�G�I��cs���挤����)����>�j2�.� XBkQeE?ƿ��f�-�t�����TdpZ*�i�Yd�o�M^:�r�\\�+9����$&���W�i�I��Q�cxIs�	��N���7t��=�b9Zu�_��uw\U6���9�@襁�H��a�j{�c���}�p�\FQ ~i"����U���F��Y0�˺[B#j��x��k��Y0��:�0��^�������<����&�����
�`��U�\�^1��4�>%F
��O�_>X=���Y���xR�^N�8#[����;�O �Wޯӿ��R��e�ӟL�頔u��ӱ�T~�~j���E�C+٘}v�]���*�����}����D5HR2�+��\����5����s�`�3%7���N��:��1��e�BH�����:��Z&�V�k��#��YdKS���y�.���B覔����~���<�\AyOն�۰'ޱV�����r��y��7�qV���奒�@SvQx^il�ZW)h�q�{�y��2�I��-0C;Y�Yz��e]nHь8j��6Z��!����9;��8
��&������ѱ��~k�g<~~�
!Q�7(�m�	�[���*�w�]�����K;��"��95�z1�Ү]�0b�&���n 
��	_2�j�d�/9�H��(��?����e`2��_0zKZx'*B��Z0��uZ%�Il`C�)�ۇ��t���8ŗ�D�.�e����w!�ެ(��<?�b��ꆗQ��C�U��&�3�x�ܕ�1V~�����a9��y�сڙ�J��{��_?.kO�t�N�iBL�H�/�u�dB�|j/�@�Y�͚�W�����"!_�0BX��#j�26���e5�	��h-h�����<ͦ��c��I�#�(����Aɓ���e��J�U�6T3��H����9VD�F\�����l���y�)Ov߸B}Gp�d��* ā��r�@���d���+��t������D۸*�����Q��Ⅎ����/���Lũ��q\	�}y;�g��j���G�����1�vn.X;i>����p^q�Băk��МJ�e�y� �"��w��E�n��Np6޶2|������;��!:h7@��,p�Ğ��sD��R��_��OX9ů�G9�S�}�'�9V�yl�ߺ2�(/��:q[^��p����$�W����2�b�����i�Gc��?I�n��+:���m~Y���Bj_h[�8v��T@,�pWۦ��`/�B�+p�$Pc�Q�LN�n&���}R�ݜշ�,_��c��Q����Md��[�>����|'�Ѩ�C��\�A?X�)W<[�#�A�O�2�1'�������a�����t�j� d��� �� tIr��Ӝ�YۃPZ��=��x����8MiM��?�<���:�����z�}���slq8�)P`��թ*u$���!g�S�(��U���T(K�JL���0��7ţ�1y��wh�����&!�l�wg`�	ڛ����AO@C���ӣ-�78�`�Ho<n�<-�ʁ�8"������e*���p4*��Nc� ���^^��ql�aK���\޶>���{�8���3xt8]�%���߶c(>�Z�e�=�dQ�S�������K�����:j�wL����� �WWhnX�'��dSb�P��%fQl$������s����7��[]�E%�E���؟ܜ�)V�vr���}�cete��\�j�#�2E	��OM'�qE�������_i(����7zH�c�ɋ��6��QN��[�4��J�/n�� ��O�����U(F_N�8�^tdp�����P�U�Ĉ�k�M�ˬKe����6� W�ӝ �|�c<�nzi��ͽ�ܣ�{u����a���B�o�D�r�nD�l���"�@���7t�����n�ķp��f{�Wp�g�@��/���Y�.��*�O�=lk �k�ğ)�ٺ�E.� /Ɔ-8$P��� �;ҫL� ��6'ℙMya���W���w?)��Lw�8&N����g�1�K3���L�Ѿ>��33��OƟ	z�Ѐ>�V�豋�5��5�h���&�l���R���T�!*���'��\.�?�_����i������ �U��~���"�ƉҨ�`|�q){r�do�踌	~��+�����n�~����k*�^x���k��A��n��������y��OW26O�F��e�ă,�\�^��\L���A�#�/ے�Ir���%����,6-���>���[eܮ+Q�h<�n;c�4B�WO;�Px����X8)�k҄C_Y��������vZlS�8��H�x�Q�:��u?�\ȉ�4ޢ�+U~�@��'�|�Q|�ނ���s'��'�n�'�{���L��0����3�GZx��� ��]($�Zx~���r�FA�(q�Q�V)=��o�l����L�|B�n%o:�6��Vӭ��5 �Kz햨Ĺ�f�t���"��T���N!'fdx���2qN�K�H� ��Z�P���8mt�7C�4�!�/N͸E0���G���;FB>�C:�[J;X�J\���D�b�\�,�g��h�:E�?]������M���Vu�U��t�{���Zk���*I�7#��c#��Wc����$�S^%R�����m0kq��gpu;�؆ )B"6r�4�Ɓ�#Iߧ�n��cD�咁KґQ���H�D��^p�� ���G��<�g����f��	��d�z,I%���Z�jpI&�CC��+�
:�J��{ڳ�.P�m�(�lSFx�/��  ��_C��u5�O� t`�U��Ђv��a4:O=��7|b�_�6r� ���Hݹ[��б'U���I�*,��U�X~c��ٻlU^w�I���u��!�9F�I�q�RғU[�3���GV�?~�q��O�KmMT���*M�=njQ�Kyt��#����l��֩����Hau����Yur��,���e
PhF��r��r��u7�.m9<-�+
��ys,�;}���.��y|$E[F��+�P/�{58xacv`�T�4��_�}��us���'6]ns����j^߻���~[h׺Oې<���x3�0�"Ϯb�_�D��K��6�9�WNw>�>�����G��}�BE��w1� D�E��?���CQ�������Q�a���闎 ����