��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0����_���3�b�e�款ҽ�$�rWV�%E�/����z�XB�klL��z�7	Z�sx��	5p'��|�
&��I隆��!!ߤ�*fv�)�l}
6	0�V����(׿��f\ǕK�"�~�0�<�Zs%{���z��M��<�[q�;�NI���@�bp��3.�D �%$�_h	~+���F;t�o�[dVH���B ��\�2��mL�$�b�"0D��K~�\������L!cϓ��Ō~_��A��Zf��ű�H�\�[@5�>Z�^�"�� �O�s�v�+�ql�D��.�Uaџ��h
���8�h���"��I�HZ_W����ū��Ѳ�f������ԛ��?�6�<��x�d殳��� Y�	X�ʘ�7����*������l��V�:	�7�k�m<�҆��\88վ�C���ڿ��umT��4���9f$��4�i��J'i���Y噼�V؋p������O��q4��Av�
�[HKL{h��������U*UൃВ�c�.cW�ǡ�AlN�<�\]l�������Œ���a�%l��6�O�B�#�$d���"Y�����+	>؆d9�گ@_�Ѭ
Z�|\�WC6���B`ݳ�9�q�+�&=1#�C.�>(T��
.`�_0$;�Vn�NO�@�ka���U�u�[��Z_+�3�"Ϝ]P�����`��Z14��W�ǹD2�A�!S����%��wBKRwIVf�p��q*�g)�����T��K��i5Q3��}�I/����������Ϲ�����B��K�|��xNq$!���o)��/d�P����ղ��������L�*Y��f3+w�X��ݩՕ�;�:��md��)	�?u�b�g�J�N��R!_�C��D�3��Jp#�S֠�'�e�S��+5���0_ySLo ?\O˃d.�������ؗd�.��W��px��N0�)5�e��#8)�1I*˫�8GX�L"�1y�<N*Ւ�
!"��� N�w�6��NH�Cw����j��ǋ�ApED�B��_�=�O���¦�g�y�څ[��Z����i��=9�$���3�z�b��K��q���P�Zg��V��I��Y,@b�wYr��&�,�W]۲���ݜ�־X���������> �Z�c�@f.A	KV�e������F�V���h&��>3��>�b��A�\����.[=H�nŭ]�� ��*1 �"�_а�d�]�+���|�ʪ�[�f�Em✃���x|٤�W�,i1�0��c\�=t?�m?�g( ���MG��rj��Rí�E�XF�I���:�j����I�KQj��%��M��pF�x9��k.�o�ugT���i���$o��L�׻�c3����iu�Z�s��,�	�V�Gp@q��T�<�D��]��f�y�1�L7L
��Y�Y����O���}��7P���}�C8�vl�ݯ�8�\w�tk�}���Hs��rLm�����=&@ ��5���@oћN����9�i�G:�'�y�FD��9�\��OF�M�F5�Ԭ�ڗ��[Ĺ	��\���h7�����<�=���.C]�8g��V���ĺ�ҏ��E)�(n�Џ�8��}rh�|�Y���9���g	�NZ�o!�h��^�%���_߶Z��/�7����KO2�J��^t>����&PR#���R�B�"��Evt$�>Ro���no�VTz\EC@������`-��z-h�K�pAژga �E���Nş�W�1�=���C}�e9D�.���F0)��e>�����0�f�?=_@V��	��w�8RF�c�`=�ճ	�+�PNՃtT�'/ʠ�����u����[�Ʉ����?�H۩��'q��)��Q�?�|yE2��* 0f���G�o���n#���ݍ�u<X�?#싸�M4o�?Q"S��xR5�
S��!���TB������o*�j<}���t
n��<�	S�'�YK��N�¯�
�gV��@g�6��i�A��"�Bસ2������eѪ-����wV�r~�
��߃�G��s��+�Q�c�숵��݋y��?
-ˀq��5;iEh�T�.�u�����A���iP� ^hP5���l��~�zg��u:��k�
��ԕɝ%��[|�f5�l����e���Jxi��z3���4QUg��7b�Hiκ� �yz���2��A���T=���#ڂi�is��Ic8�pm�ĭL��ט/�D�c!��zzX}D$� �Y��Y=��G��ˉ�]�:�����r�YV}$v}?��-�2)�DI�_g47���ʾA:�O5^Mh/��Y��T��� C'X��eկ�Ë��t��oY�4G�qց�{zY�-:(��ib��[���T{z�,%H�.���Q_[b�y���
er�����YXuR�!kwn��~A�Scl�t�2^�@+��s�K@�1��W�C'�7ا�fV5�݇�P::^6h�\e�%�Ϛ0>	zF��!�=>�?���(�n��Z�6��P>��\:�&w�T��m��-1!2�K�>d_��}iOW�����h[^cʬ1F~h��q���Q�����eB��t���խD�T,��0]���������j�B��=�s�����Ȝu�s�w��_p�U�ޖ�6�/'�`�໩_@������S���X!N���fL�ʚj95v˱�AWo�m�1���#�7�8�V$J�P�i���f�P�8�@>�.
���U�n��++Z�]}x����;�-|�N؇Z��_$b{���/O��v�+�Ai��{�l���&��&Մp��s`)�!=��1����A2ʮ�!�n��J��s���35m���f�ǉmw�=R����{���!ݳ�,�1t�i�su���}�[�jA2��:��5�?NB�|�"��b+S��i�ҧ��"c{Ͻ�v �e*��\�7��ɜ���g5k����-m��H������r�����v�5���6�q؇�Aе#9�A.�Q���Ja��@�����G��� A2��7ݝ�q�8g;��?��>LT/�n�Fb�m���<��-������).I=<F�Mٴ����a����M�(�sP`��﫜�sA{��*w6�(J��2���
�d��̘�u*K��R-ᮻۏKD����KCg����O�/h"�%�D���:I� ь.�AV��e�(�����#��Wa�۪�7��B�^*~���@�tVx���MR�Ն���_w$1/����X T>���ݘ�s�S4�Y�cC�|�*W��l|�vĵ��x��f�?]1���e�����������;��kq
�Vlv�΂��0 �Ns��{y�U;
}9���Z�'-ǅQ��@�:y�c�������w�L��\ͭw��&o�Y2�py���T��^݅�.�\�H%>	QkHx�A���v�*���I�܌����P.�s<!����fӚ��ټ֚:��e��g\�.�+X��3Ҕ�D�^qW� �?i���Ib�إ(;�y�H����	k�ٻ�C�V`P���ֿ"L�U���+�����s�<��M)�ۼk� 9��LC<�#�ׁĶ�|*�>XH�?'D�!��걭�-V��A��S�Q�m�ű����j�����(e��љԟ�/`i:.���J=�����z+j���JȒp1�&���	w*\�f�s�|IU ��v�	!��"1],�����W�}�	΁��P�nvڻm�%Y���i8�J�d����bw^	�G`:��> �H�EC����d�a��K]���fU,'ߠ∛m�n�X դ{���?R�p�g�EFI��;���{}��,`��?���L���>y���d+�q�[��`Z�w9 >9��acE�EN�@/��h[�����D�Vƹ�߫���]�C��1�O�Q�3?1��D֕�G�P����0�GN�p;7��Y�jm ���4�!97��_(��>������Vw{+����-Ԑ#ŭ.�8"��H�T,�t�9#�A��m��T��|a��&�R{��ڳ�5SxO� ��q���D�'K�(�]��de���V�_*�d��Z�f�'�N@�hq�8��z��-���[x<��r�K�
��J~$P�;ց��;�)������~��C��4��By��[>�t�V�l�X�d�y-����+"��C�!O����p��g�:���5v�Lkv����"�I�JVX���3�	�S�����. w��3s�F�a�Q���y��
�f]^��@��{[4:AұF�����P�A����:4]�¬��;�~ϚPMCa�KӀWH�Hz�YŇ�f�Z���2������/��P�М�]�j����x�X<X���zz���D�)o���$�ۻa���[<98B=zt�_K�#��@
�C�V�숫�ܭ�㽈}���/3�5~:�[�T���q�>o�0�B*o�@�X����Z7����y��#�=Ag�%9�N�M�b�`Ti.���+�˸
[���$*�=����t� ��j͹N7��k!�����-7���v�7���7�f�x���ңfiЯ�§�xUAv#��7��l���m��^��g��~��₂l�̤=òy
���I8�^��q�{s��PJ��̨_��+��2er���>a	^݄P`������=GBE�-^M�H ;�1C���Ө���}�>��N�������w�{���|<�P"~iX�%�c9Y)��nǃ�����oޗ���I��G������gB,�q�<��&1Y��d��	?���A����9�E�.�k$[r�Ue�Nh�A4�oQ�$kN���ʺ�ܚ&���4����]����?��������ȁ�-��no�FHxnk4��mG��z�6��<Е��A��-жq=1ir^K��q����`�2I��FZ�	;JOw�u"^�"c�m�«�j� �Z�B�l4};�����U��������H&v R,��b�	�	.�B��"!*����^Uby��{���Mq����O��0'vu�&��q�*!K��������b645�X79�.E�t}2`]����	��)�6�GU.����#�x�+��a�f�ߡ�cŶ.��;�ɖj�j.Vk�мS~���6�mO��<✜�PR����Éߋ'�M�ؐ�pq��n��pj�� �v��B8YUG)<&��љ�1D�WMa^��Dl=tvVIv���B����}?��U�2MB�\�����a��@r�ȷ�������o�[��-[c��L���~��u�礊�VKb#��z��E ^�!��stDBgc�O�q�D�/��8e�q^Þ�̓����#�i�G\)�o���D8�>Xy��g�G\��m^���S_&��j�Ga����OJ��F��ر�{�<��b�֜YŲ(�+�$N|g[�")0��7����(JB����u�˜�@��t�n8W�.�jF��D���{�ŗ�*2�'�й�nC�{�^��c�qa놌������Ό¿��i	�჊'�m�F6Q��=���gɫv��?*�<��0&wwn8��c���WcΤP��8����+��2��9��Rw�S���T�ZI�e�p�xa��u/�Әd��i�ã¹�5�h�i���I|VT/~�h��\L�$��FB�6���������i9�k#Λ��\�M(j,�V��`$2ΐ�1O�.d���W����o�+�����d5�6��H�/�]�.F;t覂�.iyrdy�y��2����5�ӿvC��9�_��Bf�vm�@3����'.K�`���0��]�d�a��LS�/p��º,e�2D+Fr�a��������
eC�sA!8���2Y��>P6o�q:�
�׫�GsB�I��m���R�������Bp=����Y
�3_O��@�J'�(�)p�=��4�j�.�h��*]y'v�^��N����ڳ����e�ulܘ��y�9��������g�6�=��A�ǲC�L}�$�p�� 2��� I�)����I�/�*|��{z�R����_t���ia�tv��R�EQ켷�ʓS�>�.���KULs�y2�AD���俔������>����hj���``nKO���Xq�xV�m>m��ֽȼ��M %j�Lӣ;}��
��_h���\Z%�_e�����Y3EP14x��Ld=����-�O\���$�齧��}��lB���"��W�	�'��̣��CFe�!X�Qʈu.��6P�F�Y�F�j�Ϳ��F.݄��^{��g�۸ '���R�~�A=E�K�u`(�0m�G�i�|�P^5l�H��.��~B܂�.�����/,��d�I_K��� �T��O�)L��%N�xϕ�(�����<��ɑ�u��du������PR��QQl˾6�sz�1�+B��M`</	X�E�G���Ľ�%����T��d�~P﫨���n�0L�]�������_<x=��/Ol�|fa�!4�����41;y���К���Ǧ���0����7��U�%��_6���'SGg���pp�?�7�-�6>�'d�N�#��FK<~5�F$��O� -��܉R��I�@Li��t;��>��d�����GP�RjD���!t���u��Zi�_�x�֏�8oVb�V�ƿo�j���@\����-�G�J����n��[3!��V�����>�?���c����j���A	��c��V�U���Ah-ؘ;d�G3���ja:�>��SG�Op�<á��u֩��],����)�T[x+�[�o^>V��}O#xfN��ލ �V����q�U�߳�UK.&B����ͣ��0���ة1�����ȩ#�#�<��k��S;�2�o{E�I^��N
���`�����]��( �B�B��JȊ�YQv��"/�5��Ui�x���V����O��shѯ����o�% �{�34����ɍ�F�F��m����4�<&����_�9�R.;�����,�F�sۼ��F�O!����S��� �<��`n='��߆�g�:��B1�Y�B��dǨ-&>8~XZ"u
�1D��x�m����Jw�,���Fa�b�ǽ�8�4�H6���׸62�p�N]���k���X��-���2B���CaM��M#09��`���h��}B�=<����W�{`x",�b��j��ϯ��\``�Om��Y �6�q����� wm��@���&���qj4��k�H�=�T�27%�F�n�O�m��r�!|�� ����O�>��W���ABh�M��R���z#����{B½�{��)� *���z������!��I�=;�=WZ�AZ����h��Px�2\9��o2���Cav�*����|�@�Bk@��|�hD3я�6~��0̤Bl��N���'���������0=Gذ�O���ޓc�A����b�X���R�i֎�yܘD��v�L�k.�}dq�����Ƽ�q�hG}�9��C,���L���.(�߻�$嘞_1 ZTH}�^�D8�����]�9]��cj�;�BF.�7�#<>+�q����k	�JvCm���dG��dj���/��@�@�~V`��p�'>z���Tn5���C�鸼����9�LC����|Qj��|��N�b"���Dq�i��pE���|A��(=sen�G�+��R�V��N��=�&�(k �ҕ���7��'м����"�����K��))e'��GI*�/@6�8N�3B�o�u?�k�W��E�b���I��K?�P�`�Ґ���9t9��6c�_��\` ��e���9�#y���!I�h�|X ��xR��r�);��y��똵a�C����a#d
���wxU�F���=!�-�I86�PSN7P�.:)|��砙���ȟ1��&w"r�6�">����H�l�l��2e��_B�kƭ]������',��I;7��>�?=�%V���{����I��W�?@=������ �΃��Q�8R�m�\�ID���u�Mê�̕^�����W�� ��)-o�"f��u?��_���t��~��D� ��Bu�|����3��7�� D���-���TC���XfBXd[IH�	t̸o;ӈRG)������ql%����<0v��\aH
	�t5j�y�=��撎,?�>t��fx���D���O���P��Z���ĜK�|7�i���o�ұ�Q�9�e�^�E����5т벆�h}d�s'�e�߬Bܦk_�P�y/�~)����6\*Hg[��e���7�i��N�n���Dn9�.���n8���&&���<����{\����y�>v�zG��c��h�I5?�]pG`�'�>n��ֽ�+�6���� 3�,��pÙ,�q����s+ �I�y5	:�Ɏ������ǻs�V��EOr�W~�^ʇ�g�f«˄�"�;��YN�	�Kw���O�l3��	��@K_;y��,�fj�c�,pS;�T�|<�`2:�E!��m���O��9�Avnv�RVf��#bϪ>^����P�[���O�vJs`�3���X��ʇi4"TS�>�0�|fb�8�si�>Z{)�V�5�	�$�]ئ<@�I7�A���"	�f�`�Gj><�jL�;���T}��|�def��(Ee�"y���d�}�����S������mz&՛m�g/bQ��h�0~��ں���_$%X�XЪS���p+\���}z?T�R�FDq�-���4u'Z9m�%O���!z�O���H?���$" ܍����A7�ӶS���������a>eh��-��>��dp/Yy�:k11�L�d�P�O�����%�H��Z��]sd E
����i"�@�Gy������.b�>�ZJ��(�ܶ �Y18�Ԃx�
[�Fu�p��I׼�F���GY��,���`�h�HM�jS�%(7Ij�g�1����e�G�ʙ�,j�\b��������R�im?ɕ۷�d�ZmQ[���_�I�(�6Լ�ـ�4���3���Y����"��Ҁ��?��V[R����E˶;�!�$;饹������!JB+����H�Iɑ�3��h%�����=a�����0%����@0=�`��iɪO��o������y�j*��<�cFL9L�����L,�
��0�l<�I�H�_(!�DY�j�r]O�_���aజ	G���V�mO�SPM�Ą�}S������Vϟw�Z��,��63c������4 w�3_�1�Q6����v&��n�>N����A_���I����a�3��b,�56I�/��4Lɚvqam�Nuؒ����&����
De8C�^>�~J𰜟CEwtF@�3�W:�5�����,�j[�q�TcŌC�Mn#W��*���q�JYD!��rK>'�I�m[I���MT����	�+?��oޕs������I�xʺ��������ɹ���-�J�=\JKꐷ�Tgڰ�,@(�/wU����:�x�X� A@��}����Ay�y�@#����t�Q5�j���[lAezA9[��<�X?�%Y�q'�;VD���q��^ �T�������۶��*�E�[�k-V�pGO��r�f�9�o�����7��Vl&��dr�X�f�2L��ؠ�܃o�cgx�d�RY�C/U�t/�T����#� r*����#����������8�%�9)f�:(�V+�A�|�WN�.q�(����N��o�tv��!��f����q!��"#i0��4�5�}o$-�!�Kxe��~�w:���$�@��"���G �@�_?0�D�1�CK-�2�c�.����ъh ]qUM�J��m`^�By�8�3�,b}��)R�j�4޸Y��KG��+�WS��Gi�:�n:j<��u����.'�&v��,vSS�TR=�ZiW �����&�+)�U:=~�	�_?("�pV[���E|U�KB1�1iq�;����H�P���|4grP<��!���a��眸[:W-C�Q=����E���+F�1o�7�@���F�剨��i������5����_�"�#GK,��iUe~��#�4p��	b�����(���c��3d���7˘ˊYdV�:Լ��� 0�SlnuaBN�`��V"�E+w�Y���D �v��ʟ�4�
��I��d±��|�m����+�<�1�)I5�G7���$9S(�n�l�}��x�j/;9��gb��px�m�fܵsm������T�����bDp[NfKK���A6�yp�:5E�4%ݷ����;8n1����@��QD?Z�$�1��2a��dka�NE�Ť��.\8�RJ}�O���Y2�C�:&d��zQ�P[�Ȝ��~I�%$��g������o�P�����i"����"nM�_eo+H�]A��[o�EUQ���#�`yK��r�
�ã��A�܉���F��D������-����bg���q�S�R��t��CP��ͽ�@����B wm����grR+߰m��A�fB,���(O�Oԝ�?L��SܢN��Ť���m�l��w.	��Өh�yp#A��`�`�yc�|@x�����ͩ��+۴�Q��1����*��_&	|O����<^�ɢ]�tzKJ�`��W�eڋ?JKլ5�KԪ6�����hA�<�`a�˳UQ������������tp�ȟG�����d�O������v� �i��}�2�����vAuX6}�\��WPX!������}�AjQ�Ā]��ğ�S?���z�Fi��%��S!�WI���Ih�������Y�s�X����QҚ���9e�"��䱗�m��L�)nfZ-��[���D���s;�$�7��iv�H����[r��P@���]n�K�G5�>P�����������]��7)m~H�҅.����5���
霷���y
 ��؟~D傿4z��'|g�;#-b��A�yk�Q���*rS�U��z���&_�~G������2�o���4�Ŏ*2�&���]"qF=��Y>Ʊ���� <ڀzi��sq|��(������~�̽%�1z'�Λy*���u�?u\o�b�q��> ��\���l�zU1%@��6q�4.`� :������AwW
�k�R���f捇�^���F�����<���h�=k`����,���蓋,#P^�ڳM?e	\ٹcV�1�^�wtZ��8,c�5�\u�ޱ�O�s5�w��%<���\w������a�E� ��ޑ��Q1Ѫ�d��|��'�9ɞW��1!�B�%,���C[c���+��F�K(ؤ�P��J���qϸ�9[RL�h���eh!��.A��(@6}d�W�e�O��
�x,A!��AT7j��@�k��-�����Y2�2.�R*�AB��L�C�գ+�W��~��}"<�k�t��@7�q�X4s����ڋ,�t�B�O��f���:�`u�3�=�/Șl�o��],[�DQ�h���"r`M���#m�g���5�cO����O0�=K��39]Ց�b�Kt�����2��=�Fh��@Mm#���LȀݟЮ��*c�EN������Т>�F��Y�V��nh��6���P���N�W�b�*�D����L4_���}p%��,��jp
�ڡ/fתּ����&�&��V���r���~m��u}���A�=ز�K�?��/d�lgUKkS^�l`��"�u�*����Fۏ+��1�C��'�I��0Kb���mb�,��ql���U�J�"�P`v��=|�cP��R�V+U7$2|�*
�M���`��M��K���(�����8��I��*�[@�^T��xP{d�^�n	��lc[�ryE��˚�A�AՊd�3r��J�e�;&����R��7��QMli�S�?]	K||m�"7�;��\��ta$<T /�1�͗!��,\3[�Ƙ��p�ys��3�<��|�/���l�'��f�8�Q8��P$!�wč��@��
��MTդA��Y�6�alV��U7��k������2ԎE�X��j-��;\P����O;�Τ����Ę�`۽! a��}Z�
r���9Њ�u@����j��#n�u�Gͅ���<$�v7(�M�Tg����1�t���V �2i��\�U�)��,�������Sf��ڹZKBkη?gL�Қ���%�.[��j�ȉE'"In����g���.3��MZ�u	r�ɯ�#?�}�!A>8$�!�z�����@������v���+���,]�F�������aM�:�B�,x/,m������w��-s��O�g8薿yX�����vU�͗r�1��g���{��������D%~�����f�"N���c������"� �8PDDʗI�p�9����ѓy���o-�/���}��`X��W��iQ�Ii��<�I��R��;U^̆��ϖ��c����m�%6������~�N���3��=uFzP�;���O��N`s�ɴ|��Xϕ�޴T�ݘ�d���ʯ�ٔ���bC��0��X�/�X��������$+G�ע��ϩ��]�L�s�[�@kfI�d���C�GK�)0��<��4�Y����N�S0��a�Săeq�\�w�!Mm��"T��/�r+�|}�;�t���YB����T�WS��P�s�A�����j���;U���̲�0 �^����p��*(	�D��s�p\ΩD��/���� ������_���N���L��U��,�}�ʲ�Z�/cm�^�I�_��8^궈�3B�<��[��Z|�=Eߒ�,;	2Kc%�����'�6���<�-X���<�[�:��,]�y5���l��R4ɩ�D"E�Ŀd���0�x��q�<@T��#����* /��������>�s����'�xM�\�M�l����G�����*��Fs�q4�ӛ�UTe;%�ZU��A�97)₱S���!Ŏ������q;�d�eg�b%v�T�4A����e�=������im ��O?lzG�A!NX6J4Ѭy���RZ������g@�Ԝ|6�*�񣿷:����xނ���W�!ih�?�Kj�p��4���H�K@:���4ԫ�NϤo�T9�%جGV�k���r�ԕ~����k�)G3͠H��p �`��=\�E�M�+0�r^[�*ڑ�=�$��gʻ,s]�l�+�1�^��L~y�EGr��:�:u�y#c���:jf�]:��t���ڧY�!-��W�������<�kx�ɯ�,J��t�����uo��b��=�����G�s!{����.�1b�;��d���2���|�F�Ȓ2J�ĺ��at���/�կZ�M�j��)ka�()n;�Z�E*@0��ގ�����	��p�`G&�w��_�I2a�mI�:i�*�"��K2�C##��W`�p�T��]#6��A񂭡�&�fUQ/�
�qmyh�� 
��'����)�Vz�፶�dS��;I��AY��q�_#�0Ӕ���ӧ�>�g�{{�nJ�k*R:�3���uq�r7e��j7�`���c�=�7��$��~<
$�M*�F��o����<�4��*l��qI�`�����M�Ԣw(�Ñ<8�ŧo��`���dx��$Z�l_�T�G�G�]]Y�3�,T����˷��	M5v��;Z�eA�(���ѨbP^*�{X%F��y)IQ��}@��Ԃ�6�)�UHb~!3U];Ce%)GMk])������ő\Rm H����f����L��5�SP�rMGI��f$��+�Jj�iѯ���IFSg�S�B��?���V�E6(�!;��FVG$^�c�2������B��Sky��Z�<��c�Y>�����p ���`M~{�rד3#Uis2�a��4���^qLO��$Δ)��9")���T-�ӿ�zZ����8�+s�p��U�5Nް�5BP�x������~[~�H�ǭY�����P,*@/�o�ع��>���x����I�-(~�Ȓ���MŉG�^��; Y����J�=5�L�����|Y���07��K�+�
��<������^��d�ˉ=���&� ��pw�c��R��Β0b���̄��K�X���'���	Ё�n�H�i��+����J�8�����༚����ű3"ڕ��.�q��(�J���Ö�S�#m�_�6G�Mw�)
��ὡ�g���U�;]��٭�Iÿ�G|�U��1�@fz�;�׿�WCcUe�BB���d)�ef(c(�%곑�I�t�e,pb�Zn[8W�r��s1����gk␕� `���F����wo���r��&�P�Hjc�|乭�$���b���e��-&�{�̫��G
T�PU��Z�nЩ)��Ϸh_ݶ�:=��d_C��D���eii�LNKOZЋ��M5 f�Q��KW�S0��EL��:\�`qv�|j0�e�U��~���ۚN���0{�"�*�"�}�z��j�f�
+���y^�F��B�*c���5��B���e�C_D���E2s���:�4��͗����N�.F`�������������&�d�-�B�X1��@�ą�h�7�v�+�o���P�ؒ�!#Gh`��=������d!�"*�8�r^t|��%}p�yW�����p��H#����!*Gxs��O$���u2?�^�jpc�7��⛥3�q�m �vu�6K�^��^22��9�U���S���+En;I|�o=B���CBE�ݽ�@n�؛���DH�$��~_�&x-e&hI���&��Oy��܍�m���ۨ�� 33�rLʐ\�%<$=��9�[���
�$ "�*ejmKv��M
�T���^�CŞF�ExH�ѴM�".㗒,$@Ȗ���|�NOJS�x+�;80�Ǩ�i�h*��cQ�<|-]������
�<��β��Og=v]2�NO��Q�~����� �M2��^PB��>&뇊����>�Tμ�uV@�ۏ�F?�p7�z$�c�H�)h��<M�w,��wg#T?��Ȗz��ӻ����+L��5����:et�| ��}V���]˝0�1
���T깖(F��P˻��8�w�@�ev��%�qq3U5�EI�T�O]�
W��9�!�r��?�>
��իR��T��<�	�:>s8���Τ����c8����j v���tPbZ�$���'(!q�I$�7�G<��DL���Z�*�&z#w�	g#��WA��ʽ/I�&�K������� O�mf<�N��mJ����,��k��	�����!a��S����h�N+6���(�\��h�i���r��T�"����^J��k���g(+��eH�uE/�@r�-#V�5�4�v��ai��[�P��S������(x��r�1�(�݉;�Z��i����@iL�I"D, ����8������G�cW뎏�xL�K���>�W-�:�$��EQ��ڒ$q�f]//9j:�H�g��q�&�i3M[#��b�\�@��ZJ�0�5�<&�1�wE�cw]"/I3�Ȩ@4��{W���ec��t�����E����o��B6�G�=�ҺD�C�@�fq�Tcx�TA����<�D�ǌӟQz��ڦm(�7��>�ے�wnmᵓ���5��]��mI�_~�#����W$a�s�@��	�ޟ$�6�b���.בY2�ܯ��7�d�����B��0��Bo��r�I��,�����ÒT�9�������_������j:MF�EI*R���[�R��:fz!w4L"��j2ސ�4����ď�p�h�/�9c�Zs*pd'��E�PUy��e�.��¨wx� �(Z�gC������Gt�r�#ꇽ8��Ԙ��a��/�j=��C}*�~�#ФrOߏ5���~�ޚw�\�`%�͍Lo�����-_B�R�EhN�U���zezx�8���B�\%yJr�
7�YL��xX�����S�l�ʔ��Ə�S Q��"�
?�'uc�d�gD�/o)�����7�����ʄ#��(�X�K�L��!�b45�B�b	P�y�7D�yA8��Z��]M僋b�x��q[m�<^��!|��c�U�%�VOC��8"A��zw�������.@�͟al��jc	�:l1�W�	��MvT�W�H}�x�$?Ȭ db��I����Q>��,t{%[��-C�����9��]�srs�0�!�3�hn�s��F�\�+�Ji�i�Ԭ�R&@�a���_yX?%f��շ̀ǯ���@*�T�42Y�~�ApfEzwq��u\T)�/�W�^��<(|��Mwjh��0��2!�{5`����W�S]&�9W�.�nG������=����D}��[��ԧ�ݻ:P(hl�B��9�l��L��8O��c���ه�\�])��`�%�<�aKE�Y�b�cZ����mif�mȳ/�P[�z�&�A1��U�^�+�ڑ"4U�^�+4�8~�]�<&K30�]����#��V;�>��<7����Z?�m�gv�� �e44���d�!|��R���8�����jό �8$�ȉt\�9�O���ʺ��3�¿%6>F�Ga��$~|�O,�yd:;C؊�b#?�+�(�7��
���t��;,*1���g�Πw�O3{cС�`u6�=� `%Q	)�&����ڹ��%\F�����a�L}�{�s���F���	��Ea����)�yzOr���PwzR�<�s�z[�^i�Hg�r:���x�Y�}�tm�%P���MS"s���qJ�,ڜ��4p]�C���`AM���'�c�� } �־�m���Y��[WHy���X��=N�[ˆ��fxE�W�J�5\��<�{��Ɗ��3�	�����eS�1jc[���Q]�=��0�Ao���Vˊ�>����[j2y��Y�*�6��(va����%�j�K<T^�Ia�Fdn�+3��i�T�{�>���?�hH{���ƅZ[�:9m�zػʲ�n��k���붇3��r,�R(&fڈ��y���<n������vIЧ�Ѿ����m�5�e�9�ҽ�͉͆�=��K�8s���9�&�j��r}c�'I�~A��@,ב�#��"4V�JS��g�^ʒU6ui�N���R��Q~�b��#�Cq :�	�򤦋��)�jNn>�#���9=��������wG�s���4����y���Qa�LQ�8YIk^�F���`
Q�P���&�ʝ������@Y9l��G_��� A��(���y0������>uT�2qˋ�7/�w�[�@�ɼ��#���N�v����o7�i�C:�|E��c{�^DXm�;1i���8"���[XS�p��������oӰ�0м������S��"�����g7�o7?�-��jX��pb��,��,�ۣX\ɮ�5#gN�0��,#`����>��2�F-����~w���1V�
�(�
�����P{��ݞ�`�Z�	�|�vGr*��5�=L�@1}$Uڡ��e��erQ�j��vU"���Ct��wR٥�	��b̑��v�*�u)�*��Ԕl��d�:�΂��p����7�N�u~�3�� �&�T���/5P|�Q&�zQm����q)��D��io.�C��5�i�F���x�.�������?�ejy�Y�U�E�D���K�%7啀��|��ɿ"d�&���)��<V��H3�٠c�ׅ3���}�+J��u��tAέ+s�'FR�����	�m{S���v�#��ެ � c�A��u]u��K��>��}��#x�#�:�ƒi2��;�`[���'�ZdK�[������J)�#��7H����z%k�K
F���.r׼HF.��dAX��R��Ah�)*Sܞ x'��J�ΙS�z��mA��C˃E�VE#�٣��V��5Sz�$Ӣ�x�N{�@P��	���O�D�U�O��jj$��n��Z<�q���1:� h҈f�Ǎ�vcm����S�k0������1��B���K��[Wi��E�2���L֋�u�[7p��l�蒩 g`.�&g.e	��^ǳ|��甫��)E��3o ����撙lAɖ���r��
�0��t2��0)/ذ�9��->��ѥ=����}S�n�%��k�b���.>)F�fG3���jW���kC��X�5z��u����j�(>r�Op]�;1�%�=�!�0p�2�$�r�e*�(���Bب1Wad6Y�#I��ࣸ�?4��F@%Pi��K���]�8�s��MbI�sj�;��FW����O{|��7�B��c��f��g�L����(C�tNol�������w!��nv4ϾAL{P�����K���H�D�K6#� �l�����"�%����~&��f�� y��-�W�X������t}�QQ�\��BC���q=���"ʠ�Sn��˷G�Q�}�&��t1�A7�>V957A�S�k�H�����H�h�EIQ��p�}����d� �f�J��cLl|�ֆ}�"�:[�J�@��dek������_?�Þ8�i�+� �D�X��F�#�"w� S+K`�h��ȯi{�2�L�$w!�G�Ú̝�1��(�����F��� �}^XqBz�eM�r�y%�a���4���af�Q���pv��"ohf�#%-R̪�?rpc����
�G5��j����.x$Y���)�vI�,>����������O�:3�\= *0=���D�I/����z����t�23�o�Z6�f�f#����㧦����<+���x�7|+u���F�ݐ��̡ �,G$��Q{�k��z��\<���,%�H߫�Bk^'qZB"��r7J�di3�n1��n����#,A*��)�;�����L��g�,����v4�.`-<>2�w5`�b�� R��;n�ڙ�z�Խ��w�5˖��"�"��37�e+O:�j���\���C�Ƌ�6v^�pp��i�钖�j1��������=2~�����x���H>�eT������Z$#}�|�v��v��-�r'�6�G`}���aG��"g����~�o�V�岬����&d�-G������b�aŖQ��{|�o�ƒv�a}>[����e	B�?A����*y�|�;ȥ`�-r���of�&��]��O���V�9=���>�Ŝ�S�K�D�e�~e���
�y#�<�p��tۂ���*�g�tp¿-�o��+^���3V�t1����^z	 ��4�p��y+e���K@Ck�p_Q^P�$L�p�A��vw�e��>��bl�Rv����PPaNt"a�Jw��v��+K�����4ڥ���t��hDVݺ&rK�dJ�;KD�Ј�P˫�����B�y�.��K̊��CS0�wl3L�?��d�5¥y�C_n�*��o�{�?��q)41eM���N�*2���΍��4��!w�K����u�ȟsx��Ht��r_�Z���|�52���du��'A;����(�"@�Ƒ} ���<�@oX�*�h���m�,@�zh��xc4�+�E��[�0��<^��M`T$ª�T[��f3n��ϥ��<\MO��*Ұ�������N��H�j������6�M#���'���E����A��g��#Y+��֟�bO}��.�ؚ%��H�K&���oO���� v}���땲��QNl���oOO��7�.3IV��+!��E�)IsR���j�������v_/@&r�o�R3�f�f�i�r��=�R�Xy����ƌ�
��h�1�l���^wF�#����ݞp��i1���z,�����Qz���2��V=�e!Q�L��8%S�L��y�k@�����8����bpѻ��@L��6�m�$	3&1���Զ�VG���eI�D3X!�ֳ?V�Y]�vޫ�A��Uw�gʳ��N�l�b�-�nS�}�aB��?)����)���P쇬��X(i�>"&R�!��SRG"�<��i����E�����u��-t�1ў�[;H�R؂�Ѐ�1�� �����L񅷁j�s{���9v�a
?m����s�����۽P��Y���9/������>����z����w��9���۲Z�^�6Z�FjR�=���:[�ݶ4���ߢ�'K�)�I�1$�㌬�4P��HR��ʊ�y���Y:��c-|�o�p� �$;
��X�����Q13�5)�c�E/����h�~���5�����bN�S�f/C�Y!tI��E��G���u`u\8�%`��3)����q�}U)��7������$;��kڒg��k4��:\�� @ua��r�`�����w׹����an�����
ދ��;Vّ@l+-8��&���\�>]�>$
g��ƺ�T}�kD[,��/�����<W4a��R�����?nh���d{��G�&
�	8Bև4w-0QC����2W6v��U�;��<r�@}��'�C��}�����B�%�Zo���&~G
�uU���&trl�u@��pW5���߰��/"�G�O��*���lr�Ù>E��#

ǡ��Q]���uz��q��A�/?��uz��cY�W6E�@���qob��#�R���	�}tVRct�L���ʭDv*1�[�!2��`��^w2�^�wqΖv�n!̒��%]�E�g*rs��+��,[I��d�۱0B���c	ݪ��9��~���n��km�I���e�dc�<�G�Z ��@b?F�s!h�j�m2�\PG�Ft���3n}��VXT�Ϳ{���b�W��qp�0�_����`q.�%��Vw��-�U��t�)��?0_V���
��}�������Ra�i0��J������=p�[��f�hlU+�c:���;w�=���m�yeW�����1* 9������ɜ��/��O�	�w��*�sJ�M�h�U˞��8�G��6�x 3?�P�r��SA�aq$Ns�C�W.��[I�/$w�p�rP�sSzjwp�竌.p�]z2�	n���~jw�L�;�O�%�3���wA�I�m/�Zt1�j�\w�\��ѽ����	@�8F70C��
tϚ�Dl��؅�����<ꡓ�T��D����9�6�U��D%%wnJ�(�$�=$�@�ۥ�Q
���+��F�e�/����E8�A��$�dބb��ARN;\~�;E�
�O����������������)\�V|�J܊g��ĂS*mA�GJ8�&���|�����H�of+����mL:�k�V�C�g-���f�}�o�l�Kإmm�,��8��A��6��RQN+`�g��q 3��(��]Cw �����7��d�z�/a8.�=P��_��Լ"� ��.�*m6�� p��DZ<w|�s,cٍ�����
5S����r��x�C�������[n�����P��b��&Tx�F1`��H�2'�g��)K�B'�*�_�K��~���,<}��Ip�W�Q�\am/Q�Q�Q��R�2gx�! �\���eb�ŰU�Qg�D��Ws����]&�������&!�����J`��4d��yQOŌ
"�G=B�c�d��M�ІT�X%u�tJ��a��t�M����0�t79L�Ż0f�S�<�NRe�͑>�s�:`x���$��o��:_%�'r�(��cs��=՘��z��&�d�t��VD=u����|�;.`3��<�c����i{6*E�"Ё��f,$�ī�g�;��i%M1}t��-�fx�c����0�	��IjڳW���_~�rM��6��p�g,���L�Ad��9M�/��O �u�<�B�L�dN ���Oc��ȋ�9h��Y�<����z���� "�n�(�n�<�
]���j�΀)���h!���ע)]��Y���"+0ٜ������=��7�KϠE��X��W���L��P���Ƨ����7���r`ưd�1��G�|�m�X��,���]�0u�T�o�j�%ZC��<h)���\{��0U'x5^�β-|I��]��4Y����U��}��#����J0����F"e|�W����B-�w�J��N�������"QMȍ��e*���'ѾH
^���j᧸��� 7�#�t��s�}�*���  N%�Y��q��`iv�$x�9��� ��:9Z��F{���=�p��e����[��V�^��M	d��u�k2J�P5���"���h��c~�kje����z*���GMp��?uj���46�x���P�thVdo��+z B�H�#���W�Kq�cy�f��cE:�E����c"�����̤��(ۋ�$d���R�I�4���H����H��!�$��F�B�����,5Y���au���������2D+�Z6cc��O4��6����Зe�)� �<���\ ���J8zW�։_���\��}?�*!�	*�+��5.V��C��k�T���쀤t`�ð��6�!}bt� �\��:
�a�QB��#�*ϋtf&���?�n�����O��}ɐ�w��S�BX��G�o�e��3(��.���١:�v�ޮ:i,+�O������ۿ�e"�ˎ.�݉,B�(�Li}��������ժXź�q���P�'9���<��*�`zF�4�T�
$'���W��J+8T-��'���_Ǐ���{Ё���u��-&����l&�	����6Q�H�gn��C�Ώ,�z�r8}�*�랛�?M���):�LG��s̮�miB.�r`�[ېbOP*Ev������x��R��'�x]/u�����î���+V���zG9�$?F�F�@(��H iM��`�Gi��DK���7���2?�F@��P�	ф�`og̉�:�"�q���C�.1B;�eQ�:��Wy��N���)�JW�! �'/���$���
φP?�����>��b-	�p11�+o�@y=��"������O�\�CV���>�ώ��8P
u�t�%��D���xD���4�Q�P����p������A�f�l���:A�Ԯ9%��1?�������N����$�)&�k�cl�	����K緣y������۠�^0�۰uߴ�U|��R�7D�#���F1 ���T�Il�����-+;*�#�x�"��H��j��-�j��*y8_�^<R�!E���X����~�VѸ�u��n5�|�%#���~	/�N@�5I�X�k���}
�T��;u=�d���]V���a�/�RS��>f=i)ቓ�v�k$�bK�?�IQ���5�%z��S�ȕ��
��>(���-9Z�X����*�񗟓��!!"�sȿ���%%�'#��4hZ�ꢓ$gx��xb��A"�N��_�m(���4-���P�[��	x�t��_>����}ŀ�Ō��%j�*}��	���xi�g���!�/�o�
�#�xY��Y3㳠��g! |��Tr'�&}d@Ǔ��R�lnN���P�>�:l�^'2�zu3��)��[-����&Y�Hԡf�;�������}1�ڃ�=�����.�aW�����]~�M)!�Dn����M^�&�4�Z�1��
��_�R����DQ���UL������N�����o�N�/h���� �.�H�2�5�U�8�IE���������
�x��W�G߀*�p�ߝ�f��;���G{��3?��A�����F��y�6/f�ו��kJ�L��o蹷�.1�
�0�J㡃i"Pc�Oi�����B̕�Q �(4&�� �� �L92A�Kn?����b�D�����ӗ�kT}٤��� |P�h�`7-�.���9��ح���;d�[)dʹ�/O��O�;7�\�qހ%q���/�;�E��H���-N}�����&�æTٻ��@s����v�V�l�D1C��o����M*�e�i%��1��V������V����X�b��3^��~�S(�����.�u��=� ��k�֫�4x�Fi��/{�Y^�τd��4���_�OT��-�ic"�@��&����u�H���Y6V4�]�d�I6[���(|+
���	-���YEt�̝��U	\Zc�����Yp̰.�c��]�v�u
��l2�Vm�w]���^M������y�=@��F��Km-WԧV��ٷ���W�o�pA�P4�1�W#�cm�4q�:W��ˋ�ڃ]Lo�`�f`��k�+;�m�y�M�4��u�Q���8�`a}u`9�q���Tw���^�o����TbTdO��Q�H�ޞ���Hz|��G����w��e�n���#�Ia�q�*�����ݶQYc�(j�:Ϭ�pN&�%�(��G�" �{�&P�˅ܒa���6y��}Ŝ*�	��fB�AE~�L�.J�.lwG�ǮmcO���$�&�P�+:Z�a�f���k��ђ�Y�_{�4��
x�����'��4g<��&3�d�1djl�|�/e��'y�v-�BQ@��X/�����\=IO�aWFȍ��YDH`�w�x����M��6���}P����ڣ��!��}d�\mJ���Dߝ��$
c����Ω#�Cy����~��,a��J�T:�%v���!���Enqa��d� �9'	x+S3#p�KP��@�;ߎ"ټW"�����&G��A��������I�X]��R�*P�/�E��Ԣ��-�Bl�_��B�BYn}�74VÔ���g�m*�g�����<�D�;�L1�>A���"���3?�G� 0@�ĝ9�b|Er� 9W�w<�3w�B?��l�Ύ?�=ѿ;_nϠ�b�R�z�_#�^�C� 	!6�k(���U��ՠLTGp��#�s���H��'K���~֕�Q���Qԛx��@���8������^���{M��ܖ�ϙ$3<��$�S�v�m�W#��$���u��tW�����PHnv �_CY��ܺ��Ōv$�:���{�)�����:C�m���-ּ�)&*8%����aGh$#p9~�l��b�c�J@H�F��r`�G��?^�v�.�^x&S	��;E��I%�Y��F��!�q���h<��al{���J��g�u��;�Q����5�9Y������"���ࣇ�'��*7*+����&�r��R�ny�9F^[)�_+�T�^1��i6j��Qc\�Ɓ��Y-���%�M�D7��
�QG>n��N�p�z!�ͼ��'G���(�#km�r;����}$zTdF��BuEq��P�&��}�con�A���|�|91ʴc���w�0�ތ�����R�ZLW�<q��.�D�(��؛����mML�d��&���w|/V�#X
3�7�� H>�nB���\
F��=���P�N�?SI[�'����8�,�m�m��04>��|�׋�{�9�l� ��.�sx�R%�[�^���[`���P�\b������j�a.�x�a�1���S�򙍸d6 [�v}��j:=$�_\F��>��>��xޜW�ܿ���6UX����O[����m#�G)u�睤jc4q��q���7�r(�Er嚜O�xĊ���&�$��/=��/�sUo�;ǋr�2�fK��O� D��F�&����T�51&�p��;+F)(
P���S} ���;�$J�]P�.҇Z�x_�A^���� b�F5�)3In���V�啔	"x��~��eJ��,���t�Zfh��E_c��-}N�*\C��u��G�ĩL\N��j�`����T}"(�=�cf���x
��/4;���N5V�!�
�K��O��ܹ�t&Cۃ��<�Wϓǝ��s�w�"��݇��k������FR	�䍂�c��6M�ı���3�7Z�?,g����<��?;�<׋�Cy�?�O�W�Ygi.�F���$��3v6@���M��萰܏����=}�����E�6AdYb��GX�Ձ�A���W~{��V?�*`\0�����o�򣂅���酉�J�v��GY0�]��7a�7�Je+�lYp��&CF���~�!L�T���8�`����;�������ؼ�.�V �㲅5�e��%��K�7,��,J�=��np)�����F����Y2�p�~E�h!5(��sMZâkm�/[���P �����#��i�:�+:��C���2��ӷ.7��?B��NK�j��͞ʲ�W�G0����v)�4��Ew�����Q&eQ�Z�'��u�"wj��`��k����3s�������Lg��6��qitq��{�`E�_tʔ�<��HwT*||z3t�Q&)���E	n�O�[l� �d��f^^mrbF��U�����ܗ:��y#��sGͬk��?������4~$ܐԊ9F�1��z@��qLoE�IbJ|L�]nBКV�s;Y��v�xз����`���m�f�q��H��9��D���3����}�^�e�g�-jߤ�'�*�v�>H�BE�Di�'O�q9JJ~�s��� �����ʼT�'<I�7��r�����?/�GE��:`"9��J=QIN�@���%08�m�	Qo6����O3G�ɧG�4M#�5.e7R4ͦG{Aڀf �:k=+[�:=q'����<��q��-�C'��Gq
�j/L����{$��v�k.�v�k9y�+�h~��ٹ% �dE�����A>�TD6w���s��k�^/���c�ȤuL�٘�`�/C�޶Y�	_s�J����f��(�A��@�3
W��]���~=�?��}	����V}�}�bP{�K���\eā�݇�h~����u�ߙ9	M\H�B��(�"RLl
�-uc�Ӂ�v6�u&J��v2'���x*2D᪏yȹ��\ �L�\�2�C��1��w]c�Η�v�
�!�+c)�1���v}��ݣ�q�i�%^,\ʖ��F=^�)�xi�Ȅ&hc|t^�ӣ��I�4�@��S���$���w���o(OW���7�T�3ܧm���o�p�8p\�5���U��t�2�%vҨ��Ԓ��WQ�%��
�v� ��=X9 4�'3p=Apg<e��w�y>^����r��S � |�X����Z����b/qF�/���㱢�'������qe$���WNG�N��ʐ�ןY#Ǻpĳ��� E`E�2����Y�-��5-q�{��5-�n���x�$��H�m'��#�uq�?!a8� y�@��Ă�̕�1F ;�C�X�]�S.�םG�KA�%k�ӿ�u��Y~���c�%�0p�Vܪ���5;�g.�J0��*	���x����`6fQ��5z�8[!}S���wni'sewT��Q6��	��UV��ݮ<�~���3��U�^�MO<\��f2<��M�P`4��#_}z7������CrO�h��(0ǄF.�$��Β���h̅i�}5f��$�t����*b�� +h<���y=ճ�� K�'/����L�oQ:��.�5u�����r���$Oa���FTS�<8H%KW�qd�)��E���YQ1��)�S����]�0
+�ס�[o��^�535n
��p��8;�0�-�CK��Ƈ�|����w����%rT0�̡��&e��H�8�Q��ps���w�����-�5�l��������1
N@zK�v	��r%��P_�]��l�7A�`) .�2���Y&PDtz>^H���p�ٻs�*�!K@�Đ���=�ߙ}�w�%�?A"Di�9`r͏ ��ْV7��R����5�0d_���Ha�?W�7ך��%-���$��d�SG�q�xj�ԗ<�������Vxu��@*�P?���'�˟�6z��2�Y�32�iy�|���we٬)߬.��ׁ}S8 hO���8��2s�־Ay��9�(���u
��Q_�W��l��4꼚*��3`-�,ɠv�C�n�a��`���z�UQ
B�F�7}#n�e��k�҅ qu4�f��&���ן� ĶDq<f�M��
��;X��Mʽ-H��`�<�����|O�-sU�(:0GXk ���I�=�~�d��1Gf��);�-^�+ڐX��=4O�]��+c>ݏ>�)�Ţ�	$��0��z7��StC`�/����l���bvS��]|���i��Y���FPZ���kW� ���V�U*�-e��P]��B��c���TQ.ǭ�ճN�ǹ�����R���-��0|-��������k����TOi���m�P�
�Y�6 �{~
B�9�6���x����o�`2��U_ljz_�i��@���#O�"�����I�{�a��l:{��?�&�H; ����Sɺ����ٲ�9�͡[a�ˈ4?]�W�U��{	.��!�K��J�4�	[L�����W>Q+��w�B,%���L�pWW��iV�4����a5P&vy�[��WS^v�]��g|��U	ֲ9��о��-���=)	�5�ڭ)����)�Y�Q��xR/�T,b�W�pJ��\������T��;#��{�tNT��u9M}���)l��H�hfw����8�D͈��k�
;m�"b��_����!�+{�)`�<�iQ�������:m�����ϰi.��G�g:�- Z��c��C��?2I��=��v�掰�m����07��Z[n��5c(���ֱ\{l����:���/�H�>����2���T:���X��Ӂ��� N7P�����)8-*ù��IB���=�ǩ]}/���RU�.�� }}�#�$)��6h�fx��t%LD���6w&��4�3���궫&  DNc"b&��`[YD����a�Ȇ�C�V�m�:���%�2�L���}3��s{|k�F�f	���R�5V$����&�$� �A2�%��OȨ2�j�~�.�L��z��[�@��K= ���������6��h�A;r��(^A��.?Y�����,%/؁6
�m����.dv��W.�>%ӻ��}��G&�!���W��T��{	H����N���������qD9�]L�����{) q�Ҏ���4�*�UB�r@�����b}�&�A�Jɣ��S�Z^����P�������T�|�¬x�¡�����f_�j�Q��Ӝ�{�dޙ�-b�$���J|����̣�a���_A�*����8�AϽ�e)�~�C�?M��^������vNi��o�o2P?�%ZLB�X'��6:��uě��7�����]�:$�P9Avs��nR�e�A 6w%X��B�-�E���$f��ħ�9�h��ǈ5�� �� ��sA�MEŏ��X��5i��:%�r�Y���?^R�]S�j��k����E��	aN���jʸ��G*��I���DZ�
�p��b�S4p�$Ⱦ��Z���
�<D8���8(��۰��������ۻ��p:���v����(��,�ahCQG�ϸ[���_z|^�t�k��c�{�%~��l�#����`҈θp��8�vS�Ǒ�a*v��<%8`h&e���7?����]ۚ��8�_�{�/�*w_������� �	�[T��_�f��^�����Mv{����,���?��} \��WѤ.`Ё�cs�x����-�ӻ��Y`NLlǋ~�K-�M�59���TB@������k��7��ng�}�h��;�2�`b���k ��#�x���[Ȣ������.���f�V̡����s��5�T���3}� �W�J���1�>����hH]��PnrED�-_븬��b��?-u�����*X �y�B�E5�˧�ϣj���<gy�N�#���^6��
r$0�3��*ׯ�L�����8W��;��G�k2%5�f�jH(d29S[l	ˢe`*��[*� ���:C?�BU�#\>����ZBf��c
�m]7�-�P#�w��-G��Sб6y��Pj�-J*S�K�jhqy�?�(��
h����^(O�WR�{Y�/!�ق'�E�ʬW�5P�}����#m]�aMѩ�}���^'泑��"�[˲�p�U=o0��Q�w��8�/��kB��:�,��"숄�s�g���T�3�!%�ξy�e�n�q(�+PC�R���xk��W�D݋M�Y�p�E�T��Q>C'�$�x�o���s"V�0��|8��1�bW�!�"y��3��(�6��;_c��Qw�fex�4���4�������T��r��`s\]b�Ǘ�Xf�� ���)�̗�������<2��\����KE.��컗)��:k&�̯Pv�W�:�l]�ف�쑿���5��I���4�~��O�xha1M�e�fz���t���=���H�l�&C�o%Y��|>�"e7�XQ2�v�X�d�%!���d�5�;Z�Eb슄	#�������ou���2Cmeԃ���9�! /��޹�f�Y$�u�F�[A�`�5rgm,H�L-:s�}2���a�sS���>������D��i]-�y�0cʹ��?��װ��Juӭ��1��VQ��8)�4"�2a����?|ֆ����	�\b�ڏ$}vzE��͗���ss��k�*<�q@����U����Hf���\�-k���z$�6���+�տq�d&��9�/��yo^ ���5�M�x��I���;�¢��Wʇ7�v����-�jp ���S����__$eh�4�M+��iF�}�2��$ݩ�<�G���<�ˢ��*^ �)�bta���������c:3�.����S��d��tF����г�ݙ�� 2�]������B<Wj�<jR������_���r.��q.M�tɆ�5)�� d����C:�P_���L�E@ER �3�R�ڒH�D,BQ�&��űjO������/{�ϙ\���qK���']���1���Z����eC^�r�;���[�$=.�l���7�6Бѐ��A��0o�o/=�G��OY�e�_�ˏ�완����&;�k��,����E���v��Ƶ��iN����~�ƯzoV�-�ܥx���Hr̋�W������]k��P�ws���U���km��9-��ac}�o�V;�6R��.F�F���5�ue](-E'F��"�s�����k!Å -UR�d.5e��x
Q�K�h �۳���lcY�����N����ߜ�b���1��|Dʨ�]uK���梈'O;��Ozk���n~������r\�[ln�"�1-��j*Q�	��p:��~6��)���#/���^���N-�j"�q�y�q�U�"��Ewi�t��s�2s�-���5m�&x��]�I�6M��������ŌU����M[f� +������{�j_=� l}�(j�>q�����}ʑP�X��I6 ڏ���nԢjc�:���$�~��V�]A�-�,V+�zMi����
kB�ڇ�2w�,�a�Jb�շ}N4�%b1GeҽΒ>dS�����HQ�)���"�(E�u>�?�ۀ�4yb܄~�wegl`p��q���ȟOvz��yB�`D�ǗJ�͝]89V�;���	�K��Š�+�7<�Em�0�{.e4��R�U�D�&�Q������^8��Q��BA*��6J7��U+_כ�\'ܷ_��?X;'�����!�@�R����E����x�lc���;�*�����̍�� )W"��e[��,A�L�I:5�î٧���*�́�ܢ��]*(�ʟs�!1's]L�Q��?8���V�}����,���}7�a9��ajK��eַgl���m��,��tZ9D���k�`+�w�����;�Ɔr-`'O�#��V��+0���j��U��S��%F�MPW;�͑�o�y�V�'=��Q�}d�u�S�����j�8�3�lA���%�p�����nl��z���! �-��_�a��$�����I,���K��IK<�Xix*��?�������!�i�<������/y��wS�`eB�����VK��F)]ot�����
*��+�CV0mx��V��á,�f����h�!U�}��g����!�D��m��������
�;��nb�[P�k���fA7�)�m��i�oj����?�m�L��b=�_� ��b�X��Oى+��*?���#I�1��唨��eyk7��]��L���?���|��z��G�mTAJ���_�����O��xR�9tǑ\�_�
0����	�l+Jt�H���9�F�%e����~���E�jTw�4�3|�A���4y�_�]:}s�
� �sC����v|������-������PTT�;��-���d����G��n�ߓ㔝�μ^���
G�p����Y��L$'�1����ރ�2�d�uU�Ix�`���Ƌ�/$� ��\��)����)����+�3�@�uBrd������|����+��*���o��Q?�h@~|2_���ʭ"��wƃ�@�K�RXq���r���I�3� �dWP��c֞r�;�ؒ���D<ǃ������R��L�i@�<��zV*��r��̕�3�GB�р1�'ә��$4�H�C��R�0���FX@Bwj��"B�A��#�r�XW�BS��ȯ�
I�fz�7gD�e���������}��X`ݒVX!����m�^�3�ep*��x	��C�s��ݮ�뵷CA���ӟ����%���P������������8�c�c�W�^%��W�S�ĭ�=�!��#��!5A�m�yӓ3\9���`�͂h��u����=W�KF���c���gҧ�)�5��b����e�mT�Z3臊ѳ�m�Ẅ́M9R�����jC�U}g�YP�i�{�(�C�B�3�?%0=t�H�Ƙ�	��>ɤ�t���"��O�]�$���1%u�r�Ƌ���iJ��8S�ǖ���_�)�b��qs���f�v��I��E {�SX_ӯ�s�+����yd��С͆��MQ@���U�N�]�OH�9u������M<}!��򀦑�+�� ���fL�y�����`��V�\���Md\���@�N2�8�ͥHQ �RoY%�֊�����c��
g�
��Mr�.ʣ�=Eq��u�~Z[��ds�L�Q�X�h+jAy�?��WG@Pd�5-3���\�V���_���nx�ዣ��0���Bo�c���S���eFEڰ����.
e<4I	�_�n�hr^�Օz�L�}��=�0���&6"V�ZB.�. .E��十jbh^؅��{��jwL�T�tQ��3G�}(RNT<��к���B�@����
���6,!��Ӵ~A��FFO	�T�&q�Q�T��aO�Dx����@b��}���=��X�';��s����E1ǛG�J!���~L��@����d|��*a�/'m�!�dJ~���q��{�d^�Y��|s�3B�L%��gE�3f4�ZT3>�͔\�2�L��:�
�P��L��x�\�^��`�)�J��$�oI�bG�)]d{�+�W;�g,�[� \����:6�()βr^Lٵ�!S�գ�����}t�s�I@0��H�g�_�Z��a��c�'{!5C"8�f������2�:�`�p2�._2���?�x���A��sE�p%����͵$ӻ�S��}I�;�Q�(��'Ҿ���]ԣ,�e�Jit�F���w��y����\)ό��"2�\͈�T�OR���	�T��qy|���b'�b#�9��><��C5���QQ�;��1��mO��w�F;쑠��&�٬��?5<����%��
vN}3��S���KN��?��6���w*\VR�<���ޡ��D�z�i'�/T��+ۧ�4:�Dr���<aR<I�_Ś�ÍCz#��>Z�EÑ�K-���9�(t�Ӻ�[��j��ǂ��e�Ҁ?ewZ�:�p���m)�3��\0��Yݗ�w�(��/��������Ո���="�ș�i���<FzUfm�m�WA�t;U���K���Ϛ�.A�~��X�b��;�@�e�������#�?�w� �'��'y\������HQ{I�G�ȋĺ�M����v[P�>�ȟƤ���zxo��*��S-w�㈵�r��?�iЃ��n���2�w�\�ʫ�E�ST��(�JIm��\D�py&m�#Z2���kh�E�� x���J�.i{b�ܾ��f�qD<��	�gtȡ��I���'�K�V��ۉ��W8�,e��'@��Z�xW4[�<��6�C���j�oK�H��"���k������c�1�Fn`1bg��@�����lDQ�/�u�N����7\�����^�[���_[t����4�A���ZT谋�a`����"wo��(����A��GA/������J��6�ۉ�D+�1iLx���\�,�k��K���ɲO�4U:i��6��#��(�6eP�bu��&M�eb�G�Ӈ�!`����2���䃍�4�S�Ly<�5�˽���پ��!heB���|����x	�^��vP6�;�A�0E&�m7����=�Đ���VT&ҷ��uŠ�=2a�;n�I�
a]�EɈD_!H�{��mZ�~4��#I��75K��`k��P��]�X1N>���Z���ϜR+UU���T�D�,E������^�hk�c=�̽�J��ڻ����Eu���u�Y�5p�M ���N��T 9�u��+�So��ŭ�W��%��?��s���$�)C����m,���N�/�sd�g3�|��#E.���τ��f�`��
���L�7�%�}�D���T���x�q�\搞�Y��[�̙�PН��$p|n�b�v�mh3�u����ϧ�,�����-���[=uO��YK�Ak�j7��,�H5���ņS_�g��@>~s6��8�<����z�7��|""�u��n�L��¤ǞO��a����l�%����~H�KlXY\�XeG&^�-�D�.�r��|K��!�.���2b�$���}Zvv
p_����{�Y�����v�s\��t����cƏ,��m,lc�r���pC.g ��QϮ1cұSC���%B��Z��M����|f�U.�Ʌ �&ӭ��hK���IU�����-�}�>3�<1U�5+?����X����?�2����!�;�Z�� �3�ا'�����XI�8��
<���H�x��/���C�!���z�t�⃽pJ���G������J�;;��O�u��%6��PI��ٷT��H�}���#��p����RCpu�s�,I�� ���A����{=��?���d�Q�|u�9B����ĺ��q�}k���K����	���GR6��;V�tӴ��w�'QD7��4��"��9��\���GE�u���B�U�d)ot$�&��J�:�&%[�2��=�xN2a�tL^Y��L�����R�),�A��[]f�*�5�+�8
�t�D���a$nɎ�Pu��%�Ϫx�RJ��j��#�(�դ!!���7N����M(C7j&$a���r4�	t�n)q����ӊr��p�(!=���>xXF�&�����"�o�Kӗ��ד�~��WL_���̑�F�F�̞k���^��f&��=��19�I�A]�����T��4ܗ��)�F��Hx$(�ȗ#p���8�L�� ��ֳ�Z	�D�L�i�3�M��p�~�4�'*X9aKN��� �y�"'�аcuo�R�e� i+��	A���\�T�)j�*'��aϨQ������/ѿ5�GA�k�O�E�6�ܱ����ɒ#i~�h>HCKV�JS�O�[��|s:�bÝ�����W,{�a�����t��4��r��H@Lz���G-?�a��"��%�C���ωF�)��=��renך4-����h�--C&\ƕ�~���=��>�ُ���ߍ����b&۔� �FW|��TY�ל>�����uI�8I9�E[��/��3��T��� �e��P�D������؉��Z����a��κ��a���r�ӁsW�E�����K�X��ǅ>�(M�fOc������R�
�o��{�[��!q�Z��S�V?`;\b����K��Md�e���2�;SX�*��B�E�"s���g��Y��{��=|)=���������B���D��P��{� S����x�h�r�xh|�dET(*J-��g�j��ҝ���Ӛ�$[A0�$�TP��v������_yB���-�:�X�\3�Pz��ʗ���e	(O��U���*�^�q�U��-�"��C��T�L��_��'�e��u�t��s<��`W���`aR+�����,���.�4��
�f0��<����2t��IUU���y5l��v�QF\˓�k�4�ۧ�ɐ,���Nf��)c��¹v[��\�3|�� ��9z���3�`�y�;��v�:-���Gb�0O�
�/h�ѣ	����^g�GE`�l|�A���1��4\"i�C!Q��{ѧ�
�$���4,��W��/i:�FdK�4��O�g�ݠ���[B��bqsh+>����:�1w���!�Bc�k-�H��$��0�)��v�N��Q� ���^:�*��]$ѴqO%+��l}-h�z�e�F�B9�����o��������e%�~������ex����^j��vj?RI΀cY�d�a�f�U���2p�� ��:��rC!�s�+�N�6o��������P������$��\eRd��e�p���q��S�@/k��d�f�K���P�нM%��/��`�L}3�(Ὑ�^��b��Ok���A�S.����16Q if�k�!��	2�o��4��X�����jQrl^~Q��<��A��XR����S@S��j��ɴ�RH�������#ߣp��\��qr'�� ����:�"zc��Dv���vض;�ݢ�s�e��(Q�S��P�{���Y�~fJX�`�O���Q����ۖ,�g�ݩϑ)�d(�k���q�������l�QO=��1J���U��Ts9KH�\>:.0e�T�}�����߷/vy�U����B�I����Ժ9n�	p(�� h��M�?i�?��<�>:9]H���w]��}��V�e'I�J֘�T�3_����C��="���|����k�`Q��R��,�YL�*����N�����Oh�;��93� ��
�0uF���&�3�������z�|-p�Ъ*x%�-�AP�ԉ�4n:�� ��\��Z=�˵�y�Y���T�2������� ����JJ0;���9�4"�jɝ��s�Yy����FB0Nϳ�7�V+�Z��	��R��8[�J���\�C.N�W�o����:��`jz2��T?���
_k�tK'���Ȁ���F�γ�P��'��ej��K�mϏT_�j),��G����+䮩���W1o�˓�w�j���ul����>�]�7�gNu����;�0�%;Q��,]aӈ~t��o��5=X�r����5{FH�Z�p(=��j�����ɗb[2��d��ˁ��p�R
�ά�f��ҥO��{$�m9�Y
I��	�7T�6�'b��[��T�5F��c��{D�I���vG�&9�O{p_��~й�<�Th_�4�qy��3�ȸ[�m����}�:9�w�n���{�?��}��3T*�Y'��Hٚ��|�iy�����o��w���CJm�Yֺ��~��9v��kf���Q��y�Y�TT�,>���6S�Ҥ<�0�y���7xF����{,�i�'�.5Ի^U6�&X���p�O͹�pfv�E��n��rpaH�߉�֔���{T&o��)G�q^�#�[�2!r o��)@��쌉J�']5N�����E:6�'7�{��R�yjY�?�ڍ��m����`"���4j�8<����lafr�ɰ.��;��|�[��KTEXI%�?B�K8f�A2��C���[1�+�\yM��ߪIh���/I6�3.H/��o��E�Ϗ>�w��ȑ�,��Zs��qw#y�)�2J�y��F�A�:ZM�J��/��TA>7?�_���yxN�C_�i�U�U��щ��0�ؘWi��W����O�0�h��P��-����q��$�jk?���XDvp�����Ǫ?����~��Xm^R��^?��N"޸�yj��f;hv^Sp���e��]�˾E_�H��{���C�`�0hv��Q/�@V3��tc�z�<=O]T�&O{�%� 96Q���f�O ^N'��9��ܜ(� l3���+��J�5X��Y�{z��?�G��bZ�z��[\E�;uZ���<��6��ďX�N�kA���i�|��8Bpb�ɞpUE���n*UP	��7���\�js��&C�T7-l:��W��)���6H���H�4������K�0Lx�������(�X��>���"m�j�
O�-�;���3��f�����w����i|�,S�諻I��AV�^���<f�.�����gd�����P�c�F�j�Cj����툓&g���5��}��@TU������t��k<�T�=o8bEW;Gy���py ��y/D;���a�Yn�[��ĸ`�������Tv�~3xkb{G�Zr��W��}Щj:�k��#�{8��x�b�b������P���ts�l���S�ъ����!�#�̳��R�cl���N��y�5�ذ=��qI�o)���C������c1Ů<���9���n�����å)=oK�'t��#���C�x[�~ CK6��E#8k=�*o���]��.t�&-@�/���L�8&xyT>�m�a�5�b5���>9!`5�r�� $�7�|M+ Mq��p��?���{�F���k�͇*쇻2������C�Rl;��D�M$��a�C�sX>)��d�Ud&5�/��n/�r�ͺ�ѭz��%���UD�+�eU�8��,ACD��B��:�J��'6w)�F.V����+(�2:ZGCt��'��ouߑ;�" ٌ��LH�7 �$���[Э��p�7\�,��s�� ��*ߒ~v�+�� �-���{�Sܥ�973���1m��R��u��,��}S���8��>j�K��8k�4$}�����)j��<���9��*�a�: _���-Z�}����tV�ɛK/�q�E�쐮�l�RU�C�ٯG#xq���*�����B�r.­'7K}������e�{p˸�W�8S�v�[L���;�:��	B(P��X1OBm���V�#��
p���#�ɇ3�����&V�ao�3��9R���tB���+�{�5x��ѥ��E.4�ZZ�d��X!����*Hc�S~��-P�ǫ;��U��jLd �^�iD4���K��	�6�e����W���������2�(�9�b
��+�Z��tб��0���^WN>8#�y������*�P΁ݘ�=ҡuW�C�:��fU����
k�_�@����>�
�AI�2W�	+K2tZ4�\rý"}� ALv���t�⊇��)�Ve>��Xq��tr��2ˉ�j!�}G�x�{��'m+���7h �w*s�6ji���� !�w�LPO%OĊi=o�8�'������q�/�5:�c�-�Id1|����q�1���T���z_���^y'I�ޮ���|G�lsؔn���S籢�2U�E[�M�ZV-f�~C��7P�&�u�[�lh��`�^2=�i�~"�;�=B>�w�V���M;y,��edp��P�Pz��6����~i�tVB�2¾���gA��3�a�@M�ߛZt��Erqh��%�*��1�ΨM��IF��%�M|]�@�P�׏}���������0`^���iJ[b}`?��7e��7��������T�;�DC�v>D���fT�qdJ�\��sf�m{��4�&"'��Ҽ_&�RE�]�ad���﹕C���E��b�l�?�7`��"�)7�+b�1$�	 ~M�蜝Vf�.�4��*n�Q��:S��q����@�+8C�yP�0��� ?�l���
�>l�#p�D�Q8V�����U�LU�m��*�|P�o�r��W��{��� g�� �j��r ���j
��
��&���,���?lJ��$M!�\���m�;��dG�0�s��ɱB�="�����x3����Q��d��̅Fҳ����LP��9-��T�~ex�u�⩴�.�L��r��f��>���t4Q�qM�+I�� �O�7�>7x�ρ2�0�z�Z|�Z��X����?|<Ȉ��k� T椦��/>����ZvkD���U���q������x��N����������5fю��٩Haұ$q�]˂ٌ38���Ǡd���\wK�ƿ����R����_�WTS��jؑlk�G���'�J�G���`?�O���0A�����#���q𖞄� )���\H���J�R�R�VPw�.����Jވ���t՜)����}Ԏӏo�?��{-,�l�yb�w�j�!��I� ��2Sv�ϱN$��a�I>�j`��XI �{L��r��Da��t2�)w˳$l����ͬ��]����-�I��ñ���0N����]y:㻢q�?g�ӀL~����o�@�Ƿ�\)���k��#N�ƪ*!���ָ_�J˂�Z���/߮�	�o�3��
���m����k�X/�SE�G�V�(�6N����s�>������@p0C[��# ���Ea�a��so��ϰ/����H؎B��$�I5�S�W��ke�s-�V��{��bS��qo49�|����8��VG���dr��C �d?%�Bn�?_W���BzB�mkn1\?��|�7O��3�%Z��U��7��Ck%:�Œr%l� ,ѷ��M�Ӯ� ���������_����������QM�/��rDaG�]����mH� ���!|۲h&�oOpޯ��v�d��x3����W�vp`��I7��%A�Ħ���k�x]���0�Ett�m��˖a�(�қ¼���"��P����ۀF��Mt�+ (RC��%���t�� �|�uN�/��w�û)���^�%�{��ؙ�����ygg�r�-9�.*w�=C�Pz� ���d��d�NRN����Vo����〹�$�;���x�
����k2�����ӛQt�Ȼ/�¯���p1ə�ܣ*^������qP1M� e&������!��W4rC�4Dt��?�� i� �'K�)����Q�0yd��N)WQ�ӆH�L�#RL�d�'E'R
��v����_���[������%� ،T=J�|�ߑ��᭸nQ��v�"�Dm���6�QU��m��?���?�8?<^�ȶo�&����x�IJ��R'�;�cJ$��r�DE|"�;h�T�&�~�'���CVs'�x�W�N�`�-�'8E;������f���>8�EH�Ί�����W6�{+�����]f�z��{.���Pf^3���BG܍A�3`:� �i[L���B`8b��9 4�q!��b��:�k�+WP�,��c'f0��3��s�(�6�\���u`^�>@�zG]��d��?C~M�Q^0��СtQ0�bGQ.��TzWl:�yv��f������݁e��z���*���k�Dlh��s��D8k��l4�Hg����cTrQVhP Lk��~��i���=�U�N����0�	�"��^��}�>T�<z�M�Iu��+�;������:�P�&x;��/�K�L?A�QϺ1#m�ҙ���c�OD�sd�Dy�,�	�Y�~�fȴ�E;63s��\%0��f��`����L��6�y?5x.R���}��sȈq�.� ���k�����wN�ǲ	��/��-Ѩȟ݋<�<,��^�"/#)���ts�����ss�6~OJ� p�b�A�hP<�׿s�"�x����kɹ+X�������c����خ.��x�}�PXċ:�H�Ef�NB���&�����4o�*k#��/l$��v��'�=���	Y�qxb=�Ii澖��#f(���q�"w�!|��Jk���xPQ��m��4��=☃#�up/E��b����P'�����h�r]���R�Ѻ~�(nꝷ`ͧat��4����>�y�~#u��ky�����_
S>�<�~�ev^�lV�W������?�G��;t���4�R3sgN��够'
X���q0��|�?WUL`l��(Q���x�f�':��!,Ζt��f��|�X��4��'���a�DX�(Z�ekN�*�-�C6�z� �<�RnJu0ãk��W9�����Z�b�)1����-K�ףhOS��e�5��uC���fY8{�@�I��_�q���1e�O�5ͨ�/�Yk�2Oʅ�8:��2��Ս��=^JQM`�QY���Z����_��f���B)V4q�V5�"�O�g�G�mY� �/z�7��Λ���e�[M���w���(�0�[~s�IZ�T�H�)�=[8�Iw�4�征H���vҋ1����-r��
i�q�<�֌N�õ@����ӎ�6�|Ms�1a��x��ы���� �'(�9�%)Ahf8�Y�/q�<���l��
$�8v,�c��c��b�Pq�ӆ8�c�:��r8}������̗��$�E��M���2��BEi��'�c�O�(�V��&���������Q�.7��dWW�'�:������X.\��OCSM�2S���g�ZW�[*�b�E�E��J����'E��/y
"C^�ŝB�)�&����I�A|s[��H<�b!���o/�AI\#���?Z��R���C�_�#���؝��:�B�����+Q0��-���">wN�
B0<�2:��,�J�l8�,�d�&�jip2�~��]��u!��((�>\r��}mA��2Hr�]��3ȫ_��חt�1����`��� ��)�[�r�b����m��s���ʨZI��Ÿ��.��� �:V�Ju�XX�_=��h.1E�S���CN�M�i�ew�%KĈ��[a������<up�#z5Ӊ@N^�f�}�EH'��	�ѧ�iME�`փΪ��5*�k��l���-;h��Y?7�O����kҙ��%m��}�.����=�2�ݤkJ=���S9�<SJ�>��)y ;�Z� ]�cZ��Q��Z��`W���
%hl]3�/ס�OM���`m��q��'�5��:��w"q�}U��&���%��"�8!��Q�(����KL8X���?�[��A��,	{����Lˏ�`��A@��(�P����A�.�5ۋ�]�6�;[����_��c��� 0 nd�D[}pr�G��<���-����@2�&c�
���S>`�7[~U �|����l�l�9���Z�F�F�����NL�w,-dL�u�T�� �N�\����:�/Wa��&���%�z���K)A��д�t���G��XH��[P����3�G���y1Z	!<�/��n�ns��^��l�Q�s��Ŵ���e�&as��Z�UX�J���;]ϛ����OW���e<<�j�Ҫy��&Fp:)�p<��"�����\*�2���gۙǀ��,aGa����n�b&��7):
�7�Z�JE9���W!��
�k�t��-��������R&��dsW�Á�_.��Ù�fM$�|<���P�]���=��r-�#ؑ;K���"8}龨�(�%-��V�%��R��|�i<�����.�g��6�P���C������J�Py�~� [G��'��c��P/�6BZtS�7K.	|j5�/��R�>)䦧e��ēs��bACP?7�ɑ���y�S�u�I��QBG��.���!�'�8�l8�ވ,e���`y@m����L����yL���1��o�I�:7��;ɥLm�t���t`ѐ)���ƨ�Ԗ��B���"e]T$�q�5T�Z�6:��	�4����iP#:�I���H4L�rH������n)a�q��ޘ��"H&���>K�Gz���/_ԛ4�]3�M���k�q�f��O�e�e�A"�����R*�}�{16ʋˬu+�ˢ�?[��fc�e�),S$
�[�G]%�E6��1Z��ktW����,�]���`���
y7e!�7QuD��� ���.�g�i�k�˼���s�x�����W�ȕ�>��Tw��j��8���*�ɋ�(��SrdE궼ل���A��vs*7��]v�'�j�y����b�D���.`��8��
��^�)n�e�I�Dq6�g\8��ZAS�0V$���H��0�q�^!�����J5�Å�p\�0�FG�}1�~"�O�d�o�A���r������X_�Н�˦^wƅ4����x�a�Y�x5��\�=�C��S�QO��H�H��V2;P	R���C�营d��*%�=mJ�׽��cB2��6��A�i���'Dڀ)�����)Ƌ�i���#tD�8��&5k��cl�6���i�ܺ���|��{ ��.�r�.
���`C�	N�g�@m,�B��:�&�G���s�����JPYBq1��U?:���g����0�0uB�a@�I�L���;�R���⌠��_	�+E��U�SR�%?I3�'Ǡj\�q��fj@�ͻJd�Y��x�~������zpGd�,�׳n*���:�j��Ĳ?���\5��L��֟�k�P��b��Ou5�PHv��ݚ���I�*FA�D��w���K�^{4~HC�8�6�r��a�CFH3�V2���}�Q\FF���X�*	��@7���,!/�)mC�k2o櫖7b�����s�SI�H�w6:g����b��7�lC�	�ƇD�7�F.j-�Y��낈6d��#ت�Bc6�����p�E��x�b��\�������7�Lad׆b�3�7���m�SԧK�F+b ���ޛ���R͞@]v�I�3F�};�[Ԯ�n�s��zg/aa4�}_�.�������2�EEao3>��g�M��٠�NM̀��vv�N�����ҳc�NV�Z����j[n)�<Zb�Znٹ���hJ����I�=�9�&��y���h0��˥��u���Y�D���#
��`lD�#M�X�m>=ѽ�s5"@��69��'}�3�R�s�⡳�j�ڰ=��{U
�a���%.�	_EC���T��W��	�l�����y�N�@�umz��K��ej���n섎�	#�r����Җ�O�C�n1��#�Qu3�K��H�&�:(�'��A�ȕ�(�Fq�� ��N\�6i��a�l�O�G1W�>KR:���h�V�kF�&!��v�U�3#
i�D���2`�����FJ���R2и�0]�ER�՛��׫����~'`����}���|_4ܗ���*�/�[!���Hb-�A�G@<�HB5�$Sv:�B4���2�c���P<�B!����Z�\|r��=_N��\�Q��ro�����@��>�o�ڝ�����M3����״D*�m<"�u1��d
�����4ֆ�2r��Uo����-��N�G�^J����F�K����?2�wn?US���Ҝ���sV��w��4�$R*�A��)S!���"%I��'�:,j?��7�m9�E\�甦����������๺�Sc�e������^��S<�l����5�Al�ŵs]�Z�s�*>;��&�*��;�v3�N�մ%�'�����>�"��-�g�?�_ϴ����Q�!Fx7͔6��ف#�9��aN���L_K`)G���r�W-%�� a�s)�%��������w�� �A�h�,0����A`��T�:�-CT�����
��"L��[�I��g�Z�:�]�w<��^/��kiF�+��+'�xUZ��c��N]��&ǈ(��z��7k�|a��Caٴ�`7v\,�T��$\@��������}��Ї{YP&�!y�z��4:l�{c'y�!P?k��g���6��YQ*wMS���dB��?_FI�hq E�}-n�i:�1!�lgGEr2���^�u?`;I��=g��M�K�d���F��.�������h��AoM���?ڳ�]���?*;��xϑkZh[Z�\���3��4��I����!:��Y��:�5��,v�pUs�X=2�4��I@jHЅ!�(��.#��`�Qϯ�J�3����|���L;�G̫���Ͱ�]q���e#��(:  $����y���������x5�PV�g���!�r�:�{�xN�(~�\Qnƥ�_��w�1�X�+��{��K�ᎍP��+�	�W��lZ��]B,�K���X�:������/���T�hk�F��1Z��� ���|��C��Ryya4�c�V�}SaP��s���]��������d�LJ�Lp�/�O�J3�w*'R~��4G�>�!a�D�`�G�`�f�;���V��;EóM����~�/4��+W����4�@���D�X�Q���Ӹ�h#�DW��3���
q�>j�R�p�E��4Q�a�R�C��|�)���D��$v�FczoL��q7!�®5U����w�5�O���Ca��A�"�-�*k�w�Vң�f�T����iQ���>����گ��!�%)e�Ӽ(�_��C�>1�mtK'�%y{c�������+�$!&Måw����}����d�� 	������R[��DG��wMA�}�鄯���O@F~G��0~k�"ܚ6`qPU�яW��kUk�;!�sqe(�T�R8��|�u:5�w"2K�d�{&[�O��������y��]˴0'�G2��e5\�>��uyG�gɺ� R��ck�`�'?XP~��)w�̓
��j��Am��Y�+�
�����ZPA����_eKm"�];���D2�.R,S���^�V⅍���]/�<muR�|���@��`���qf�k��]�4	'qŸ�xZ��;g���$1��fm��9�D4<���S��4Y�.Ê�nR�(¢%K�����cڨ��a�N���0a}�j��N#�u	��\�*�;~�cs4j�Q9���h��n��qs2MV�k ����3D0��	���Ї#l?:����-�RA"��M��_w��S���wrR}/�ּ��D�y�)���L��ڰZ��9o�3O-�{�N�kT;�����3M�)�NC&�N���z�@�%�f.f�1@�|�m>��S3�@t������G����݂�W�$�����{T����p�iBٽ�߮s��w{��׶3n�9�E��Q���[!��g��e?����o��j�*c�7��W�_��1���׊ԙ3v:ӧ�5��R�X�KC虂��I���sD`䘳"6U��\���zh�Kkj���I�i<t��Ɛ��ЧVᰊ,I8-qw,^�ǀ`o�<�$#�rq�)ol'����\�S��~�,$b�Z���5�/9���Y���t�/|[-�	0��G�{�q(�3���x�ӧ*��/&��K�N��2C>�/k�# a��CLL*.��F g����v��L�x��AK4��Z���@��f,�?�Xf{&٢p�0�� �0Ů�_�\�Tݙ�C`�x=H�`԰W ��]�T�k��O톑]�7���2�=U��L�{3���>�s�+4}:1穮�G��o��Sh#I��?1��S;�: �ќ�R�G&�}������Yj��9���z������o����5s����6yU��������2�%���h]:�!^�-��SF����
�lYս%f6���)�b�f��0<��4kH|W��a��y�U������(��gO"$�t%*3�au�&���ޓ]!M8��gb���4TB�j�)q$��ɍe��4����g-�-r�߫=�w�0�!Y�;i��F֥ꗌ�����{�����.��~b:ۆ�X���C�ǍT�q�wu��A�Ʊ[������u.�#UhK�3��Y�*Bc�F�*s�ƩSD?B8�`�L��7L`6x$�(���J�w�;��!@�#��U�Al�i�b՘�wv,���5�/+J)�7U����k�c:����D�[�Y�O�
�b֒<�g��5fr֒6It�w �0�������Nd�Bk�2��`�3�'�7�/��GDِV#�=M=@=tG������t6r���A�1�غq}�.GU�X�[
�ԍ��|ّ��U��NW�:��O�y�W���JE�c�]��}�<w������x����gx<�buQx]��۽��n�jύu��L�������4��?��$ʜ�b��o[�}��zL��P��Ԯ�4�8��|�걔�)����ΈK�����9�g
�E`M��8�!�K��H�.�'2(��{�3$skb6����d�Ӊ�>bx:�� KA98q(
PQ6����D�_Z���xJ*�2��3I��-�e�z�~]�L	�y�����s��ȨT�\�o1<Z"�>�x��������:�Db��d�������k9pLAbi�ABg��]泿y��k0�UW[��qZQ��3���zj�'N�ÝL��9N$����f@h�s���s�5¼�Z�l��c��2I�t}]�/�+~�j�*��i9���m��2��N�DvRϣ�������oq�tELK�@I�ӡ�	.�F���+n~���6梦��툭�Z�%��`����8�}ii͙.��q	�j��x$]�M��qԙ�R]3tط*�Fj�^ud��F
[��cи�vB	�����)��OE;�a�z�=L�\��
�T�j��v���ݷ~��B�*V�p�(έ�c.T��c��,��ׄT��^�-͍���I���f�~|�j�11���+E���.>1�t���S/�f@�9f�?江9��1,Z��W�V�ӭA�W��lo4+$�S����)��ʙ̘��`�Fc���� ˷oyi������n-�z$���cM��s�Q�T�?�惓M�X^����S�7���N��0�b�,�	�����*������=s�n��C��	ox?k�K8��+$!�Yd�V_���c�=����k�aO��_tJ���Ľ2N=��:�y_P��q��a%z�3�#>�$觴���6I��b���9Bh�|S�ͫja+Y��p������Y�dRK����;P��G��4���4�=�y��E!�y��9;^�L��kdݛ���Si[��$���Hh�Xz=������%T��K��T�"���qT�@�u�oZ��_�'5�D�Y�:	}��r���,�HM��h��(	�3k�^njs-�ӬA���.V�9!8C�`�8�*t��@Vp?��|:���2��@���2uŪ�����/�U���|H����֐h�Ǻ\��͋�������,.���z���4r��4���oX�6eG�8B �.}�RQd����hxA �-9���3ܙ�x|]���Q����9��1�
��z�$a�a�9�.�D����|��\ǍlҊy����]���G)���[nK�;"d��L	�h`;%�G.�䓘���nH�������o-��&��}>#�շ���.����Kq�k4]�����fR	)���^Pf����UT� Y a���뜐[�!�= s|O�}߶K����iF�9�$�o�S��s��Q����.�fڋ�:�QP��:v+-sN���(v��s
+�o
`	�
�d�e��7
~ Ǧ���E���Y��	����<=~>�r�;r��)%�Os��(삁��TM�|�/��/?�3���yʓl��X�I����l�$#Y�h��������PU��r�<�3�.���A�(�ѦŌB)$�GX�A��iy�kx�F�y���A�W:�~u�'l)�ì���Hf��1Z�*W���?t{.�#�l�BR��V��� D��aU0������.e��]�f�|lǁ�mr�:���Û��	lH��Ó�0~X�8����FOu�5;�T�/z���$/w��!P�|���?���h�nM>���:�w���k�w�7�� ��.�|⭑Q4�tL��K���`�� 2���[-F�bc��a:;&nV�ԌX���@Y��!�&��7bD�U/� �A,�&"����7oV�1���y}8vzG���}����H�s�Nc��Ű��\[p}Ec_�<�6����J�NG��H�8^��ⴻ	I�9]x�C��m�e�r9,V�؜Zކ��d%Ӌ�))��D�$�����5�pl��"2�Sc���\��'��*�Ӽ� ���BO�$eiQ�+��-��׫ݢ�@���p|���D:���ڈ�2f�@i�ݑ��Gq��p��)��1%(�Q��nhy|��W�gLI�*#c��251�t�Y���i�%y�]���Kg�AB�qN`}��<�ix.��~�8���Ayoǡ��e����2���'������%��F��rc�T����H�I��j���Ɨǩ����Jۮ3�jn�|Vy������o�Xok��{�k�5�&Ԗ�D6W�x�b�5Ź��m�ZzD����%���8ѿ��FLC��8��8� =q3��D��'�+@�Q#�"E�H��M�S"�\Mb�v.�~��Qi P#P�=�K������Wq;bEq_5��_�v��|C��t�ϼXv���݇ɩ��~*S�ccE�K��$���d&��5htߗ!�G�Jv��D�e)g��}yLمeO������)�Q��ʕ9��QRr��C~b���VG߃$Xg��ϫH�c�v�Ɵ�~u�Z�y��z�p�~mmgE�~Gz�/rk���,��,�e�b��@�MȢgh��=�y�=a2�i�	�M
:0���nm�n.���_����ˣ �S��P4Q��Lۇ��M�W싔�ϼ}(�Sx���b7���0�O� �?�_�<^� ���\����N�S�s~��Tpw}����ՒZ��spr�\�F���4Ե��v��X\u�*��"���c��=�XGT�J�܈���J�P��=�2��Ub=O���|�C���A6a?uX�ռa ��f8"���NS�d�q(W��r�Q�n����q�<�AVw<���2;�/�+4��..묷5�Ԭ�8k����p)j�o>��6~������ɴ��3O�Ԁ#������ <�&a����s��q�a�#@��-[��ķ�:&����7�2S�N��_z�q�D��B�s�u�����]���1-�|$m��};M�t�h3_�cRj:���$�@�U���(Fa��m!]~��7�Q�Lt��^,�X�O����)�!�6����W\�-�R3E�D����7o��&1�]8+U\��!}Z\�G�7ݺM ����8s�I�T1�4fj�"l\~��.��4�%�

��M~ ��b%�>o��W�S9�Gڜ�Z�����F�4���S�|�Fjp�Z�5�-�oʧ��j^�'1����f�X&�o���C*M˹��p��T��2�{�G�*]4�8���oeC�?��8��y?�LѲ=��t���J*��^�
e&5y���m�pH V��I'΋WM��罉�.ۭ�64kUQv��_�>�[��z755���T ���MM$o�A�sXg��>��4J���K�uɚyc��� ��W��8��8�̈́w�i��<v��O`G�S�ߩ"@}|\�I���biO��8H��)��n?�����'�ӏ�hqr�^�I6j�k駙/N��0�D�FP�p|������Ns<�_^RIQ1"������2;y�M�>W�kZ�R��#ک}0�q{�[t/��4!�犏}Hs!t�Lξ�守�NJae�����Yj^G2����L �Z�۱W�8O M`���]��ǌ����+-BO�M���)Z�Ҳ� k�TA���h:���7���;Y��P�v*iw������i�ƴ����or�y���t�}���®��7˕�˖�'6ծ�~YYsC�j�D;�m��;[L����?�.s��)XLn�C�b'Z<��⋏+�u�eహ�:��
��|(�N�V��1{�"͑"�F����H;���Ă�oܳ�v�@�2s/%~��B)0��HS�(��D��c�mQ����h�D�GW�w�1~���hy�ck��$T�� f�i��Y�e�6f��d{��6�+=�le.��14��s��`ڒ���zW��_���a�W�ˮӭ7�gP���uu�s�m��;���sl ;��8��T���P @*Vl��uoE�u�������������7y�޴�9������DUZ�DaP���F�kT��:�3\�����iSQ'5J����� rV�֗=���D2hU��i�E��!T*�O�LӴ C�7D�I��؞Iչ�l�$c�qc��!P�?(����y]}0�}"��Xܡ����ҍH�k�ŦBx 1��U���XP�l7$9�Q��0�\m���w�v/l7��NXr��7�6�� �Ffi ̰��BpCW7/���Q@0޷�"xy�9T����G���j�>��-�E�w�8��*Ǣ����)��!@��b�lKX@�*��dc��(KӀ|n�,�|�KiZ�8�gm�Y��؇���b&�	���5�\!�ĳ��}8(_Cd�8��-���3o[ҹ
�O3�38�5��V���5��5-y�&x]�_4�1+�p�QOn�����/�W ��i���w�������C��X:���Q��|�:�L��	D�R��Ge_ڝ� ��2,O����}�-�s=�&#���{�H�	�6�k��B�~J�b���I[�0`�+�,M*\2����{�M+��4��y`��X���~��#�Ӫ��U��K�nWD&����Q��Z1)���`�pj������Di~0���u��,��t%�-�zi�]sB�^\�'h��㞎O����P�ykj��hr"�-��}��p�4����(��N��nT:��������h�U0��k��/�ǆ]O�@�Ԧ���R�q��y��;��N$��Ԫ�*<��\7 ��o>$唢��ؽ+��g̝<���NYM4X!`s�}���i_��=�������m�ѺU��j��~q�����Os�*�:��Ϟ�4��S�P��!y@�_����6� �2/j����*p;d���	�����
���?���Mv+|�F��;|N¿�ך����7�c�4�Ue��|�ãwz����ς�sF�wО�EpD\������́51�Ro�>�o�[Ω{n��"J��������87
֋M���e*�k4I۰f���Z��.�|���X��,��jw}��3�2�e��Z@����3X�-@����縙[+��d����+��۵��$B�vOɢM�D>U>PA\7�*�r��vdb %"����6$�����@��lZ~��Ʌ����6��LQ�Gr<��A����d�D���5y�����V�����򦱟�E�l(|����F����##�P=i ����3����>��b�i��i�����ќd�j�P�X��Ng7k�y��Sh�խ}�c�J2ot���m�[H�����G-W(z�n{SkSy�S@.�!��a[c� <�2~;hƳ�a���؛�5�h�0	�"9y�i��f<u5��u�&?�m��<�|�7G�~���I ����\���i�F^�?�)���+�En`��z~����B��Uְ�� ��Q�0��-%g�o����e	FY�%��L�J�P��!ZЄ'�mH��8����ߑHz�QH�Ɔ��y��\�(�~L�1�_[��ש��D��!cϜp�v�uTaV�;�w�����dŨQX�Gb/�6���QľF�iۍ���,�����*�o]� �y�� �D����¿��=XGA&&&�x����q��Ӂ��J����B-Վɹ�N����j�~�D�|_��]�f�v��w^	�w��
�F����h���rϩ ɖ��:�{��VWZ�C'�X]Ȍ"���Rz��;�Ēsf�2�x�x�ZBk�r�#|�w �����|��#�ht&=VP�����7��L��ؤ�k	�ht0DO-��R"!�xJ�$Ey�HM��Cr�ep[�jq�Y���ѵ��kC"c��[-�n�7�'��*�rexs�e��u�;�L_m����:=#��e�,��]N�w�Z�t��^F(�����s�<�!F�Y�<��TT�"��})��{M��t��+�q	�JR�S��YT��HD ����HY?�� �L�C� ��� @&�����=�MA��E@���YO��V�(^v��J��5�����C�Lி�����`#|���}�M��{˴������]S�J���Gu�����W|q�n�[G�4w�M������P0-�+y��S������;��X�c��/ԇ��ʶѹ�?����v�`��K�-`�����=�l��C˒ Z��X�- �~K�\c�5��ڲ76nK
�_�":��=Gk8<}fc(�m�H��H�y�?�u�&�x���Fv�dq�[d1�9x��dNj�C�B�wK�8��T*��0���#	��c���ͮ�*^�Fb�2jPV]�����4�� �m�G&��9���V��tݕC]�6��y���	r��
���s `�+����W����V?&��⦻��H���d~r8�
e�r#�\Y�@~0)�w]��:��Z�Mfw���W{��s��#L��T
���bH��jt"�֫PZN�:�M�;�E{m_"r�["b=�B�1�I_F�?�������'�ݍ��Į�-���(�?��;��X"o��U���Q�%w%�@�D�V�Ԍ�m�L$�%N)7.�����F�c�2�8���`�.HL��ba���Wt;����H�3��\���J���
����Q!Z+U�A8f�%�h	<_�
�� ܢ4|�%3�V�s`
�k��K�������)Tş�-�?o5?����HE6ae�}`аX��U�3�&�'���H�^5�4�E7 @�}��ܵ/<k�_vPG�/��p���������~�>}���a��]F���	,�����}/�.���xL�0���%�]�B[9�����χ�d�°k��R�`9��,�S��7,&���,�:�ԝ�A�0��!�x�g�Ni*X��Zܪ�Dz��iC?�>}��*�+3����Hcg�/:��F�|:AX����k���?�nM���Jv�>J�
����R�&6�^�s9&,X�k҆*o�m_�J����W�:��ߘ�����u����1�+G��`-D���lA���$���x� �K,���t��2�'؁�Vd�D-��Q�I$��8�+��L���:��)VY_���ՠ����HJ#�ya�يR]���#%D�Xh7�5a�<ݧ���=�E�Ū�!��o �Ri1�a�v�t������ݩ�`LN70�xé	���~�f�/
RY��������nSm����J�W�u#���n#�59dN�
8u��J���:����0�K�c�X�w�����m���. �ppVȓaT�s��mިvd���hd����`��<ܼ�C�QD|���4����������� �^�Eh���cف����#��Io|�餉�X^&w�Kn������G������]��m���R�$���_b�]���4���\k\��>�	���n~[Jy�\q ^�T��֫�"���XR�\o5�1^4Z00�~_����R_)�m�6�q6la�`��jݎQw��Rti2�P����.��رZ+�)qe���W��W�Uŧ���1�x5�uJ�T�5����s�\��0��������VPtͅ�%IV
�\y�P�*_^$w�6'ԅ� u4aU S����NUʇp��L��C)@�H�`X��!@Q�~���5��s�l&H��n �S���.!f,}��l*46���;49��d����bѹ�h�'�x)�'"�1��"�E����5�w-<���`,W�����RZ(
�Gs,���ݍ�y'������#�7�PRr��/z[F�>�+��s����H��"Y��!�K������QN�Qd�(���-�F�~�r�5U"�xl1d0��G���������uW��uxG1�4}��n�3���x�]]6�c�]�P�9o�I=�voMT��!�Q��SL�<͐`�v�����U���3�~�^}����� �u�\�����'��/<nfH��`/T��4z�f��/����i-C�犽���4�|�o)kO��d������T�E������p�t��s��G��C��ZcK�i�ӓ����N��K$p/-قc^*�;�H/8QƢ(_N��)�ͻH�"�_;�pӼYԮ�4�0�O	��t�p�7n,q��v�9q��ڽx�(X_��+�u��v��+s#95�W�$}�Ͽ5�<���D�Hj�����g�q�_�{�}.�4��k��.v��'�j2� ���Q�Ť��7{~g����6)wT�'�C������hؚ{�ǜSP��%��c�ʸj���}��,S:�5�tZ�����,C%-(-�ř�b|;��H"9��C��x���0��]Bq�^����E�Js���op�������mjF�qp�t|	%k?8�x�����v�4U��ܔ=3��-,D��#	7Z�t�u���;�5I��l�[ I����.��0�je�M��l��R��#p��~�)�x+��.ޑs��d4�j���&�f^�E�L�ll��5	��KT�rwS[��S:=	&5�Eh ӵ!n�A޸�P��us���7��y���C#��m���<B��5k��X�m���m��/Kݝ�*�	�;XE�'
��}Gy���Y��z��$vgG���~$30xfD��;8�t�0�����g¦�ܵ��"Z�"ϠFh]��h}2C�W.� ?�-N�P"�܇�>u-����L@�b[$ȳ� ��2���.`a�2.N����o�h���� �q��F�2�l��K��]6v���%��7fH�I�Tew�.��.�2"�mS⣃�R��?�B�0u��P��}��9���`U_ !"X��۔�8�#\|gN��Z�0P	=�1U8Rdq��0���&E�}^5�!�oqy�2~C���bu�t�A}9��I4/ �V�)Z����jѹ��9�T��#�7���P�g�}�����Y���Q�R�U�LK�Mf�pH^�*?[._@�� xsJc ^!���tj��_��SNQ��7F@�-n�����K��h��)ʳD.�Ry�G��/��	,�a/�.�9�`w癨�7Թ���.�&�#7sm���?�|�usd�>)1�H�CH9��+�# PGw�x��FPo�w���T����?��c��&05�~��hH��`%�Z������3�iZH��O�ggg$�Y��]��&o�Y?9�6|4˲�2n�h�nI���!19�4�8��ձ�?�.�4��YOE�Ǔ���$}+6�m>�.��3#Qp��\��,��= 1��ѯ��9,,-���d�C[��e�%;�D�	R�����1���x��+P&�.���cE[�Zg��s Iϋ��1k�OL�����Z}X���V�K�Q����85����*w)��Q]��p��]�&��g,�&�Jv�G CU=E),���;��H"o��@�-�%�;�"�E�N�e�f����A���XL&��V�Ylѥ���d���ZZJ���J�"Va0�9�Ns��d<K6brm~�����F/��'�ی?<x�E�쑘�%sh�Q�z��s�򊺣�T�Ft��-:�����-n�e��ٱ�T�	�xvs]����,3���� :�C_�T����]��Z�H�J�Q��E�P ކ(�h9�RϹ:��4YQ+�?�	0�y��g.$bĊ�+�>��p�K�M����ID�����g����ҷ�C*kD?�H�vR�v�u�Z:!4�i��3��j=2L�U���ɧ
�g���ޕ�P�0-`o��P}E@��Y�k�X�rص�{�h���Ӈ�V4d���F�:6l�ɠ�N:�$U�N5ocA����~�)A��-5�fbT����G4��" Esg)ko��p�I����v^��n�-��@�%�,�SL�d�w��Xm��W�DƂ7'rg�X�ULc
�m���e@'2��|��l�ҀzOξN��>(�Ov:ƣ�'e)KV��r�(x�5�]�k�&�/�"�ϻ�	�/�U���+���!�ļw!��v�������<~y`D�#�+�˛	��l�E+�i�L�%��a|��3/$���[�f��஼${�,���r�¼S�J
0�cO$n]��A����u�#����M�Û7z��q\2J6��r��G~d��o{ksm!i���T��)G�e�魘O)�@�.�̦�t�nv�|���$���cR������)�J�_TE��(o�H��32�~�h �r��uׁa��Z͜z^:'�5�2\�4�"�?��o>g��j��������{� 3�G�6a;�s�UT������P�� �'M��E�~K{ڕWln���rs���V�oC�6� �x*�,G?�	�q?��C���/��c87	��o�Ck�x�=�/g}@^N�9���Zt�8ғ�}�\:�
D6�� ,e����U��$7kD\����,��E���2<v��!��"�ܵ^������0�8��e2�C��c�?+� �F�� + w�a�c�su�����.K��U��9G��9�8�\�4\�O周��uu�fՅ݁��ϴ*�k�]�%
��R�
�&�8��Bc��:.���<@%��qC`ۆNn�����[6d�2*����&pt(PI���!�����]<�߮9���TH��S�ظR�#t���T��5^7�gpZ��������LZ�D)����<����q#���2���+�ϑ�N�+�%�N��%��?�pȦ5�J�-�~ؑ�DA1��+�@�?��;dӥL�qe��F��o��y°3@�[��<l���̲I���J��m�in�E�eπ)Vp����ot�Q�F̎�`��%ʢL������UF.xnH?rk'^���C(�أ��(:F�[ ��b��1;��	�\�����I�����psX�5/���I�΋�>9�t|�9 j*1��S:�np}h�u�Iu{�����C�4�@Ƒ��.�#г=����Yp�s�UWo \w�
���R%>��Xߘ�t��O(��=R2?�Ċ��?�%b��oRx��w��-z�ZK�]��]@.��M���XB��G̩Ŗk�]2B���#@u���(��ŞFN��t�l��P0�,��C�J��Q<>��|��ci��u�rT�``_[5��O9����x�f�v�}�(� F����5Ǯ�W>P�i�; Ug&JWƒ6Od ���.��Z�Lc� ����9�U,q�t,���u�X5�v��c�Kly� ׎j��'['���ihUS��?i:�	��V�2}�ui�g[
؉��Yマ^1 �%�<��+eB�:#|H�Y'����"����h�/��w�>��"�4����E߆aC��%�?���[ْx��E�	l<� �4�A�����:�'�4jr]q�(	A�н��{���vO�6����1+�ƙ��ҹ�p�}���C��c*$��)�o�L�e΀螾"��������ek�V֋Z�(�,8�Jp�p�F��%���lŵS���+��x�~�.��UI���^y@L�[S3�H(�#pm����0�n����L]T�m�����n=e���K����*�J��Th��j%T]���k�� ��#;� ��/��|���l
�g��.c�<��I�T��IBA'�&	y|���[o�M����4�����ԓ�Yu��!ԫ:hl�t��'D���G�������4p��DG��T���ߴ����f�����u��P�Ø��CH��?�lHsc|���Y�bp�1�T��fqm�OY�t�x�,,��K/k�p�m;%Cu�r����0X�{4m��U"��:�0�i���ĥ�\S��c07��jpk��Ӝġ�Ne̻$�䩤(K��SX��[��oq�I�6�w�k�O�Z\�{(�����H���39�� �9�P����E�?��_�Q���B�&��ȷ��G�T���,/�aJ�@���C��Kx�s��}����_�t�� �R��{�Z��W����fg]A�"ɴ�Z'?�	&ېK�z��׀�7�B'��|b�X���8��a�;��"�$�����O ѻ.�C枈yA��Bg������j�I��������	��Uu��b�`�C���S:��o���r[�'��iy#�WǮ!\�
���a���/ůg
r�>(~�_����w�&@��kЭc��j��b'�yU1o�ɓ��%e��>�1*⿄؃~�E �8�5T��|
���T!<t�.�K^��~�����a��u�`��K\�s����n���A0�V������渨�e'�\�\v�F����NO��,��?��IK�q�n��v@s" 
*��]���nǅ�����c�
еl��3G��&�4O�3ű5�چ���v!]�����RFPr-3D�L�R��z���	�ŗ�>�Dl���ᚫ]�cHD��8�ey�,fg�Bͩ]aM�a�A�N���ȼ&m�Av�n�����"��U�^�X�����h�s����|��yc�u�W��{	�"�匩�=Ȋ(�듥�lKP��2�Z W��Bp����Uag7���-�D�_U������S���7�R����h����dNk�]'�r�6M����t͂�o6B�7pa�ޒ�ֱ���+9����q�ی���C�D���ا9��-ظy	�̥��o���d�_��ɚ�$�X�L�J- ���@����O�A_�h��	��w�?��B��n/���n���E�G����U�BP�?�[^�^�'r�ę	a�>в�	PE4?�����Ջ�?�?�PF����v-��:�s��!�'����R����˰�j�����u�7��r
�uH(��7~A��|������B,Q����|#r΀!���-{������#�@U�^e�I���j�������9ՐY�6�-�j���P�3��^��S8+�ت5Dc%�d0�!2���r�
s�cʤ���uC��p´�6-�^͡��/�����뵛���Vz�){=u����������$��Y�U�蚙ߥ ڜ`^pe��x��*9�e�?���8%5������s��=���FH�%>�k����c��i��H?1e �� ƺ&]��W�	|dvjC|$���]�����M��{�c��s��+���*QT$��<=����#������IP{�W�A��4�\��v�Ӥ��x�L�e�W�݅��CZ�`h��	����N`,�ő�>�ެD�k&�Gc��|����î���+G�#��<�u���a��.��Pw�r����p8e�>V�Rz�2(�8K��5[O���ݓm�t��%l��-5�����~X���6Z�%
[��op�G�/�o(.�,ؙ�[0�C}�	�R ����m��
#����͓�Cw��?�B�U7_�b���r;>f܎�e��WwI��hjk>ǎ�>O2�ks��ܟR��ݔ�Gk�^]ѱ��~a�F@Gpivy1e��&s�wٴ5Q۳盒Ktw��%�?Xh�Խ����+r�5LסlL�栵*qࢹo�([m#}v'��J���*�V��HQ�<nPX(����D�*y✲K$��p��I��w}��v�jK�^z�i���@3v���
|T��uxɧ)�ￅF[�$��=`���*@e=&"�&��u�E�D����p���ǩ���y"e�u=�<���'2x�!�pp�{f��X1$�(��&C��q�s��.�H"B���Z�O������X�g�'Ι6�iX�I~��`��<,}��6>Ci�� �o�=|TB^!-˗�wx�������~��q�]���"	*��x��*(!՟�̂��b�lޢp����MӰw��bc��N'�"��j�Kj�_[v�D��Ɲ�z" f��m-"�-�s&�n�K�Kp�ƒ���3�9/Q�S���ju0�^i&�����#�ڟIہ�u�x���1�o~�f�wG?��ysu�"�q���`ݴ?*Βm_�r ��ЃdBR�*����S*]�np�6qP�?�b�ۓi�1���EX�95|�E8��I�����^���q�c�) �/J�$(H���Ƀsu������IU�Iw���R�X��g0��Ǝ���J���]d�UmA���7�Z����~zcy���
S*�p�&{z�Z�!(1�jr�u�G����*��m FӠe���
շ&���^@�,>�۬_>1E��5��'OI�w�sI������2� �!�q2��~
v�6�O�1L�?����7�'r�IK%��Ea�ֵ*���G��[�D�X���G�#9;��ne�H�1SRҲ$I_�ľ�2v��~Tb�ف@_lz%�AJ�D�q�qR��|�뮨V�j�=����t��G'.Y��Do��׹Q��G:�4t�*�v�<w/۷GW�y?��9��le�A� >DI������Hej��Fg�a��G���'Zz[������$����_g�+�4�N�I���{Y7�<p�ie�{�;/@��A&_F�ļ◤C���y���Uc����8u����h�/a��U���K�6�G-��T|�Z�8Xj��C�F��x�~���;�
ot�Ę�PQ��c3fT	-�b1%ty����B���?�̺��+4K��j�*��<�FV�V�#ZCh�c�A���
v]�t���CY�s:b���6�pQ9c�\�S��hwt���5�� mpN&�8�X��j����"J��~إH��h֯s�����={�G��G6�ͲD@A�j
��m�ː<�8h@z}6Ҿӂ6]�����		�̓�X�x�Q"x�U�f�9ݹU�ˇT��ǹ���y�!1�z%��J�����*Z�iA���!4�E
�l��X��c�Fk�W�?��������H��U�|Ϊ�TL�U����Wg��JsƗ�-����7�c6��C���>�����6�^&�~֚�ſ?	ɯ�̕W�
���ʹ�_&�~��k>`J�YK��/�]�[s�h��W\��l�<Ō�I)��\Q�y{g�s)w��EC�vl5cD�l�ҁ�K�J+0靖�lp�����v�(�Tgf�@!�;!O h^�DQ]��ee!M�R�ʗ��=���`й����p���������wt�����&�l:b���W�J��Lge^C�����T�.�^o 9wG���X9��o��3�&bȌ�۝��QAP��.\S��P�"�-�$h������ _
����@�}y��r���U�������g��Z�-�L�gGuV�s�H�J;�@݀Sq4����;��R�/Y|�o��:��c�E%yn���ҩ�S�w�p�1 ��3�6�Yȧ*sy#8�&:/x���׸>�Lb3�9W+p��uS�BW�XQ�׮�������%���ѱ���L�����պȆ{'<�-��O�;����vFX��K`�&'���ă=ܺ�H�:�Vo�j�u]�'�A��~"L4���I��͐)��h>���3�Ǣxf�ZD1�4j�e�3^"qm&�����^#K%�Z�Gh�.G��; �2���r��A���n=������]��O^3 ٿD-W�V/�C���鉣�ڀQ�����7UV���|Ҿ��D�;V)rہ�@g5_ :�&��Ҷ�#��b��}�:V\��4�D��V~�H}$�n��c3��5�J;u��Т�0ȉ��� ��Fɪ����:+�
(���k&]��1r��[o������I:���%7��?H`��\�k]��E�VS�|�J�d��\	Iy\<�/1����P�3���Ɇ�P��h�^8�8���W�vn}����gp�ne�`�v������)w�߾D~��>y�793m���% L��O�`GSV�m"^T�

�;y_��䪵)Ųd�^Bgl±���GB�wW��G�#�K[��=��o���)�Em�M���R�of�3��҇�Ih.��_KV��-�;F��;��ģ�ֽ��Q8F�DG�ʆ���[��_$	�!S�͍���Q��'���!.�,!�֯��Ln�!p��s��~�ۜgP/�t)�͑W�LN����j1�މ�����L�g���>�s�@�_�s����q���
03Ɏ����V& ��Q��{�;�vW%&G��������3�I`$��V���k!��D�g���o�9!���W�%Pau	}��_}�ɯ6���t����d]MqC�vC@���E��P����͛���W��ߔ-zqp��<�N3�<���gǻ��Q�c��D<�ANB�X��W�E����-h��́�u������b�?��҈O��lU¤C�@+Uq�t���B1���pH$��{NӶ�o��Q��	��{�j�v�
؈;;���
�I�ݖ�P/���$D�S E] ��y�U4��V���}
ŕ	��Uv�q�YtԱ$���D�}�i�9�KU���y�N�*�7i�n���T�h���$G�k��������u8����\@]wTA O-��d��b���3z��d?�-F�mf����i%�}*5n�`�����ԣ�P�79��(U�>(; �s]4妥�岬%�C
j���gsұF�h����!�������Ƞ��RbL |^�9Jk���S@mueF����A���͈��mW��H|B�7v�a\��\#��J�lp��aCQ�Mdm!l@m�j���A;�]�7{�B���q8g��( ��ʏiT ܈��(w��go����Us�N�ڽ5��C+����(5�R�W����τ��/���Nm�d(���5��Þ)���F��v�O �#$RN}���C����q�7�2�n��r��ZRb;���y������$m�}B�;���Wl�>��憽���#�����ǳ�h������M�Frǿ�\Rd� t���g<����S��^�m�cń�ݖ���?�r}��'�SG��v��Ɋ�A�Z�Mh��w��9���=���S�Pͤ��+��@#�z���d�8X�M���z�'C ,l�v7���D���д������Q8$`�EUqA���vGO8��}a�J=O�&�a*D�@Ƙ��iH~W��\�YC�$�;m��{�j<s�I݀=���U�BË������3��9�����	���Npi��GO�n�t�Iͺ�,����^���f3Z���X��$��F�=�8��@+�Yu��;��;�A!*8G��A̤iiZ���~�8�I�lS0U���WHxT�Fd�O �J�WE���Hq*�I��5��!2� �ڳ����!U��"",ɏ�o-7�Me*eJm�E�/��;�a"�O@�/y�UJ�`�l����GE=k0g��҄�X�\]�=<T{U�f��\�0��W�zO�^�^��"Z!CLh^�Sg�*�I2i��,��z���.-?Dm���;���4U�%�[�kB�Sc�3��H�����z��D9��I,�̌��8-�/"l
}PCv��e�;R�"(8	�d�î/nX[U��ݺ�B�s\O��pߍBB�v���>��7�c�8��;�����X�������IA�����T)TACFg �����Ђ��ɂ�.�Ne�[]@o��>1�jN"��$'���ͪey� ��%U'=����)�=�"���@��>�PKz�4�]���zǂ9��A�by7{tG�n'	�k�}WcT���c2���8��_�MID��T�I�O��>�,�_g"T�j@�(WV=�����n��)�q�����zi��5>a�mb��y��	�_Ak�>�����Z�^�eK� �0]���j)o�C$6o6g5�]��M�Ƞ�u���u��o��!�oI��c�F(���L����!-���φ����#l��nY��wH���љ-�R�%?����D9��:��5j�Q}����m���,�͍�Lִ,X}��y5JǓ�b��Ǭ���0� (8�^�x�C��_?M �r���Ő��"L�̿ۅH �A:{\��)K���~��������j�!����a'���V�
�a��<ˣ���q-��}"�� Eԯ]�?�9zc#�@�������JU��
��g�w���c�3�"�f%~��*��2���ʹ��L��X�A�h����)�m��\�����{雃>������l�L!����Ȍ�`��������ƍ|C.���D��=XP�\G�'��}N2$��&�芷�ݜ�@Q��N��Yq�ȗx�eXTx�vl��B��]��C�w,<�#%emC�gu����َ����έq�%ū��<����U4�έ �6e�K�Ύ��]�RyNKtZ3��d�T�L6���ҭ�NӖċ�����ŋR��~�����[�M���5�/���]��0�E8p;S��}��k�}U���!�/�l?a˨��7�݅e&T�4���ކ� =����ؐ*B_�t����B��X�G�B�%x_�Z0��֨�
7�n+j���e�L�9OFl���͞��+:u	����Z�W��9;?��?�ݩ�B�J]��9�ب��_$T0u�C\I��O���m:/�,H�s���b��Ó}9?j�W���7�W���X��P�d�O�O���֙A�Nhԁ�'-�g��F�ų����p".���C߈3<Q^\�_����
<��{�wо�)\�H,+3:�u��ͨ3y~G��V� �9���U=�Ɗ����p��y�>J��:���#%�ok�����xAU�V���U�H��M�T���̤4�S��S��0Sw�\��*��2S&�s�9r)|!64kǠ�b����bY�X�F��LF�f�ǎ��xt�@���0���-:%+�f�O���*E��Ñ� ���ٽ�����DϧΓ.� �Xf�"�y�}ahU���9b��mi_�g�}��#aC�6�{��'�#���m��b�� ^F��-eϟ̊uZ�e���n�� Zkw�����)B2�@]�P�u*<B�B��TZ#iL0�<���Ӭy9�M��m���yr`�b��JM�ukNm5�\�82�V��F��`�v�H�c�r+8� G��]�'X�iL��Er�����~V�],�+�JE=f����-�ȿz��_)�T���.�8W�Sj�?|�e7J�w vZ҅��4��#d�3���%����|M�h�tޢ>�t�Z���#Osy��7#ެ��u0G�Z�Vn;Ѵ�)��ǋ�.И���+�	��զAUQ��Ps��=��훖��F?�$�~��d�`�VJ���L�G~�yզm\G���f�|�4�I|��.v��PS�)�)��t��� ����E.��!�5�gAd�M�C}쳍�ε�ah�t����K��Yt���1(R� ����Ke�D��B��@&�w�I�b�X���X(G��'2��l����zR�
�Z˜L��\�@�pdz����Y��'/7ɶ�y!C�i'g�'���)Ά�.C������`k�/й��?&��[�wf@N[Z�8*C����ufP���8$�����vWkuo)H�e�
�`����-7?EnM�D���5���=.V��mlחP�C�A�+�3������#@����؛���ϱ[�����I�Y�"��  ��٭,"�x��`&F3*��W�	�Y��u�K�R�{�����KS�1��#�|ت�w���= ���_��dq3�J�k�t�9%���YS�=C�V�{�|3�.c���&a�~+x�U/9��d�U�3�U�o�X�g���1ⲅ���7�rϨ��@Z���1�oA'�.(��\|��}.c-��$�3��:Z'����C�<��c�pX�%���o�{��I�t�
�v]��|�>�%}�W|O��G��9B��@� ����MVr��-e��t�_yAJ�`+������ZI����H$��D-�1�(6�֓��%��f��;�����Č�+h��[��6����K��K:���.{Y\�ɕ��6%f��"��
�$��ȓ����
:o�ЕX�c͠S*����s�����i18���Vk�]�3|سW��������	t�0�71\�'klf�w��=���)/nE![�j�B'}�7�}.�������s��b-�39Ƨ���Rq<���2C�(C��/�@T��M����C�;�B9�=r�h�^�ϯ	벨��6[�2���)�A9	|�8r`�	T����ϟ�N�qB�?� ��<���ܲ ��0h��҅M|tn���ıIP�����N6yFՃ2>�x]KY��S5����A3��Um!�P���Շ����#�dޣ3�nkr�f�WCе����&�֥��K#���d��tR(�� 3�J�����^�4D� X�$�ַ���G�x����[�Ғ��_H(����e��PZ���n�%і�~��Z��h�<�؞�Q�9PLX����8M��F[7}���p�
q�c�r��C��c�l"���G�"���]��j���e__'|�M���9l��ԛ9�x=��`��i���_Iy'���i�i�$�Y������˿:ʉ��44p�}g�yǝ�� �HI�̹���g ��m.�%E�<�fÉ��'�yѿ����Ү,C,Q���;�J��ӽW!��}̋&v��d�I��<�c��{�@M'��J18_�R#tP�@eeek���Өm�"��a�����Ns����&�
�.?948$l�y�e��F&��"�������T���
�������d'��4Y�=��+�yOS�<�,�e��	�P�����G�wK�z��<�  �.�8U��;[�aȌ��]�C?qdU��
�{c�S� >�TrJ�-�'K���!�9��)o���w8�χ�F��f�{ӟf��e�v�"U��[���ߠG�qz�H�Շ��FC��M\�ؗZ��$�c�����/��C8ݩ�HB��w���!҅���y��+Ο2M\�R�E�U�;{u}DV��*�.��sM�y��Knj�ie"�}od�XA���:;��AQ;�]���U7ܮ��VW\�����6}��B�LF&&�?=�c�7�t+��GI}����A������"1����u�Z��M6"����m���/��_�3Þ�������gǴ�i�`��/�7f
�~��,����/2\9N��u���u`,J���J���������S�z���\L����qAk�\\��>-h�>�+"���SN���|8J	�@��7}	�*~��nz�*K��l�s4�v��ǩ�ԙ�ҩxw������k�V�bG����᝭x&�D�&����凣���`r���h�\6U�������'��߽�ʓ�l^[J�.�	�b��3Ɏ�j}�v�.g����ع{����L��F���s
!�L��ME ~�դ�n�ݿ	�`�D�߈�ۼ��|R��=T��������n�>k,��}Q ���D�ͪ,�t�J��M�ڒ�쯫��t�i���׬��N��)̆$�!j{XӉx�R� ����YjzCZ��G��I�%��q���qU�jBL�;O���C�m�M���bcGZ}���i����g���٪-vx���i�N泆��B�A�0�X�19֯�1�nO�{ţ>?�UZi����''�;O�W��AN{���-"���m���	�a;�o�wU�`�r0����`��nh�d�݌������������њ���I$�W���m�I�%��� h�A6\9��G�<K�k�����@���G�z R ��O*���U<%���0�R��ЗY��'J`(��1_l�����{L��;�-�I�ga��s*�-W�^�g�_+�ei)Oa�G�Y#Fj./)��ԥf��e����`��ID�wE=W�/|��v��v�C�om�ܨ����cN-y����#Ϡ��`>�s vHHol�|h:�K+HM5<F��c̀�9�Wy<�7ä�Y���>:GjJ?�#�,י$0��6*�K㯷7�HDn��P�s��Qp���ܬ�v)���R=�����虓�@ �T	�D��m��y���$-(7S���I��1˅�ќ�T���.`�|�"�lp�"��8�O�X.!�4e����9t^��`(�����=��"ظ�r���V	����,{y3��FH��׿�1�0�z'f��?h�u0ٌ��ԟr2s\�_
3)4�>�t��Sd�Y��}�#����8_�φ���G0�}�Û�iB�w���*��� ��Z��S$.� wԼ��˛����S�����P3��`�����vo� �H�ZRҽb��f�σ_���4�
_�6_è��H��%��I]�\;E!��d�=m����3='�Uq��)�P�諤���M
��X��uO�����%`54ѻ���]��;׼Ȅ���rHٹ���]�V�)��%d�| �ȟ5p�%�ekjUm��(0|��ր�/�i�s��d�M+���2<�j�����C.�{կ��ӑ'"�:���������H��,�A���I���x�LAtm�;�8O�GT�n���h�O�#B�/�3��<^=�S������p���--�9��|�HnU7Fr�28�OU鏲�?Oo�](��S�9�X�P�-�i�f�~�K~:�BMŤG+m�<�U\�1ӆk&�<$�Y�%�"�#���tj��_�<�]sf��$H�}e(�VQ]/|V29%$�Jy�����gMX��{�+20�o�-�����zX��y��o��$A>�C�3<�g���:\O�����Tq_�qU�)�{&K|Y�؎dښ�v���l��I^�
�e�;�E_�a$�m*�Nt��-��b�J�2���H�*��U�n����B�w�%zS������_�po�q��C,������3�5��B7��Fp�&��O_���c��\BO8f���3l�֍3?��qK��Z���Zo���B)
�+��c2�ڠ�`D֛���R��eQ|y�;F�͇f���1��^��|�3����S c_�6�����w}t�2̷�]�3��萒���s����o`gv��N�c�hەP��[�鷺�e3������0�>c�bҦǼp$a�]�.�݄��O;�Q@���d9���h$�h�x�l5稨&{��j��L��49�w��Y�[Ǩ`�&,�����p��F4w���q"�RJz�\2$�0���z<b��àTW%�>��ǂ��bI�xv7�E�d�#����*�>��ŷX�rg(lqA��{m0�}�@C��)�v�(�H�Y��_�:��f��%��]%����̞�Q!�?�Gk�Q�$hk���^a[z69ވ��_v��[��KqW�)3�ji�H����l��H�WU�TmG�����������L����Cn�qL�["�7��f��A�M�J29x4����;�E��x��!�oA���t�����=*��^qX�+���~g��,70X�$NA⽝�$�]ñ�^�u^׀1
h�W��X�c){�M��۞�=��ս��R�-�߂���3`<J��B��v�$X����Q�N���V}������Ȣ���Y�Z&Ӫ��* sI������;�-�l�kɄ�������	�],�E��8�`�a��3�ql�QĴɼ���������1���Mtȇ��)��F�� �Vcm;r,Q�gݤ""�&Z<�+p�>�6R��`§����^��]ж���L���U��a���$*@8����Tm��܄���"��w"�>�w�nKٖZE�x$���|-`��di�t��~2I�=2zс9��yo���cN�[x��/d�3������>R�9/�Z�H�:���O,5��x\�I�?�MׇIEhK�?��$��#H4"`��ȍ���ƽqq�}�`U��9�I��'v��t�i��E�tE�8�'gx�l��|i���%���2�q|�r��q{Z�mS����Oa�����
�\E}�-��`���ku/1]�R����8F���W�In�G�����>
l��!�$�QB���u�D�1����1�t��ᐶƣ�g�����_��1��8az�\����T��Hg��eb�-��G�w���JoB��w'#.Hs�����k4�t�Ϳ]��ް½�W[w^6/<�����u�� F~�!k�bPsJumi�w��Y�"�00��\?Ow Bzy4���O���*�A]C�"�#��gO�������-�vђW�͖�����gЂ��tt ��V� �+��- {+NW�� gM������8����{�(����L���L����)�u�Ye�NU��Cu}���b��m3"�}%*
�Gwݑ6RR��:F\������������	U�OS�4���q��n�k�NK�6my�.K�覧$�i�_ׯ�)����#fOp}��|n�.F_J�2I��UX7`�G�&3X�誕��5_���З8�Z���)����o������<��d�fߩ	Й���o��`:�-)h���X�`�p;�ูA"��L�L"���;�"@�[
/a���#I�l*�QR<rt�[B��D26��9��t�X͊�юt�H���,����_+�V9o�
j�d�h(	6=����X(����t���l�um�����3�X�{��nc �cF8��p#ֺ����,ٱ��!�
`�D�p�ҸȴwҲ��n��u�K�
��?b��;4pC5��ޫ
�~��	6+_�<�qd�fS�x2�p5R6�H �
V	���O����L�r�z/8�S��r�$@!4�Bw����z��@�po�-�pN{����x^;�4���GT�� G�DE�ف�yGF����C��X���5G���_�`�-}$[��+Ϲs�by1b�s��Umpr����]6�8q��d�c�� ���y|���R+c��C�2�������R ���.��z��У��&1�q^�<�Պ�L���kI�d�4j�!�xZj��@W �>apJ�d}V��ÓF]�-B�~nv��;�#�;q��u�7��ZP���-~[�T0 H���Na��\�g~ �5��C{]�0zVe(o�:���EPኆ�)�J�� �XzM�T7'��U���e
�1)�������`���'�ΈRMO�*�i�@�4&	v����/Ru͢;��Ҍ���wQ�F���3}���p{�$<�YKc3X��+n85еԆQ5�ݵ�ss*� �q*�}dh���D���7�\wRߌi��>oJ)�x��1��E{�HrU*���̜C����_�a���@Ƽ-���h��k+��@���p��%5M��@0�d�v�+���j����B���)x�Y�]Mk�b��t�7y9��h��@ܵM��O� ��(ht��*����/��6t���,�`ۗe�r3+��Lmgo�<���(���Ĺ��ǣ��U����5����r�{�+�Q��Me|.��Q	����[��/�F�E�d|��&_H}i��-��@����4�ꧨlη��}����������&�,�*9'<�d�O�*j�p�Y����d2Y�h�X�֪1��6P�;��=���so8�޳�d�)�Q���_����ŝ+ɥ������f~�	tZ�H"�z��%����X^���F	Z��B3x �K�f��f`����S���!��ೣv�V};5����m���;�6  �
(���q�nh���.��潎-�r����y�o`�@�9���9���� �Zz����K����OR泖asX���.�6�'�+�ˉ�cLx~�w�V�ev��Ny��c�Dz9To�n0U�8�m���L�㹢l�_8=��4��m�5!��#�-��ߐ���~��e}�%���P��v��j�BPeM�6/���������'�~$��Up��}&�q�<�e{��
q�5(����{v����Wd���o�X�t~1�#I3����hh������˯�낈��'�
�3a�%'�K>=4�mF.[e;�/���1�<h�4��VO8��I�j0�G1(X��=�Ӂ�f�NO��f��B�*^�\z n���~Ÿ�#�J���^��\S�}�lzE�༬,
��[p�x촕��o!`=c�Մ�7���,̀9mu�=�0�̵�rem5�����.O��MN��m&¼{4'�f���!b��X9���Ǎ���^|�8�,B-���A�VOH�L�10���Sو �\��z1emw �X�R�V\%��O�{�BK�.T�Ifz����)��sOr�x�b*dl-�1��I��ؼ���x��EA����RJ�o���dД�:�$B֋��OY%x��~ɦ���t�\��J�P��^ 
�'�<���|4�6e�Tӂ���S,)~6?ځwV.�٘t�A��D�}����+hS"�C�.��s�����Ͼ�rd ��|��}���	�I^����I����t��	~W0@5gy�3l���!^�ᣃ��6�F:�$O��x��n�����w�Z8\����/��(�S��e%�vXǀ�u��¼"Q��;��G@�	̹�!�<��˂�%\�	�[8E���=�8�'�q���l/��ig���H�Z&n<�J3���`#��NJt��T���E�
�ʏ���1R{�I�j~�N
��N{2{������-�����W-Y͗H#BVRn����V��-H3�H#5:�� ;k�,Vdw-9|�q=f�K�G曑��^D^<�VLQ�l�n���M^7�]2-���L�sD��!S�.���=��P%��К&��ʌO�h0B���'����=�C7��k8Nv��I�$JM��O�e��]T�t��ʠA��t=�%���.�Z�_��?C�����?6�C���dzH�=�:C
9�柜M�I�5	'���
a�o����e�V�����������m,-�u��'�?�Rx����0�{hj�H��$�"c���7��KP���yn�8��1mb��ˇ����l��"�bd����m�2��o�W��{��!��h��H�D7l�@ۦ�c�eQ�K�a|����'��vP��n�u$�X�ٱ�
O&=�k?��� ��$��ڄ��VkFe4|�k��E����������j�&E�Ĩ�XHI�S�@�G�Ŷ@5M����dH�3�@!�R+�٦#K���J�3F]���Pa��� "�o��G1A��/]�>�J�Y:Z���o5>��=�J�L�4�+���}̱��7��3O��h���A��i�:���0Z%���&�3��*�D��n����f�{*��f��O
1�oꗩ��Bסh.ƒ-\0�X�
f�{�+b0^~�0VR?\�����q>�V'\��u�>��x��<|��+�ف�D�[=��^�.T��:�V=�'{|q7���n�1�i�-/V���r�4dJF��P�`~-Z�=�cE���_�N*�����i���3tL�I&���
ǼI��ж�*+�w�'������]�s~��C�Ĕ:�u�쵎v��o!�\��3�U���4��*�O�@	+^�V�k�(Ts�:����Fp��y�5���T7>V��4%��Ԁ�o�'�-�/+�B+�j�#C�&.%n��:�:əm��Z�	[<;D����f��f=�%�ѧ�v+��ޮG.��:��ݶ.ȩTae�T((.l4�V@��#�8�Y8�~Ena�1��p���bl��ϷM�6�jvA�x��9�CL�=M��>&�4�D��qmf�-d�cz�d&�IfbAp�� "��!��	l�����7��hk�b�5���y�lwn�b��?��ʈ�>D�1G'��SƟ��16~�kgx�����P.f� mH��.�������Kk��MY�R�	�ik����Y@�^�a8RC�6�C�ۊ�L7�%�Xm��O��
=:
��)��p�{�^��)wۨ���wo|�/��|RT����׭�TR��*⍴e5�TKQ��N \$��qT�(g��_�GB]|5>���E�ʛ��|�=t����'�����-u765!*0��]�y��K�o�n���S��'7,`�$qX��U���۱�Ue��0v#}er�6�u��[Nr�R7&�l��kp��/�u����)���V	*S��ᚽ�^̮5M��@�1��p��4����	������Y�b�j�a��mQX����8��é	����s��FE�PU~����"�f/�I�����"3[?T����E� )sq}p+�.
�����Mz��]�4���t�	c�u*����5E��� NO,�∂��zL�6�k�KX�
�_��EP��b�g7��c��J�#�0W��1nn���[��<&+0�J�Ynevi#��!�pzt[s�ub'k�h���#s<��ߒ���A��؇2��v3�J4��	�t�Фj/a��"�o2��l6�M�Asm��C�-�x�b�m��f�M8�C���|3W}�S4�؄S�E@e#��T����'XlA�A�q,얉UH�@��[�t{;*�H�vaw��=q���_��;��JJߠF�2���'�w�_�� Xԓ��G�ˠ�b��ٶ>�<�T�V<Z�5�ƒ�7�ro! ��P֗uM����q�[�W�.x5;��{*���+2���wJ�m[�������0ϕ�&�PDe	���q"�����U3dpy!>�^��K,�
�f��,�K�eu=���1yKR�je'L��3R�Z^;��嶎R4b�`P�%m26V�2��������eg���-� %����%4��O��!����+��kH��ܵ[E��4ΐE�}���Cd&ȱ�U=t�Xf��	u��VgD�[\���P�nq����n��pGo�x�c.K ����r�?��`�"Pzq �d�6�<BY��6.��􉞾�[��ѩ�q�[��D~����r
'�Zr�� *�Qb�h;䘗w�Ţ��	�60Ѹ���o�}�6;#V�?�$n����]��R[��l)�E�wW����]��u�z�� �*�S����6 |��nK ����a �Z!S���,v�F������8�sze�wc'jR�ܤ#���]�f���Q�g ��	t=fP��K���Z��F�	�0����7���8k9��g�Ү۳�Cm������5�P�GߎieA���;�E pl�,���j5Џ��]�T����3�/k�aG5�n��JuoiR�_-`��^_�P�V����?N����/����p<%���r)��|�Lf?�H\���8:�L���Z��J���.��i �rҧ�w^��u�Y{Ӕ��2�<G�#�Oȡ�6(e�,R�O|{��}c�Zô�o�e+)�&a*��7�Nf���Q��0:�2��/�W��i�L�Q��4��K��Yټ�@".�5����G��IQ/@�>�_BW/�"]k:��(��V�֑��>g��5�L�6폒��ʶ�2�:4��Õ��j7���)ϻ�v��~	���|��.ؿ����;��u_뱿����ȯ���U������.`�FR�/����7T�����MA�kp�W�z�,5�V��y	d)�^?,��"2�VPȟԱ��K�z��i��m=�("m6����S���7����oI��v�xO�^�g4�(���p�A`�=��1̌�9���
̌Ŭ�����L_˳��]/���i�n8�>|64���%΀����d��=ޮ�I��Y�	>��y�Mj	�\���ϑk�-��fJ�}4���m�63Mz���Xs(-�k#ǳ&�������A�$�o�5��-���+�g~�f�8:~�~Tj=���PW$ǘ
��:=s{
���zv؁(��ʤ8w�<�ͲQG��`���pf)`[�ot��T���O|�7S����lJ��,�Y"z_z����KO}�1^m��:J�W�ܡ]�Z_H�:Zr��O�+k������b�����0��+�T5����80�LL���4�Dj��D�Uc���f����.�F3�F��d����ҫ8��B�>nP��=̯��)�:��^B���Ŕ+8ō��Ϋ]}>/���e׋)Q�YzL�7yh�/�Pph���������Y���"��ί!ڏ��þ.�s������S���6s3���&e����R�/[8_����li�C�z�2ʰOD�D9�i���~T-;7	6�<6�ΜS�s���j�����n!NU�; �>p�k��j�-72�p4e4�c��Fc���4t����Ls��'hԙIldO�:����#c�\n���Y�o3�	޲xBg��MO�h���\7�n�Ɠ�#F��OC�]�M7E�Ԋ���R��gL�����!b8�4�����6�1����풱s�jiӰ�FPnQ��dxA4X�%��J$&`���X����Է+m��,�u�;��!&^���M>կһ����L��O	�l�o�<VK���,dnW��Pԧy�|�z0�ܡ�f�xk#��\�7x%,�\h�*Y,O8'Y��S�Z�MZ�@SJ�4ld��L�2�8c�\4Y��{�BncYƴP+[sz>]���)���Sf����68yc�� ����]�0ޡ`�p=�NR�u�^����[��N_��Z�Y���"���hy�&~�z�o1؝�y5�f�[������A���-7(�������zї�ix_�v�Rg�n6���
��?�:��0A��Z|�b�����I�@I�ӭ�����x����D�X���=��3��E�B]g�Yh��~����T�}��� Í}z�dq9�jM���0=�8���< ��O4X�FW��s�B���<�LA{i}��ù��j���6���=��CО�T�8���#B�@v��U�0/\��T�<��fr�	��u�}p�e�>�x'&jh6�͒7����_|�c��3�V���Y��O������ze�I�&G���!���ƣy��
en��u�S����.�$T�Jv�)�s���2`	��,	�x������a��b@��ȑ�O�l.�DC݌`��:�,������/����#	;��c
��f�y������f�e��`�!a���_}}b���������Jb4��هº;[ ��}o����*����|T�?WnQ�wV�bb�p�rSS1S�z��{_(��o���pk�_ӎ�:�vfM����La���V�$K罎��bLJ�0�<��r�nk�d�����ޝ�g1�/B��^.{2E7$Y՚��#䲎G�����o.�R�����@���ڶ��c/�y��-F}�J�O��L��2vm!��+7�9 S��k�-A�"�|YM��~vؾR*�y%������5��C.���6���&��j}I������Q]���k��=AH~)�ʍWe�b�UP�5"�T7�j�aY�] =n7�M�>�y�S��}�)�p��H��}���e���B ������+����y��jhjs��;|x����쑒���G��9&�ڴ���k�9��CL`��\11�K�Z��6��Dݔ�م��	�]�!�v�U�Q"[��v���8�Z��0�/Sȕ~�v���������QX�\��ٜ��k�+%%xCD�t!w~He�M1�+Z�)�*��d���)Ͼ�o�=���u@ls�Ĺ>�	΢�8Ӄ��-,N�;����yo�,��翬�S9�a�F�k������XP���C��PXG}(�A����nJ����o�,Ql!�'�W�zM3�7v�A�zu�QՊ�I��
Q?��$�����)�$hG*�Gh�S������~$v����(�PY�B�Y��ʋ"�|��m!�� u�1����Œ{������/�� �r��F��Dg���A�S�Կ��B8v��'��Yl�6d@�x`+�Wᦊ���
z'khT7��`;�~ht�s��=�B�O��4({�ksP:GV�>)ݔEW/ج��1޻��(���o�8�c
���
���7�^k����	B�$�����͟��)�T�'�m~|���p7�Φ���NG�{#�2�x�S�c�dgsʆ0Fg���<!7� <
�C����Kl$9�"^Xw��х1QO���^��nƜ��A=��M�茋P�6(���8�
]Ҧ�f8���_�������ۜ��n�b�M�k��L���3�?��R��6a4m�]b<K
���S�'M��]�s98Y$�+ZC
& ~�`dA,��*4��+ە���� y��'���ث�$�`�yؗ<B[䔠/*"�A��8����F��� ��"�=��k�߱�/������x��c,��4a\��S���6�=�Ù8��p8\������'ڣ�,ؙHhAؾup���)Ը�s*� �:��Ъ�$H�ˏq��R��n�ϵ�F��=<�<���ㆲQ��'��n(W����d��<91�#0�F�U..s^R�ځ��yΉ.Q����o�n��Xw��lBe�I�����x� �	yӶ	�X�G}�e&�S�B��I���r��tr�{4w�Mo�Y�$e�/D���S^Vf	�|��3�ї�����������^)}"�T�Z�7�w<�q�l�Nf�'e����};�X�3������nV�լ�߳T�%Tg��&D���)-�2�0\:^С�l��#�r��B}B˭=����m��?5�H��ч6�e v1�)5��A5I���bKlb��tB7����t4�l�%�膺ڧ׺B�L`�|h7�U͇��"��
rY�����5��aA�D{Z}Fl�u4��F�e�6B)d,'�gl���D�B��E!��Lp	導��D���}��)�'����
s������AA�G�a�a��6���U���Ei�|Cf����Ja�+=�x]�
���εy\%TYO��l��%e�3Vp �K��~!�3����y�$�D��6��̌�^�
Ag�A�2o!i~�UW�'\�j�����3��d�i, ������ \Cz�t%6˨{�Pb{�´ɶy����$��1}�S��	w��D��{>8КEV,k����H�)��5���l�����B���J��.U��rp'�iP�?�樮�2�b�R����u*?���0aFޟ��$1N�紦W�P��|)�ӵ=�J���zFS��Xfefz����\ ����1Oً��צ]�(�@�0m^O�8|�1�r���e��,|ܧ��i������Œ����@�L6�؆17;��al� l
b�jN�E
�(�HFäX'EP(;�s�'̓D g��G�%=���"�v�Cr���,HD\yː���_�
%��L�P���do|������ZE��}�5�!��c���`����E�fQk?��1�����?-�6#�j`�y��;G:�jq�|�-��yl��?SI�*0��;���>����v;g}�G���PT�U�U���iߌ��#jkƱ�S�}:�Q�ݣ!�a��)*k�c��X��ȃ���H�Z��÷Oe]S��	w�E=��<���}���$�|�o�3͂�e�ñu@��vo~N1$�{�vX�ՓF��A%@�]F�fh`8T��\�ĝ���Mӏh%/\����z���ڻ��۠��V{-�.F`�U٬f¿��u�����'FN�����:=i���6�]�?��9�rA4		a�H��@���ED�Qe(��+���Y�wte�J�[�R,�:��&�a�ۋ��kr���T��PY{���=����ߖ!V{<#EVHϸ�D�Gk���1���FO���ڮT���D�¯�T7��#%��ޯ��yS�j�8���������d'$F�Eh@z':���آi���+١�b�Ӏ���IM~��$���'F,
�����-��ޏ?z��c�A�ML>:gT�Ͷ=�iE�}��ŮѦ>�Ի�n���΃ 9m�mn>��}�|E�+�ǩ��z����<V���>l�,���~M��Θ��L���^���.�!��1�I#��)p�:2Rԏ�t��n��!-+�q?YQd��G����
qP��$����s�����~{N~��7/��B�q7��P��1?���ZP�xVyT� ���C�Bދt`{o��CX�t�$i$��"�]}Ԭ��R�p!bWp�ܾ�b�ۧ��@�ؙ(��Kǟ�'��>�ƝN�
�i��ނms��er��%Bd�s��m��"���~�p�x��t�}�>�i8�Q���� ���*��v�frC�%�ה��7[�F֙(K��e����B��压�&��%/-�Y,�@�_s�kƬ=�-��Fw���.ڧ�G��9+��,��rfH�t�Th������z���g���d�6��ʒ`@)|:w�k|�����Sb@q̆Pq�������J����Q^σ��#{��g���˼=�Ty�:����ɜR���she������ݼ���p�	�xwq`�;�0R!MK�A���qy#��tU$��i��>t0C�u�^+���Xʇ��|�n��#J�i�r"0NU��J&�g� ���%k��׎�hGV�����䂝r��ĘV;��#�u�+(���Dvop;ud�GO|��Sl'�r�Θ�!�e��oj�<��UV��ۦ�.����[�w�(c����>w�V�_�:TU@2�@YI�%#�q�6�U�WGx F)`l���m*+@��d�c���4뇌�\>1.�g�yPyݥ�����/b���a��◤v�r���O�_\���= *ʬ�m�Uh�(�}��0G,�2Ek �`�6��oB�]F�[܉V\��O��^y}cO�P�LE�:�/�r�1�i���얿�\�m�_ˋ'O�h-�t�ؗ���#n�n4�)��[�^DR x�!�4^����m�1f�ƤYrY(@k���!��JZj^���~�@��GA��v��g��p��rK��xwu?�B�^�n�1ʒ~"�ޒ�J���K`]�n�T���'hR�)?/����2�����n�q��U�}ҕ����㥤���8�ؖ�h�'<�L���$���!`WjB��G��6�� �ӗ�w`NŴg9t�P��P�+���1z�gm]=F��w\S�8'v�@ؖ]�I6`r1�����'�����[�;��3���L�W���#Ʊ��*j.$��"�dls���VJa�4.Z��Hec�p�RF�a�����:^��Q{�۩�`���^�����Q�u!��ܙN�����nP���|/�_";�#k�k:>Z8�?���In "�������4@ �}���\���Ky��!��.D銍�����vE��R ��9���q������yE�5���er�
��^Cg~��G�J����	�5���Y-R2��m�]�=8�WC�*��7ŵ���u	P.0��?�^y�ur�6L�8���|��M��w�vĬ7�n� 2��D�Gf�-̋l�W�I��fU��4'�����2j��嘸��۶�]E�M���s�����Ks}�iz'Q'X�"1����8G����U��ڶ��	&�\[e!�	$*	���?���b�l���"��T�&�v����O�^�x�킋ۍՕ�v]'8'u�d���4���u��)��d���]���ʄ�sGV_8�*�#����8��t5a�R�����AaNP���H*��UΙ+Yh/o͊�Sc�z#^5�Fd*AX�\[��)��� o3��[o;��R@����o�ᒋ`W�u��\��Q!��H�i�SO @F�lG���@����Ϙ8c6F:�\�;=� c����i�C��w�Xnt�X�<��ְ��ɤ]y��a����a�BE�D���v��x !a�w�wa���zѱ=�g��'�� ���7S�>K�U�O관X�p�^�h�'�O$&�q%�3��$Ȍ{�9\7��3�2d��B�Ó���Ҽё����koI���d�.�ɲľ�	���ν&�2x�UU>�8�)*�?�v��t�-�E=�=�}x鞌U�x���F{������^�y������&�`"�p<����� 3�K5�{��=�[�,b�=kE�0Y�	��M(�X��=����dF8� ��A9����/�zca�� "��*w�4�S_��nF�j��l���XMQE������I���� �-��˨{�9�,����+�i�g��҂��}�� H1���C\t�Z�?��aX{�W|A��>����C'UX�FrE�2�-��Ϻ�H<������C��LQ$���L6�R U�*?Z���/�#���^��C#h5I��4਌]M�G'/�)�:�/M��T d?��$k��F�&�k�W�=�ؒ�|�pZ�`Դb���b�jͪ9�b��_a���J��J�jhn���s�hCN"3�B���Fx�]~�t�A8H�z�E��G�׉��v�����s�@W�{��VP��܅��<�]�I�E#>51��� �{j�u*�Q%*��7�q��ߠ�H����$�{��Z�iAcJٯ�Aɔ�V��qLҴ]��Mh!JR�̎�o���t����5Z��B!ښđ�@���n?���8l(�]DS��v�6Xi�C_� "�.�qC��-��?+�5��L��[�&3�ݴ�[c$;�_Kt�L7���e��C�:P\#;�b8GW���X��l���+Cػ�iP�������Լ�	���b��#g��HK�1P��l>�����C�jc|wB�$v��e-��0�V��)��.Ƌ}��h8��Eس�姝�k�����ߛN��C_�[̯,������_(�mEJN��٣����3����i��K~������*�,=3 ,���j����y�L¥za�3�nm*e2!ܑ�b�A�^�+F�;�6��K�}��=J�u�>*��� l,�c鎽?ꘔVJ��:8O�ocR��nb�CGT���N
���o��a���$�U�z\���ګ'�9��<�oZ��Ī��_n����:�,����v����~ֹD6T�A�'ߢ����oи�Ò�s�	��2G_m}��SǞ�k�<�~h���K
���H=���L]̹Kv��`���Շ�"Ęﰹ?z1\'G"�	zy��=�S!��|���H�݅#���q�x>r��0�6xhؽ.*'ErĤ�4�@������I��]�2��!H��@��)���0
�wJ��_�b]�hƖ�A�T	�6��@����ԍ��M������5[��h�d[���<�?4UD0��K���7u_���"Mp�T� �]��be2��,Ȑ:��11Y�~�6{=��9M�+���$�GH^+�(�� 1|�Z�R�Ql�o�?h���S�W	K�<�(h�Kl*����laEA�	�K�����^W+w`���ܽV��N�/��Hx6�7|���~Z��	R���r�h���%1v�������&��P��ڃ�5G}��bwOW6<�>yNl��-Gο� �o�F1�|����r�\���r�87����tt�6�=����Xs���>>0b~�V�X]��/Ew��-�FZ�-�d��3$����O4����FP�L��X�*7���t�xl��'���$Ul��;0>��`h{�-� I�x��~k�
�]<l��1;�Z�6�lKH)?�����q�9%0$+�J�����+�\�&9gQ��k)��W|5X>@e}�|?��z���i��&}ڞ=a���#�u[i�xD���;zuH���Qײӛy��^ӗy�>9�OM+x��-�b
G����KUm�]��xڳsfi�%]lI랪<˝�P����{�$4zz���N�bv)&�&k̖�lQt{4��DCJ���V�dq��Mu;rW���ȡ�b[U���O��'e �K���p�P���cx`x�	�Oc�������T��ru5�fPU�9)��Q6�9��?O2�e�*B��c�J�n Io����Ņ�q>��s4���� -�]�~�]�������	�Q>-�0X���7\_���4�o���b��~3�EO�C��(0.��Yu�K����|;
���g���ձX���Ǝm-w�%E"WaW�T�����H;*�#P��a)�^�\5�� 9�}�?�&��1Ƕ(B���~�q[��K;�3>/���,����b"8���S�=����Tl;'��1|(G ��-�e�'n��~Ol�}6b 	�gc}�C~��}-Y���}��x�i|��'#��Ň��=,q�pȨ1	��-yN���bB��Z�Y�6�W��K��4:6�|�+�l�8=+���}@;'�^�x���HXSTE�b������3ҳ�Wb�a�퐓����18iOh�e&�b%��<ye|��j�T(!]�3>=�&��
�ޟ}>��g���;M:�l�����r=���P��jG��Xz��>�W��]p���ԑS���Q���:)k�����@0C�u ��R��8�a��'�@�Z�cs|e��T>�R���{�|���m���/L��)�3o���������tGf!!s��h8�lH� �{���h����)Q~�^�a,�Fr;x����s��Lڂh�]�z�6~/h7������e�����-���؇f���,a�o�FjJt�B��7N燰L#��*�B
&�Bo�����ж�,���C�I���?ה�z){]�@GI�+"��ߞy�I6n�y�7ss�{��QY�K�@oX�m�7�U�0���vx�D ]�̼�|ް���T���b;l3?�8�M6d�V�׀^�X�{��T�b�ha=#~7��?V�M�65A�����u�o�:4W�Z�<�i�,�*�n�������Hю� A���]\D!���)���qq+/ESr���x�Ta�����5`�!rتz����Ǘm�4<�M5�,�"l/��L6��̰�x�';Y� �����f+3� ��Eb6�������n�w]�C@�*%�ϔ��m$��Y��� ���)�)�����ƲI�������Ƚ���>�y^���4z,4���CX�!P��u��fOX#"oЎpߏ�F��L�F��;V@�,�ߘ��E��%@�w�����5�Թ^�����P��au��}o5׼͑���߫�;zڟ�0d� ȓT��c��n�������s��pqZTxY�1f��7���I0y@}�ϓ�5E�Vj�$
�A�&�8�x@?��XS������6,Q��_&���|`cT+���~����
jن�4 ͵!�[�x�R���ׯMډ��%�א,�}�v�\f@�9�r�F�i��t��-#Q�S�Tp��$��8������,$��wvºO�e-�"�$����<�U�I�lI�%V�W4��҄����5�S�|�QH�ι�W�8o�1�R_0|�>�	!Q1�C,���G���~��sd�݌���������+,:���bV[�����������I�?���������A��x	��<��sc#��
l;���W)�d�����ϯh��
�g�q IH�������e�Q@%8��Ƿ�)�0껓r-�e�>��X�b'+K�	JB-P=X!�zDq��~�v]�3(rG2��V�M��/,o�<Ň��J:��h�tr`�?z�2n;n���d�j���w����1G�����{&;ߌ1��>@/� @f4̯�S�(��p�/�x�-@;���3����L`/�x��iQ����ﴪS;�l~<�
/��B���'�з�����5� ����~(1��5�/����D��wDh$愮L�3a�H��OE}s��׊�48Mh~��J	�x��v�����ʕ����!kC04�6FKλ� �d���5,{�8��FN��=�hN͹��V���)M[a���p�rU�Io�r;s������X� /	u�+���!}����0�c9��Ғ��?v:*H��3-K��7aD��K��	�p��H�#�maxV�}�3k�8�~P�0���~��ڎL0yaXu���A;2�������捼��{.�ȳ5	Ϧ������Cu�"�
�:~�ϲŧ/[�{`���e��Ҧ��#�fލ�K9�C
����g�R�wk�z�"���$
��&�a�_�|揱/�S�;,�+k�������ܠ�+�;J��|g�T$�%TǶ{2�qS�2�29����CY�L�7�T;��T��r���r�w��r's��P�m��'��)4��%uE��ˁ��9����G2"�(UJߊ"����{�/������	�'�<�y
q�{ɮkR�$�8e��K8j�}�AU�?�"ӈȘ���0]�a��F�Dc9\���M	���hχ֜3��d���2SL6 qKZc�O�k���I߫ÕaC]Z�,�ݳH)���b�qj����8h��1+L�b�4��2zw��J�C8�rw�����1A	�Q;+,��׌�.l��iQy�g]5H?��������jRu�j��9��c���)	`�������U���X��� ����C���"�2Z�� \��J��ŽN�|��{����$ fӴ.7�[�am���`�*�γ��Y�a�ﵭ��eێ���r����5Y�����-���sP�:��<a(+�=/_$'ъ$���D ���į�����1��o�ij�!'����,Q����_7�]E�Wo���x�'����d��A*�j<��K�S�ABR墋�h�8k�˹2�{B���nޚ���w��,���r��L�xS��Mq9��վ/�?>�ܶs�9���h" �2����
�y-��7�����v{��o;�Յ�EմV2�q�?*VF����X�ެ�����qG�k��n:����RPT^(4Aw,��ۆ���r��� vM�9�����m�6�n�ӧc��d�����)Y��8c�k��U0Ե9��N	"��`r�퓿AYէ��2(D�^,b��",�G���zY�婜\���<҂�si���n�J�.��~�GnЏ����XW���A��g8u_I!,jO�B����
=s�jݕK��)�TA�y	��/��^݃74i���%�h�:�V�'�!��z?d�K�3�S�*�-��/x��g=vg��s���>���a?�9:��,�#�Ke���Ӛ!����MQ)v���«'��y���j3�wk�M���!�@����SݸG���l���W�Ђ0��T�5����8��yU�|0�
�qx��|\q��	���!큮��V5~x��(@�0��žY��31��;�Z�*.̜Ю�%��3
b����<P����j��E�ON|A�����z��9�9=���9
�-�����.<����M׷�`�^�é�D�٣)�U�(��eZ�5z�;�A#S�!�-2t	'Y��Pɝ�9(���讈]d~2m#�*/G�s�Y
��6op�7j7Y����YA�J�p�@�QFG����Ƽ� ;�:�#��lp�J�.2����V����_��2�Y�
?����y�}�NlcY#���sމ�\0 j�o�������by�o+�%�|� ���z�4@|B�вt��*�K4Y��F���"w�}Z�s�;�Q�va�!|Ruf��$�(͢?�UCj���#cy���~Z������+��p�!�::SMvKw=��>`d��~>��^�vS��o)/�a�;շj���<��Ȭ���D�`J�N����b�N���.����~���"�pn�����#���O���G���G��s�eh�����+O��|<�����J�8إ͐f�I�
}K�-�X�Rܴ9�/��7�?���.��`"FV|�r���-����۬h%��y�p��Z-�b�F�c@[����W#��z�[�t)5٨��~�o�w��۳�(��hv ,�|��e�}�㈢!�f�-VX�9�y8��ׇ��"�f�8Y*��w���s�4�Zߠ�U5��Zy��7�h>;��艜P��T��vGU���D����,�`۾ˉs灼�	� 52�ey0]���j�-%Fo-U�9X���I�4V��,�Ѥj
q����0�b�*$�')��ƸM���%#��|$&t�>�c�x�r�/nO��{Y���{�Ƶ�/��s���e{��% B�Z׌M��݅Ȥq!��};����&�+�m���'8Q�Oq�3 jY�Ǥ��Q�x���p�ǐ.*+�q�Sg�U�y��=�ބ���ۥ�:F��0��>�O`v���]����� rl,ڍ��Կ��L\����{>i��{"����	Uv�*c<�+��:D��Q�v�I�'�cB�	+�\-?�WT���f��M�o-
u`���-��������?��5z��x��|=��Q�a�K{�3���������ￅ8
i��l�ZU�I�ox�k�I�2��R9O�ú2�# ��R�a�\w�io�o�)�*_�;�?�<����a���?>�[$�3�Q��%*9ok�7�}=�#�Ɋ�Zn��A�j�V�ȏ�`�ޒ7[��ѧ#��흂�O�ô�Taܖ��F��4��F� ��dP�E;��֕�vI2Pױ> ����&5��#���e��q�h�Y� ^C�J<l����2�����#�X�����0�����!)=�6�5�9���RF�D)�$+�ǲؾ���~Yc��찥����K(� "��DS�������c$Z��6�.n��Κ;FȳJ�rI�����Y�8�jc��O�Q@͑��
�ix�lDE��
O�]�g9�@7+8Lp�9@ɉ3�����1��% �JT��\C�4�TOe�]��xQ@��msʾA\B��s�pl�r�̸��6投�Fb�C���[	���1�	�4' �mգ.�ܥ�!(�9��q�9���% �t����)Nճ)v��&=w/�LQ�7�&�kC�����u�M<�q~��=�PBͳ�V�@��늠6��<3�a�����.���fb�`mw��@�t8�B3�]�X���~r�=�w&�k���AH`�GM��u�c���U��m�� ��oQ�ɚs��/���QY�B��.5�Mc�!���4J����Y�v�A�ü꾛s�PZ �����|��6�$#�0vH��������~ѩ>��8;:ṷ�rG�kK������h����+!� nD�N3Q�-	���*�ִh��1�����-�<1�	���T��}�PDF��N���m���!k�V��`�`���h��2B5�ʲ�y���L�D-���`��U'�u�nQ�^����(&^G��;�� �Ɩ�}�k��s.��<��J�Dە�� �n1�-X5j�箔�)���s+��/a�t�І9�9ё�BI��"!�E��n��I�3@e�b#8��%��Dd�`6�!~#�j���}�ˤ��o�Da�~il��d�<� ���y��O8c�E�Xb�E����r�O�&!�a�Z~���Y�]3��YS ��\γ�m:���@;����J���c��R*e�ɿ���R�@�C����6�
��dI��`����ma�&��P��d�Q�N���;�5*������㴀��܍]�y���̓��<�}��KIU�0s���O�Z�2�bp7F���z��6oz�G����;5�j�nzIz҇��:_��(��1�7�o�-����!�hd�k�i2���J�%��Q�B��7S���`�$���M����y#��IN�;�1Z����tѠ��`��Q���o>�mKɴ�iB���{3�c��*V�b�M�WS¤�A����tb ��m�Ӎ?k�%���=ߋ\@�f�pst��d�!hG1S�� 5�;tޛ��'h^����[�8�	54^����B��u_y���'o;Y�t�Rm�-���;cP�'#�I�Etex�w����5���N�0~�u��E���(;̐;��e�s?�*��0.���������Q�v���ʜ{��4��tU�����/������r<W�J	lx�N;����0
_��qI�Q�<�|媢���w��8�p���;t~�F�@ �K��^I�c/�l��K�K-7��\��`���S���)��/U�4�)�u���܄,��z}i���%v�Ĕ�����F�9އ�f�{:�TX@B���%B����S�]��N2�d�.i?N���Ꮼ�(�D�ٽqu����P:���6�&E��S�_4�c�A��<�q�
7�����G,z��Q.�5+�Z���5�t\�S�|boR�S�1��9�ПҒ��4nn6.�^e�F ����n��y/���bͰ�)U�b��)"�i��'O�C�ﱒ��o�m4���Bh��� @����������y� �U������h�2��Mn+%�L�H�$)R��Z�M�1^M����Ϭa���(���2vT�(�R)��d��?=h���ar�E���7�T�*�vc���q�Ç�qG.� F��)G�ۏe�z����[�<�����k��Ҹi1�>��&D�!���Ƞ
�:]ad�g�@��^�z�!���|f��|RyT'���YG\t]|f"�`Z]az$}l�D=��Չ{���a؄ܿ�1�av���0��A-ú1�Ł��^
�?�0�q�\�b�|J�k�Fe��l-9w��w:mRQ�M���x����,���ѝa�'oFԀ� e�N���[�`:QIR��ߖ����d�c�S�H	�u�<#}t� ��G���g�x	£w�e޲�����c"3�-
Uש�֕OM���A��~#������j��BX�=�J��w�[3������!�b�[j����؎��2�z;�/h����	�ED(�n��a�	������9��{5�VW�r@.����R��7]�pH�Z�tʠp,#�Oީd'�5ůPnX��Gz��I�dR���v>��$SU�WR���W�雰�!��}�Z�Ɣ:�߻g�p��XR��.h$���R�fP/I�]����a���#SN�T󤧅�}V�b����ҷ�
|����j���m��6�a��߅ ��W�T�3Ӓ�v͌��W���'ш�2l�i-�Z�=�+O#ə͊-���°"FJ�P�Ī���a����)j�C9�����W*��+���'N	�Nɭ��i�������a�X��3�lK~��R�#�ԫ,�)�մO@��WX�B��ª��ԣq�K���^$M�J���J��}i!�Tɺ3�i�u�UQ��=�����S�5\�d>�|,,s����,�ۦT�����7�,vЂ.�����aADr�,����� #��|�
sg-�G,,ģ�eϭ�%�Cq�3e���[C��*[�Hu��n�띒,%Om-���2p�D���7���K倥��on۳�P�A�\ ��Ƿ��i�^��f�W���U@-���3�yF1�Ś2�[Q���5?�y��6�c�Nt�=4�={�޾�G 'v������Yy���a��;�t��_�ʘr�����x�X���P3'�u\�v�v.��r�;TS�@IdP!ƃ|}��|<Qpfa��a�s���~�ԟ��Xң>eJl,g�ٿS�<ܹ�����Y���<� �d|M��	_�1�\��&�a(���8 ��u�T����B���$#$��<ϗ&�����q�.������ܛ@����t�� �����a�~��lbIjIb� �yqNIs�V�s#�pYN�Ʒ�r�q�.ȏo�c���6�h֏�uH����pWCC(�a���8^�4�ubT|�~D��e��7������B5K�Xٚ��$���5��B4�p�3�l���[���㖺�~�Z�T.{Q�/]y�y����f���`j��4��Gs�7+��k-����C�F|I�t7���ڜ��'���,�D�}�&[�5��TL�UқPț�rJ+�isǄ�Ǻ�ge���q�q����s%��YuN/ƌ���Q�ǳKU����%{����JK�ET���x�9%9+�[=<R�g���ϙ{ԁ�y�\]��|V��8,!�'��Hj*"�RT��oX6�fȷ�ePuʹ���f +\}G�et-m0^X2BU��n�V{�ͼ:q?�Ԉ.	��<��W��~S��3��^�5��e�U��V��"$疘2/;C(;�������w��4 ۤu8e���X���i��w{ɀ坟���Η�ڂ�teez]�K,g���{�@[Z9��i28cA1HiB�{4i��sEP�Z�����;��0�r�=Bb�2�]1WGɜ��#9��>�!�FQ�![k,����?�!�o2+�����o�>��=^M����o�;$#��,�x"n�ϳZ��.,+{qP�X���ҽ�ȲI|�"�z=�+��K�t�{<م������Ћ�{u&/���%(|��� �4a2z�vHڙ�ެÂ�q���w�r�j��cY�GO�a(�
żyBs�H+����
 �ג�3�����<#�����Q �펏��"����BҤ)�=լdU�+�H0\  >�գ��l�r��	j�#~}폮#�-����95u�є����@�'�u�BӇv�_�	A����;2p�q��S6bn�u�:u��^MHۀ�A���1K[y��&��>I͐O�(��.nGa�B���\1x�� �϶�V۫����Tվŧ�� d�JpR4���C �l�}�֙�����4ۻ��X��ZK�s�}/,B�v`�63p�N۝'�"6�	XBeL����]����IV�\�]:d�d�*q9u�{qv'�,�.�x�d�5�7�3�� ]������ i�`ă#F�������E��Ų�Oϖ!�CƐA���͜gmِ�mnxg�3�l9�����U��v�dG�ɏ*gN>�ՊC�b��p��؎}��y��C�<�q����ډn���:�����k�nVzD�O��ɵ׎�3�r[���e���S\
B$h�`$�w�Z�xk� ʢosm7H�÷62�v^Q��5Fl��Xep����E!U9^�s .-�o�j���I!���fC�����R���0X����Kh�.`��dLi��o�d�v��I��Hd�F�w���v;=ڝ�	H5��GƜ)�Q��o�pYJV��$?��2�K�8����Mef\Q5�H�_�>�55m7��z�\����n���:��p�gV�#沁B�m���^���L�Y��]�6C�������!P9t�"_�7W�n�f)|��5�{�>�H`)�z�6�,�W�)�76�ʽ.b�aCV�n��֮�	�
0�t^��m���|'\T�t��_%j��k��=��D�#7�@lײ���3z1���'fq��xM��WX%�_���6f�����X�%��1�������y!.������_7UѦ�Y�ʕ����z\.y&u�6�Ƌ��B �M閾��3u�f��G��V�g�͝���EQ�Eg@i6o�g�ŉ,��\����
tI$5���K/֌��ǻ>*�p����F�#?���i/2�x���K�H�|���}sߦ����Pĭt��A���B�9�1!�d9��m�q\�eZ8����T�ى��!=��ע�FvEsF��^`�����E�Sx��b1޺Ʒ0Uo�\qa�6�h�m'��Kɂ|II_����O<�F�͖Ktk=J�5i��$�!��¶O�����=�OjQ3�ʧ�E3�ˈ쒫�����X]��iZ�֫^f/����!�B�=z�J6�$g���;�s�@@�9d��B��UX���Q�Ty�D#�km��IN]�4��5v�GCB�z�(B������v�he<�5*��65A2��SEu�E!�^�%
��!,��G�K�"qUQ�Ͻ�KLr�:�"��r���Xi@T%4�?!�S�"�g�MFE'�o�C�+zE����|3Tq��A1]:�+G}sH�S��u��}�S++����+��,\>�"��� ���J����\��٪<�P�Y���5���?�@
29zIV_�N� �7���A<ڹ�f���EvYL��K� 2�V������<:Q�Ƿ��1$V(��I����E�Y��jV��?밹��dR�i��#���cw�H:�֭��8�ɣ�u=#im��p�_1?�+x��!�
^����f��t��uCK.��Lc�g�kyf�ym��GG�=6��u�0	�
q��NG���F� Z}��Pgx��~ t@꯹�r��SdzD��O�acV�˼��4�?t*E�S3��xz�����b�+�d2�?ϟB.�3�P�Ğ _G��Ϫ�p*	Gz�Nޣ����I�z~��z�0w�y�'<�Gf�A�zOmd;�GS�'���*���4�tgqM�+��{M�Ye�V��e�K��p�w��o>�����X��,8%�P���ym4�� �~���a��6����k��o�=Nne1pI:N�8/͞@iy��ȋ)���:�gF3'j�.gm"�TB���nF�z����/��¤B�{��
�R�D��E��6� �=�F��G��?�&K�8a�AnO�
���%�W(]�cY��z�Rn[�b���^�G�g�#�T���*�h�����Օ�&3m�����TN�X]�27��aP��:���j���=����rPX� q�n�_-�p�2Zvg*7�V)����]� MH.H�8�iU(� F)���M�H\�6��*�2��m4ܣe?U�����s"
�N��J�;����`��?Xnvl�{{7<����&��fB�z;��ҷ�]���B���F�0j{p*�2���>�d�&���`z�����UXof����Er������tץI��ܱG�����x���3����k��5�C�j\��A���-��=��;��YB�~���d`��݁�4PY���0p���z�'�i�-ruo�җ���gvTd�Zgx����*���z�0330�O+[�vC�AV�y��� k�����-۾вg�X,0�=Ż��<�Rn�j]�^V���c�$>�mC�-���px�
`������~� �Q> ������{>K:������M������c0��d�� �a"E�����^=�ZQ�}��yY3�H�.Yem��R�K�%e nv�#�1�n�T/.�P�2�#�ƛ݅�p���[�*��k�U7�}�����5+s������8�3e���=R -�hįU��ֺr�����7���َ'N'�IO�NCء��:q����觎|p��x
�.��xq�:���w��oʐ��ت�4��ABI�]AD�d������E]�kR��a��C�MU�͊Jk~�L�H�Ly�U;����ӶP���%,��,|�
r�)��q�۟z�v��V��ޭ��g̇a߂A%2h{R����`��l�c���E����F3vCn�	2��/�����lsG������J��SYsY;D���9L��n��3�1~ܢ���|��Pl�({ڛ�*&:3��d� �7S.�xj'	)ŒT�t�oV�?Y=�8����
J'Mc`��ĺZˬ��Y()��,A_ʹT�����Ć7�)H_��m�]?ޒ�G���*N���} 1��=�
݄G�z����1�Y��]b����O3�y�
.i�PE��r���b�_��ƴ�;�b��ٸ�bݾ �?"`���Fj��:������	b;P�۹�+��z�-�͔ɿ�C'���\�l`G�0IV"�7jqdo)��ϴ:V��+K������_D���D� �OJh��OXX)f{䜆�9�.�!CUQ��.��o��)���~<�U Zա�����r��7����g5G!��r�"T�d��Q@����	��q]�޽�װ�Oݕ��c�����f_�O\Γ2��ו���[��#�b-�F�-P=Zq8a�UD&��� t��͹	�y��d'E����#�ppg�dv�,SP�
�c#K�T,#��w��q��	/<���lI��o�bɇ��h����*��G�F���6B>^��e�E�^����*�����J� �_�+>�w�l���Z�\t���ʳ�m�(iL��'^�=eL�Z۹	��?�VM��G�q�:ӝo$A�~�<�߆[v|%Ɨ�\���w򶒳�.3���rr���;�����"�V����+����b�D�{�f�6	�lR.I����)����-�����̛^c]�e��5�\\��TjRsMF@,d�YDВt-�I��@g%Z
�c)X�|&�Ze#ex�����|H����~Ww%�<̷�`�__ok��$$t{Qz���У{8%�s�^�֞��3��֟!v��'t/^Ō��3��OF~� z�ν(���d>���؎��	M0�h��&��!�:]^�����I5O9�IZ3{��6��H,�o�����B�s���-��b�WY3��&��7�U6g}w��쾹F������
�)����Z��%��e�r�Kb�s�A7K}8�g��+v��[�a)�U�C1zY�狁B�����c$9M�@�6/�����+WB$�����P��$Э
Τ�����:hT�ѹ��"?��n��b|h�C��[�Ÿ�$��By�� �c=�J.��u�R(�&t�t;T�37��t�O���2�X� 臖�|p��&E/1m��y�g+�CH�1^�m3���\��x|j��*pW������O�Ӥ�z�@��슱G���_?�^�eS�t\���4
��]����;���?=�]fFH�`Dj�a�9$�!]ab�hu�j���:��x��#U�D���.��]�:4�+���������7u4/nM�p]�L]z3���YR���Aw��`++��Y�$�W��29Qr��2��Q�槺K����^v�^ ��#��a��Q����d����R�>��3�F��b�"�T:�	I�n�O�ֆ�������>�|%>́�B�f��}.K��a�磻�u�7�Q�Դ�Q\��e��.��Ѓ�+�o�_���
%����w�1M�Oe�}�[�Q򱧁�폹�yN .�n���h���?#��_���S�w��	�b��v������h{-�jK��n��Z3�h0V�{g	[�ej��@pK����ډq$:gBt�Z�c��r&�qj�+����u8���O��)~�ү,�ͣP����j������w��J�`3�v�|
����A���'q�`���l��C[���qpĩL=���'�j�qZ����q_n"����ܞIG�J��&�a*qO�p��\F'Lmw0�9�Ϣ�;J�Na�tI1C��s�J��J�Ԙ��]�$�/BW��*��,	J��Yӷ�}׉5�\�����;O*c�:(m�F��G[�ZV�DgM��΅f|�}��b�g;5����5�]=F���:>�"64Z8|��A~���q�S�#��O�i:�V�}�t��}փ�W�_j�?;��l�̗5Tʥ�:va}�6�g�bya[c��\����g��V��H�w�ߖ���c�J_N�\\�6�'�?
�ty��)d���P1)�g`1�>ܵ �)uG\��W����r�@����[I��ԏ��o)�ف�88W���G�w����B���msdL��\&�,*�Q��<e�c��O�MX�:�gn[��Q���4��1�-���=N�L�U��Ғ��$Ӿ��r�D�c���s��}�#ͪ��k��} X�'�r��P���4gf]A4[�<R%.� ����i���
�.�c�$,��4��pN�Q0��OݐV���Z4!��S���-b'�ߔ���;�����&��y��yl�-s��q�)��#�7������0�p���	�uf���keQ��?U���k]�m�����˕���5���i+½Gh��[�IB�Z�����j��IO�[����
>ދ�4d�Ɍ�Qr�D�[�@�P��������(�N~�C�<+����IgW����ly?��))G���H��qy�g|H�&���
��n�q5�I��2�=�����uQ�c�J@��/	7��Z^���6�c?��i/��q��=-����-}�oC���䵠�2F�~M&`��� n���HF(f�����1|x��p׷G�� �.:/�)�2�|�'j�DzN96�ޒ�&e�r�
W��ܦ�
����3��1�%4�����\&��Q�Q`dsJ@ó�7<�^"�8a�G�T����S��~�y�����ћ�}*bb��YN�|~v3t��1���M奒��e����l1ܺ��:���s����a&/eɾ�f�5�ye&�(�ޅ�x���uFZ��9�6�! ����e'�̋�C��f��@����X޹���L��F��	��GY������o�ҡn���̴�w��=�b��rq`�����Tz�q�b��>�H�T��ʴ���ƕ(n+=��^Y�9����6tY.KlwR��[�]�V1S!��Pppe�UJ~�j�'D���=�ḉ�z��,df�q�����H�e��e[𰂄�rV�Y-!�Y2��h�F�X�
�e��R6D��#`�=_ښ�)u#�eX^�~�]�c�่�+���M�M�=R��@+���.՛���N��w(���S��ȫa��3�'R�m2'f~@W�)� ;c$�j�$?��{��ݪ��0ݵ�ǆ+��ߠ".%{`~y]�H�������T�k-�c�.p7�J�O5c�4�	5y8�Zc;ne�����7"&U"t	5� �� s��Y�R_��T�whp�D#K3� �2p5c�u8	�]���//D<�DAQ�^ܻQ.�QhU�+����M��~��l�#e?�"�����?�_����|�y���QZݓ7}���ۮ�wPH��*�& �~u����b�]a�D ���3����|:�OөAq��2{? g[�����܄�&���1К(�{e�>h��N��9�$�ќZ=}y���34�,x��n��)��'�>�P9�'Ń����
I��_O@��t���Fi�	�D&�h�:�&:|
*��N����J��h=J�C�1�R���i��4�̜c�k�#HhV�{�rD���MS�I&���M��L������髟<�|{XPD�i�G� �}�{C>��>�t?����%�
֟����g�kO�H���!R2�V(�CԲ5@/q|��@�2�$�z_��Kd���䥭������ti���n��iS�}�E=&]�O�7�������جF�ᲀ��~��c�5�[)�m�����]!��cb^_�OX��"�١&�%lt=�mꋣ��2,��9��ZJ٧����j�=ի��!�!�2��v%��P�サ�d'���l�MHk����/(u����J���Ǖ�K灬�#g��B�A�������]�$��أ���SHJ%������W:���)S����@M������:���Ǐ�:=/s��'i�r��mO����8t�Ef�J�fJSd7�bJ�G-{��] ���m)��K���	��*��U�	�jc�����C	�=�J��p��W��6Mf����f9�>ܻ��(�3jNd���oM�~%���œ�({5wR.�S��E�R�ǯ��C���Rr�x�8?o������_�{�f�����[��V3f��H��w�J8���e���K
������AZ�#�����U��#�V�.H�c�I7�̛oF�� ��E,� ����%��ZM6�~�!ǒ��Wxw�uOJ�Td��l5ϼ���a�և�C��ٍ&h��>AWzQ]��B��IRH\�-�ڧ[?�f��j)�\�,0��	ܿ�Fy�L���.r�?�Ɲ�������F�J
y�
}Z�u楈��͉.�.��>�Ը�3o�������Em ����c��L�w=䒰#��@Q����Xe��K`������O�h���ߏ"�����S|�Je>�⃚�3�ݜV��Et��*�I��71[^`X�F���?*�E\��ֽ�]N�( �Wf�KW�J�+]p�Z�f<q�F�*M�p��L���W�$�/�Q�y�u]�6�K������v�ݟ����!R=�5���<r��0��4P,z
�͎&]�́L+T���i�i:�|�����&XQ�X��Hz���	�/�/�#1I�x�l�z
 �h�ps5��!��c��c�F����Nx��Cu�E��Id[��^��s���̃ h��<���� ��ؐ��aP<�Tc�Gl(2t��Z�,"��
Q�Ҏ��Ѕy�b�y9:��y�<uU�*$"�>>Y��NiAί:Q��T���-V2�_W�
��;Q��b8�uɒmM���Se��c��?�-������_��3��NL	�C݁!b�<����˘�.a��^��/�<7�W@���������-C�J��y�NEwnoo8#C���.ޙ�[t(tR�3�2����b�Ռ|
�`.ct8��M6�b�X��W=d�L�#�K۬q�AZ�{5�C�	�6�6-��ѡ��
��Y�|�=����>�F��o������9v�y��t�xR�k�W�̩��
�9j)!]�7����p!� g(�����bdʚ�[ܪ&be����m�!�*��i����~��E��͑�gY�{*|�
�e�0?�0�]�,)q��T�����/R�bҎ�8���2DG�2�u�io�����O�m;Q���i_�G�8��%�-,H6���5���rN'�+=�Е#�k�$B�p�}����`����]���9������\YHC������,yD��1�YPn� ��⣺^+�é�}�A.�
C�Egh(9Fۦd"1W,����y��F�vw����/^5���!/�����B�E�=$�� x_� 5x����XSn�~u;�^2�1>�Sx�&�
�J�d�����3��b�sV����lz>D�@�[Ud����p���@C�+���YfF����'W�u鴺���P[p�	Q�+���D�E�׬��Qcϙ.����?���wc���hEh������vI�x1=I4�oV�K�Ǒ�x�#�fpg��L��嚈#��	^p?*}Ts&U�@�'Jnw߫,=�0LV����5t�Z�'u�TpR�	d�KZ����o�:ͳ��);�'|yv&����}�����fq����d���k^"K�Qo�	� 4J�������4hUEF/�������O���C�.8}�j�x�Vi�:ʚ��o�Gpu�:
�Jh3�۽{3˭-H�YFy�:�"ho��^-E�x܀�h��o�l�E'��� �6ud�����* �|D�F�
��A������)>C�~j`{�4��d{��8�B�@L�SjD��i�~Ϲ�`��SG��rM�=I`�Z�o1��s+<#����q¬��ն#Y��,U)@�<�YJE�xv3"_ UW`q�����'�a+(Q�:�IU]t�<�����τu&� �Hf�(��[�?��Je���Qe7�4�5X�@~�+չC�<���O�[�븬Y�ZS;Z���$�9�>R�HR��E~��J�=��^��Ԡ!pm:���VY�#\[�{���2�2��f�E�)�g#Q�^v�c�p<G�}�B�r�WNg�4£�)�D�;�����J����@��	��5cw���_�!��<�{�N���s�+g�M'�\����x�,�Xț뽠�A�#c�Bl��vY���&�d�򙫨U�C"�U�p>��r���\�p�[0��p�1�p��-6�%���D؏��1�2{6�9�j(����3E���ధDG;���ț�2ȉ_n��Н�9�u/��R�-~x�U�
���J�u-u"q8ٿ���h��,yj��z`o
���/@�`r�D�zd.J�Ӳ<:W������1m"H?�Ɖ���6*
�m����M.0J^4�H���	�b�h#bI���?T�<��%�؂c���G���XLl5F��|��)�u�e��֐���6<��Ͽ^tnw���Dvm�P������1����fkp���~(w��3n�������$�.�HVU���,��Foݓ���Hl���@]���y\d�����֘a�s/;��a�)^��Q)��q���g�J?��Ȓ$�����_B�/SM*��+_����iť;��To30��4����s������4��&�9sL�Ÿ|Y��2�p�H���q=���
�H�K�㚍�\P�:���zsɲ�x��`��ʺ��Õ<��b���_��LF���C󤇈�x����FI�&�u���ǥ�0������U�Ċ����=�?�����!�̒����s��׬o������M�Tg�ac Y�IgU�b��Y�LT��CF��=7�0��t��Z(��ī^yVF��]�)��k�;�p����VT��CF8�P&�V�D��/@��:�Ut3hRW˸��]�|8��r�[�L͢�e�J�<EFB�Q	���>�\�����p��Aw�����+mTi/"8q�Q1t�R!J����z#�:q�-8�Nj��1L����N��հ�sS���@'Xx�X��+�#e�Jn[�E{<1���	���9�� C9��]��-� :aSPV�̈�+V7�϶��D��wA�G�:3�0��L	��r|A�)�>�r{�^C��mL��̟�X��s�n���CЊ�{�y��\S�-_ZX%p��-,�uD����-�
����`�ńN1O̝�^l��
���cE��T��v�7�@�4��TGl���_��,�:edw?�ʨ��D�=ڃ�P����Zxt��\��5P���rWeנ.â"��D�C����I��Ob���S�Mh������5��|�j�?�O�N>�Oe#�z�ㅣ/�/���0:���s������/H���Vf�$��fۯ j�rIOg�t˸�ί���t������q��Q����F-�N���. +y�����@��.����ZĀ)C�9�96A�3�j|�O-F�e���{��W��	���A�3g)�M_5Y���}��+'���]�ƴ	^|u&֬ف�E|Ɣ�]p>�C�[M���pӥE�GU4�$U�����ȅy&@�kT�I�ۡ��!����A��X�����5Rͫ{TE|v�=_�gVD�m.�����QOY[�4"|	ȏ���j��r{��|�YfM�1�+�l���&�i���j�L.�u�7�+ ��,.2?rEe�ALV��d��I[��<���aP��T�G'�B>7h��*��!�2)��HYտ�������jOvyd�n�8�2:��U�n�����P�*Ů��l���"9���s�y�l2i{R�d�@a��x�`���T ��Ui"��r�ȭ�H��VR����b�^�t�	�*�N���U���pۂ�(3N2�����ϓ}m������g2ot���?0�K�2�������O}��� ��uZW��4o.X>e�M���4xV����D���i2��������xS�5���`�	��Ii?
a|]�3R��\�*�p�l���U�GGǱs��kھ��:�;m��5B��.���\0�bA0�����8޿��D���]�4��fꢽ�E�>	��6�����FhT�6���q��u�wz�ۅ���t�~����sK`A���`f^�M�p��m���x�y�2�1�H�s;�����42�je�������#���6�ocD�_Y�EZue8�'	�u&�����#}�h7�\�^V��k��/��V�%�~���[�P����(2���UPw�l�Z�"��JB@x��ˏBN�ū����8����>��"��x ������.�}�tK�p�/���ؕ�\Y��0��K���kD���ਚ܅����t�Sd��������{�|=�J���~T�n�[���w�L~��������q��E��1`q�0}�Rʍ����T��`6��Oz'5���pP����[M? �p K�7�N�w��I�K��!32�gU��}�S5��*m���B�p��7���{uo���yH6�g�e�����шѐ���!̟�rU���tX錃;��v���d�Fk�8,=�|�ƌeЇ.էյ[����D[�n�DP�R0��-�f��_�|!'�u�J�=��_�D��ܨ�[<l���o�r�6�ݾ\L�珍P�<�fKէ"����ʝ3���
��% ro˱m�;Ϝ�/���Ph�[��v��N�(9��w�^oX���۔_/����%Ȇa5!�R#��zx����D$��v8IBhs�X����u���&�B�fH��2����K]^�߅�2�1[iV�6������I��s#�֣jZͪ�:�{���^^�
�ٸ��:�F����3C��C�F��A �;ۻ��~��ɜk�9�"գ�psl��?��e313%��iV�Յ���o����u�"���`g�N�A3�����R��|?���a���e<c�^ط��s+vp����u�g�5��IƩ	K`�M]O���p�����]q�f3Q_M$�v��eg�őJwi2�@���O���-QY�^Ĉ�m���.t�]Ihe�Fx]�Ӥoy�O��X(����o���/qԛ�R���_6CŅ���@[}�EL>����Uߛ��&\!iv�8M9����یB����E���+��W��ƞ�Cġi�������qrh�&`�ʝ)y�0lf��Q�	/�/�� �g�d[v�N��Y��*�A˔���
^?hej���(��ͥ���<?�_e�6M���Q���#�X?0F�s��tJ���.�6�$Ǧm���F�=�6��7P����$�Q���-1�K��q-=H�E��#Un</�)�`d<���ޜ����x v���[�g��zʽJa�^�xO���6E�}H*���o�$jӝ���+sj�PG��9,S�/ޏݡ˼���D0�|��������:�b<�P����Wh�2rc@��@FПi���� %�,:㲎6�F�Le��H�
�v������%j�~��PM� ��c}-븊�AG��V$&�#�0��Q6��xN�Fb�0P��c�3�
Z�fjyܞ4D��*��5���y:��������([z�8�~ ?Nj��|���wb�u��[Wh<Z�0s:���
�dZh˾(�BH�fɿ7��;�%?����� U"|�L}^>�$�+j8g,�h��s%.ͬ�ɼ��Q�@z��&+-g~��	P�$��=���6Q�h�����Tͯ�nt��x�!(=#�%㉑�u�۔���;�n�f��_k��OJb>�|
��W�����&����q�]}��|�3���X�p��0ðdc5�Qsϫ��%&=0$�la��z�����y^;�'*�t&�b8�C\�I��M��t�q��K/�<��v;��7��F���ö[И�e5z�eRY,<�ľ�+Qz�{I4/I���h��.|�oi���Am)��.U���O_�pd���[�H+sf�#��7�`��G�~Pc�B6i��G�D����z��&)�Y9K����/��,�hI��~�/���qjVgê-�vŞ���c\����I�,h��P�x$��%���BD}����J�*�ѵ�o����T�����#?Q{�g�]v!g�@�����xO�o��;�I���3Gy�촏�k�,�M�̧��WT���޴�q�rM�C8۞&�RR>˴��(���jŻ�\�Ji�1�y�Ry�� ڈG�Wwk'l���J��`'�s��q��5(̗�Ԛ��y�b�����?;�����<n��ǟ�O��0��_���I�rj���0�罭�p�8V;�ׇ�P@8�J�P�Ot�,�\K���f0�Ϡ�|Ɯ���{p�Ot"��9]dJ��K���n_$<I�O����Ez���G.M:��d"��S.���G�cf �P��Ϧ�r�X	^�g�������u���LM���륪�x��l���Ɠ=q������f���%�[���朗�]�=���>y*���!�� δߪ����=`#o�NǼ���6��p�+Y��5�7{�^e����||"�{�Ć| �JwNpţXb��x�@� �*��wK�-cw�`[���5d��p��F�I��ͤ���o$"�	u��sI�D
�E��it�,f�TA�rY������r^0 �GG^n:�~f�Ǒ��1��Z����x�c�~���t�Kԯ�W�0D���`�AL���Ұ�Ӎs�WDr�Qn��Iu1����r:j��l��	��*	�As�8�v�RSkd��.>��C�P�̲��륌�t牒'ڢJF��2u�p�k��QUD����#�MsԂ+��!���WFÄB��M@j�P
�}�O1�����t^mA�z�Q��Q[�Z�.�r���oj��'-�b�Vu(����Y������z��P�%-�ds�'/j����u�!X.��K9y�q|#��a4����{��`���g ;����wC���1x����E8#L쟨��� d�s��N
��j��
��G�{���*�;��69�'���!>��T�Ċ�Re'A�P{"N����<,�쭡!Ɂu�Cx{7;��jBA��M�eV��)������#3A��!vz)$�G'$E�{�=^�L�l�'S����w�ʫ�oW�����p�4�b�=�$�w�O�s¹j�����S&���!μDl}AP�9<G�q�b}�L�]*�'���U0��_̔H�d�׆g���N�;�s���Ԟ��Č�o�K�o˒��k������R�&��dq�G�G�]��jW?����:���zq��|Ƭ+��$r����$�`�|�K��>߾G�tDa:z��j$oY)�3�[gRufny�kr5
�	v�����T�hRW1��f���9�Qj�v?Ij���gY�M�	�t0��{U�F�V�� X����2̈A�/z-�T�����~*�I���'ʼ�;��&��ä@똷�n5��fS����_֖�R� �V9�Cҡo=>�M4 B`��0����M���c��,?0ӘrC���pQZVn� �b'�(r�a���8��Q��s���n�����O���R������@�*�}�A�	��}Npٱ�h�eV�79L��S ���W��N�a8�;�5*C®˖(Lߡп��i*omdPiPD߿�-��W��l��7Y��#�
��/���0�_ <[�{1�B�
,�[���&����h�"M��3��/8�#5}��_�GC�<��!��PY�!�#{	�n�Ʀ)_>���bW�K���cMaW$�̡ds�$���\�ŒA4���5i�)�������{r�|�O"���|5��Ela�M��:����
���Ea�!I ��}��ݖ�p�#�R<ɸb3��o~�/Z���,�ČV٭ܔk�L��ܜ����(̤�Ǽ]��/�#Ƥ@��ϓ�@�^Z��o[t�W��^:���2Y�b�$5u/��W/T�|:'^�|'�,�ܧ�b���<<�x��~�I�A�'�7�a�i%��z�q<iU?�S�=<���w�6����ac�[}����WZ����/��%�h9
��k�#�*��
P��ߣ�.�)��Eٗ<�p���/.@��aRhҠY-����<z���6�jb��ի5�4�_,�/�a���ݕ\����"mQϖz{� ���h��\��#���j�Q,���b�G�Ab'��c��}?��,�[L_�x��E��AӨT��Y
�B��*��;�n�mȹhYv�n�q�������#	� Q88������H"C�o�j�0���b tq�Rܑ{X>Af'�?����-iݿW��Y�6�{_&���2l�C�{K�3rKz�����T�z�0�7��'�I�1� \���*ՏV�b3�cMԴ|�����T�}K������j�LW�oI��\��O�˟����rM�4jN�`�;e�ќ~�P�`�+���ԿTly�Q�W�&��gʇ�"��.�])���3�Q̂�D��W~�Uh�l�t�g]��]��d�(�ͺ,"��V��˰x�m�k�t�c3:�j)�
+��G�y?"�"��Ү	<�����SBյt��d<PS`MB(R~4 S���o
���Z�O�QD�O���!�	"���/�B�����C�� ��O'SQlx��%�6�0���S�xզ�yL �е��ro��o���� ��X���E7��s�������K#:����ԵP�X�mX���Q7�g&���e-UVZ$�ь�.��.g���q��'�������p��)�0�~�ڐ_���̓�l�HD��L}����o�����4�0_��T�_����/C}����z|����X��B#���\wD4�u�P�1���5l���Z�˚f��v��j��5�����	N0&H�D �#% T
ꫧFX����Q�B��V���<���0$I���).�ϰ��!��w/�R?g�7,�GL���.s&�S�]1'���u����%D��ي����w�n%8y�uC�=Z򞢤���`n���]�7ν�/���l02˿�Y1��㴣���n��d�OЩ�R*����g
�G ���ˋL�+ܣ���������Ii�H��`���������t�)ň+�Ewg�n�ӣs҂+�S��8�8������ W�:hwͪ�h�:Y72��FL0tY���𻓾�Nz��BT!��Ǔе�HM:�5y��p����D{��%ප��I0�3�Y>C43��姃��h��f�g ��>��
������W`�qR8������Z�A��xa%jC׬�}�S�*��u�6؆���膥j�+�T�ϔ��4^ /�j!�A�4�����7LSHJA�-Qg-j0������E"B@lX���8�=���_L�E�7B��.0)���G*�L|����׶pI����7mT���ez�Z�i�\ZV=#iI7��c�t�w.pW��4�s��M1]e
9)6��&M��z����S7�AG;�O	J2m�M�U��k�d�q�VNZ��%^e��F�d�w�ε�a�B�\���iV�k�<���a�7T����D[��h�y�#^��Ł������G�ل��S�������W���C�#��m��Fg��Ԭ7��S�K֧��>����h��hӖ��U�I8!\�_�s^��NѲ�y�+ے+�BĖ��C����ͨ��H_�/��I$ i�4���B����c)�?M��t����ph<���H����	�=t�g}��oLd]?���~��H)�b+l�)}��A&/���t1��Z��J|���\��.�w~���d�H��_V��N�T8:�U�(r�%a�A�nK��Hl-{�~�����Q�f����8��n��n�Fh�H��B�F5J����
�Qo�6Ӥ:�Ɛˈ/y�S�.����ɝA.N:����>�P�k���D�P�����XkUϚܔ�44�d&��/<}����3���ڭ�����2��E��sH������-p���ZKS�����s�c��8���]-E�b�7�Uķ�۹y�6#`e��͐-8Mc
��A��݅��y���L>�҆�cܤy��7��7��T*�9��B�D�da�uD�ĥ�揱�`���Z����ҋ�V��J���$w/�b0��0a��1�Tj�
��.^'�!�'�>��U�Ց�M|�L��P�)�O����nMQ�l\0��6��i�#b�4Eb.�I9<�R�ī����I��tx�=Q-y�a��wе gp��R�'z���2l.Y��	E��Y��6�}�~����6�Zk+�ua~
� ����;�Гx�
������4]���i�D�y����x������P�$o���p�s�r�Ҧ�@�w�^��/ �����lڿ[f�cڞ8��gm�=�K�-i��� �N�[�Y�^���l���u��y�}M��_�˺j�σ�9��Vp�%�J 7���@���i��R�{�f�"��^@��l�O�#�<}���{�N23������� ǩm0���)��kG��i�`��d>�����"�)����M����X)w���.�<\F��_��n�Kɶ���Q{�0m~�z��h�J4�=����5���/��vE�K�=�"ʌ�/����hY����SP�����	����hS�6y���$c'�И����/[e@��'��E�<�,�i�!�\Q�m � S�&KA����o�����Ґ�\�ӕ�Lu���3/��
�y�b)^�����HC��9�7���R��c��s_���"a{���C]�^;��*̀���b�xR�W���h�֕�.+
�v,�%^uE�{^� 5�J/��>�B	Ƴ��?�5�x�Ún^�}�PIh��O[wӥao�T�.�A�S;��擞O������%�6:�>�kS��,�����&�K2�?���8Cc����}ٟ�M��G�����%6E���Pg�G�F�Q�$t�~�u� (�6���Qk���6c�"Ru�석3Nig�L�=���,�'�D��Y�y�ʃ�na�D]�+����ۥ����!ʑ�3����#��f���S����Sy.�������+���K*� oR����;��8���05��	A"}8.���WfE}�QJ9ǎt�5���Ji�_�~����P�;ݖ/I,����)��b^�s���v8�3К�hje�;K[��nU«)�|������DRq���o�R�DTr���n�ʸ�h�V_PY��M�����'IM��F��n�bꦠ��i�6F,%��ۈ�&6e^ �"sD�y�cї迣��j���YZd��n�L�A��h�+�M�&�U�H�g����2����;�Ќf))�py�'s�a	�VX:��X�W9W��z0%W�'� nW�iL�x���q�r�J����Ƨ��Z�A,�M��@#���F7u��~pUP� ��R��g��P4�H�TE��X�{�~r�S9��ڨ��� ���u�{:���R$������/~�)��d:Ļ�vi�m�X���|����1�Ң���~�?,�ۨb�J��?^Eڸ��O���!Ѩ,�z$�;h�@@��d`�&P�c>�9�b;$oP�Xɦ�i�K���Ḓ��1*��$�>��A�̈j$b��9i�w�C���ft`���f�h5yb㎐�9�@��Cߕ�ʲ�YG��AB��:W-�|�1*����.��E��W��K=�SxBo���%)L�r.�u�)
x:-�����b����Ӱhrz�l}���F}�)�Tp^u��
A�`*��Z�Uy@&�_$h�����]���K\CpJM�Q�t��H�Ô��<iGȶ×��#z�dd�:o���u���.��X(i#\���� �$4-df��$����l��T�@��P��	8k\v';TA�С�+#G���Ax����.��e��	lUk^ #6c�K(i�r����ku�ؕ��O��q�Y\P�,��3 ��޸!uń���.9��;��B[����UHEW!0�i�<C��N J��<ф�)�o�%���~�L=UG�T?Sl��d� ���
8J�V�Z��3�$i�P�ꪡ��R���n2�b� ��\t�G0.뵛�$wwa�~Նy��|f�8�.�H��5s}�`�DsѺ�o�-`���C�t�<ߴ�+�`!ި罋AC�^%ܫ�/��l���.��pv��|=O�:2S�剈W�����.�p�OlUz�@8ݞ���k{ZҲ:}���m0��>�����s�R��9�`��~Gq�K��x��..i�zރ�ii#{T4e��|D����{��B]Jn�F��ωmo{�ƴ�O����a�� �ͬ�?�M�fd�ĩk9JCT^��'��a��^��
37h��)�Ā̮_�"�t�|>�iE�=PDN.o]���6�d��ҟ��&�͏�˭�P���^��W���|�DyvU-z*��޿�'��S��aJ."��(s?�
�\�g�5s�[S܄�ZK���㸇�=��2H�"9MZ��X���C�mRS����!�����h�5<^��oy(d�.G���Z«{����{�\y��^;oz�7\}i�`y�y;Yu6U�Zk��>������*�$�~��r�J��{�n%�c�ݣ�~������c`�r��)���瘖�~��:���[�ō�T�{�5��d���]��B��Dp}���,߮�OGJ
����w�I��0ڴ�T�'��+]��-�XV�|h�.��0�TEe<Ʃ�<MM��jY���B�� �f�eAEGʾ���co���
�
Y�#=���^G�q������n�m��6br;�P#�pɉy�&T��;V�|���hk��VM��7�V�w��I���K�ڨ�b��u�rX���6fp3�ٸ
g龁�3�'���uf=����O�����G���:E��*���L�Lv�	[9�7�6G�I+�?�/�X�a|1���I��f��dI�%g��{g�>Ƿ�a���"��i{D�\���K*�X���mt��å����UѣJ��ʘJ�"��m��\g:� �������ԣ���"�"���)G�v9�
փ��[���U�&z��?PM5���C�SF���:l����R}��[�}�C9�3r��A�\ZD�
&dr��e�]��8A��8��
(�����ka���R��H���[��X�1O����ި�GkU:��fr�#��#{#����@)p�kۨr�����������D����LdQKS��`�92lr���'�[/�"�Y�_��(���x�2�X)+�	�Цb�x�+�(;+���W#���^L��gX��W�r�	3��Oh�*�T�b"���3Dk�ty
��IW���ڠoCFۇ[�T;0�װ3�K|_��g='��}�;�^<L$.���Ba��f�1/*ɛ8uYźt?Zy?C�.gq������:L-<�F@��G�V�gґ�j�17��ȝ��n�T�ډ�O��ƃ�1�8� )�/#�x�d4�9��J�V'w+MqB�lٞ!���!�z�G�|p�;|���½�6�	B���Fa}Y[<C˥�H������]k!���ҚMhȱ�Z����H�ݶ��K�ۥ�{:�c��u`�ⴠ;�g�A�u �?v�>n�{¨��3��L.�8͹|I9�6j�@>��=T"�j��dm�T��e�ff���q�|��H'������>�A|�4F�)B���UO���c@TF���o�6\����\��AD�CbtG}�!����_���|kJ�޲�����ȣ�X�cd��?�P߱b��&�Џ1~�E]J��w�pO�F*�����W=�'NGz 9[y��G���I(j���N��)�C����Ƞ����k,O����|gU��پJ=	L���K�[.@�Z���mG��(`�]�q{�s�i��+����̷Gs�&�?��C^
؀^������-*���jW�z��F�[�f:?��{Āݿ��$���Y�aL�}w��8�4g����ʅk�^ןa���WCᦴ�pʈ��PW�?�qe��ˈ�
%�*Ƿ��"0{E۲�v�f�� -�O��0�P�LHr�E��6��n�`7m}�|.HERVW���Lq�܈����j�Y�d@X���ځ�ĭɭ;6+K�4�$X�Q6E�%�SŒ�T��`W��+X]KW��@#c2��(~�TN�"F� ��8xE�P���RA5�e̸�.���ᡯFKw�7Uj��B���UZ�(�Ƿ���ۯ�>�6�z� �������B�� MH���~>���ݳf���O�7GrV�Q��O ]W�tz�Ft� �cs�+�BI��`;)������:�&r�܋P-ОoyE� �OB�Ok$��``h�]xv~��x8�[X�'�)v�G�.�S�� ����D�9tx+&qu@s�)� ��JƢ���d-�X���:�e�͗2_|#��ǔ<�3�c֏HX��:���Wgr��Q��s���Ł��^6<O�
�ow���D����A��괊E�D� k[��(Io�KT�]���'�t$�%�F�œ�x�!$�mt6� O��h���v�F���o��a2�|��)z#ĝNt�:��BD��}��i<�ͅ� �A�g�o�仠9+k#zy7<���~}�s|b��	w�s\O?���'�p@M���q�W�g�E�ɞ�b��%hɶ=�7�
w��]Fkv�X&�?�8iT%����|�?f�{�Mv3J�}z�|�@�ѳ�\M�+�ٵK��3��9{�����^[{��.��Mb�.C�Eo����\J�.��[�ss��y�n�p*�e��������L����2;��+�Y�r��w��:t�8�0�[�������<u1�&a�B� �f����IB���ĶE���LU�S�?�N�)�o#,��3�ڀӦVXw���k�_~�У,���&JTF�g�O�H�/��('�M�]X�Y���k�o�ڛv�h`�[���ˈ:�h�x)LiD��{����{�xb���������Ć�A���8X�l���Ċ�W>��e�-!r�l���״4�t��� T%�n�GVJɎlȰ�4��	t����*+����(C�ϕ����ў�d������I����_�s�
�jH�@�C��@�kM�P��a�ф8ta@0�a��7���GN\�g�^���^��� _VJ�cR6����q�)R~���	"
�ne�		me�s�0��O)�3B�[=X���<���@2ߢ�A~�����`	���1R�U���O".�6���-�kyOqИ֫F�v۝���,��@����`�'��gn�0"�����-)dRf�g� (,�Ғ4+�ѭf�l\[Kl$��Aυm���@=L�ra��O�LLF�UT��E�|7�����ܖ}ƴߍG�s�r�����a� рh]�y,I��~([�:��o"�e�6���&ï��x��?Йp�
����j;d��	��e߾	Ci����U�*Ya���_@>� Ƴ��Z&��7��ߖ�0���Q� ��	p5����B��g���j��C��J}�!ȉ���)�A��b������|c��M��}����H�,'M���5��|�.S��n^O?��~�pyV0�=����Ʈ�}��G��"�������og�P�\�Kb63tz�msu��B.�V�Z��C8�<���V$�Y�m�o��T��L�;2��<�<���z���.�9X�������͕!N��9�/��P�j`�8��*�oЀ='�u*��ǡos`d��i+뭆�U�!�����Gn��@�<�?dgZ�o�UBGJO�U�+���-�c ��@�G=���牾�<��������ti'Ō1�����C~/��Y��Ǖ�A�1�2@Tn���|/@����Qi��y��9����<���_��~����kf:F�k��9�dy���uj&�fUkW
Z�$�gh�X@q[�-B𱈳��0�����C1[dC��9���ա����s�85g�;��N�d���7�Q?<�/��M>2�.:l��=�gxЉ�
��0|�>$� �{�ˣ��m9��c��ΐ����ol����ͳahO|���e�skL^��������,_�f�5�^K�����[1r�`';��5���E�H�(M�U�U��w�M	���
��6'��Գ[<_o;� W����B)��j&�rZ[k�'�<���U���w�ۉI�5��p��p ۟$%8�r�v���CX��x~�g)�5�d���ǡ<��	�����>KݨW6�ޞ�hi�B9�p,C�d������p���+l�:.��Nx8FV��DZ-��e���Õ������)G`@��M՝��)�gq�״�C"&S��S����%z9�mr>G��sT���.�/(gD�e4�)��w����i_�d�L�z�Q{��9"O�RtF���7�K']��k��}Cv%
��0�iZ0��+��x駭m� ,���}�+$Ua��)G؍��;a�X�"m��5�R#�̄�S`�6J���g0���=�_��}O�S���{�=��X�s��Z'��<9%��?i��{C�_��v1~�&]�\�^%\�2ޭ���_��+N�XG�"�+it��k}�m�v�i�D�9w��UY(߀.�y�JOc2�}�&ca�3O%�N�OaՔ%�Y��҈e�����f��K��QK뼵 r�-���l4-�8L6P!}D<���w� ���L��9��q�݁I� �ZAW�B9�O����J�G��E	�2��۶�K"�#Uo��7ʮR�4`.>�O'�&3D��ZD�+�6��o��� ڧ�ؘ��~cy�a�
OT'c���:$���J��i{�����z��M8C�Q�
�������d�z�"Gj�B;B��Y�0e�Γ�j�۠2�J%z�3���a�-�=���o��:Eatˈ��[����3C��'�L��m2c�PW��{��U
)S��$�ԍ^
 z{�BU��=0�xCO��Ub'KL�fe�=�݆dX��(Ŋ�uP�z�li?D<���1;�|���[FO�c�� ��q[���t6�`&b��t�#I�.�O�[�i������Eg�B��*7�/��
	ؗ<�ǽ02��GN C�ww�*�ID�S1=�w�F�035Vm��ǻ�ݦ��+2tj���-�r��Ǻ}�Sct]�l�V��o�[h�\�/ �w��c�ؔ�˄yf(']�>m"2B�Z�r8�������ޓ\ɓ�*��|���%��!�V{�;�lq۷�����_�eh�OJVJ�JtY���s���L�R,ؑW��]+� �0��f�K��5���`����$��ۊ)4�!ꈣ�ٯ3��'���+�2�uTN���|V�R������ٹZ�/�ݶQ���T&k�0DYK ���opO�v���[��b��?��XCё��飑{�C�&��g��`4���E��/��	Ȅ�Xޚ�����h?��m�بv��SB��Q#˄uf�����"��w��y�����-7�FN���PJ��������H����w���x7��I�c}��"kg�3`E,;��X���i��-�ʵu?����q����C�����Zw�/乯���.�fiP)D*k1S�����朥Cֈ���p�>�։��\4��j��=���jT�o�SŒpX��3�5^�,��0��Z��I�4Ïc�"/������17Y�]���3k�v�nuǫ�~�ҔK�V爣.60��\S�f�<��sd��>�F*_���x@ߤ�B����Ŀ$Ʀ�����Y�]���Ϯd}�s��-���g�Sʮ�;ސy�E	�e{V�&L�c%�MJ,��W�0��Ic�_���&'t�ڲNz����J�]W�g1�ӭf��`�"��~����.��O��I�]��P�ocE�-Y���$��}Ttc�Ѹ:S�8<�]���e���QL(��@�y_�ɧ��W�fǥ��I7����
v΢Yy�j,�?�`�X
N�T�y�7�́:�$g6�` ���鸟=�v,�E+�՚9z�q�)t+O&x~YѸ���v�\����J�����վY��o"����?�ы��U��&��D"U*�2^"TZH��{����_��!�3C5[�J"��C,لj�ޭ	?ŖEڨ6��g(|�Ή�r]�Ƹ���u��k�W\�����(��D4PX��������?��+��}4Wʔe���da�)��=N<��Z�A����j��)��B���M���L�k}_'3	C���u*p5��Þ��a@��~��QL4��}���S��&䮐Dx~g}�OC�&�i����5U�]�����@��6/��E2�R������_��|A�&��G�e�3;B/�D	�9GooRj�����w*a<����K>����t�0�zZ-�&�_�D����	�H��Z�Y�s��Pm{0�;ǅ�#�%<�+�*ޫ\)P˺��ZN��p8kp���g�8F���:��S�\�Iƫ��\�5�3���w�o�q��`#ژ%Z��|g�( �{L�VT��3i^��|z ]�d�@���K����/ F7j
�U��n�=	&E�Rd�|��"Ĥg聑u�)J?h��+��K��.zHy������=�c?K�w��;Ә����NK�dV�1���`i��-��D$�R�[+|Czyg`x>�7�E��,�#O4�Gc.�MM���`��ټ߾��w�;*�!�0����u�U8Ζ�����w���x{��=��R�h|�Q[j �\�pګP��d'n�Yva\�j�&>S�
Y��SLj���0j�P��m3�ʈ�����S�hM�
2Ua=@�]5��}�NzO�<{1��69��!�֡�����v�x;y���rv�ό�\ϫ�O��Ym�Ts�q�����\Y[��c�b ��dP��$��u�#ɣfs�����,9c���TY�0�r�"�7��#��!���}h�j���h���+dt���'����G�������hP��f�r�fB	��m��O�/v��#Қ~}'�:�����|l�N�7>XǓ�A�Y%�N��$&������w����0�*~�v,n+(ܙ;'Z��>'�d��\�J���q֜V|����Q,de��Is��ޮt���])��W[�\�ĺ������R�x䟴��x�5�_�q���[�@��O��T�%�ϴ�r�/�zʫ��Ă��e3��2��*���Km,Zd1H#h���p^yR��AT]��wV_�q�7#I�	��p2��7P���p��u��e�����8��m�x�C�� Ny����Vϗ��_��:F&�ƃ��6uF]0����?;���S�4r���i��O ��U�W�>��~�����!th��]�B`�Ȁ�`��j� m�r�"��5(����k�DWNi�Jm�I���~�$��;#�����%�,��4h�9�N��O����[�]+Zp��u��Z=��L�.�>Gh@�/tC���d�a<��e	E�����8��ꖄ�F8vei9i&���Q6�eF�ɘ�T���*�]���w�Е��rE�e�������N?X��yyq���`h[mBS�
�R�Yx_����K+J�D��׷q�<|�]P���L�Q���j�3��3S�}a8�
�X�h��g��e5-A���@;�e���p��.۸�،�6Y�~6�-���X����� qQ���,���͌)m�Q����Y�$���jn�c���h��[S*�^_^걨��߲���-�n@�SD]�	k�`�M�;e9�V#�v�xU���f�.�0�%89�a��� ���V_�-0�.�Ul)o'� ������jת0NG��mA�GG��B��_z
������e{K�R����9C���{�c�W2��f��P�S�g��T�^������@i\�S�Ђ�6?�H�=V<3�S�V>��s��i,b-�AI��
���u/}HD�#�����E��뙼=Nܾ�kDf�!V`*:�Ψ��eFG�yg����7餠u��IQ�4�f�Ŀʡ���{������fF�S�_zj̼�n�0��>ma�3�/���P�[�}��>J�'�s��G�w.�����R�o9_�K���	cǶ�]2wv�߾��+ӟ~���U�p���űg����O�勄��-N:�qP~4�t4uS���m�:���ȇ���8ٙ��y��s��ű��h�-��t_����Ag;��+�)�]s�м	j��`�!�����c��0�6�75���^��8���,� &����	sY�tu�j��=%�ȴ#ҧ�E�*0�Ti��� �B��๗q���j��*X$)c��v��[�t��2d�h)/uY^<���@�(���ejA��pj:'[��k�4�f
 3wL�5���'�F@=^"N)}Y g�Y� �D�(�ǹ%�x��p��`n�������F��k�E+��~&�ͨ$S���]7�玔	,�;-p�ÉF!�U�<���U-�dp�rq�'�F����1��y�/_@a��υXp�K���F���M�J��BM&��$Ėk=��m�y��W�0�cE��^yy��9v����fRΤj�b~�ޅ��'c-���n��u����f_	���Zk�X��?���L(5�r��o�1C����6	��<؜W�`�4+k�9�\�(���Ͽ}�6�1����6�Cet�đ��U�>����n�����"Bō Ӂ�b���{/���!�GE��$��%k����B���ȾTy����V�hv��U�8yth���tb�kS�U���x[��^C���#0�ޕ�:s��~�V��ZN��괶�mVf�v_� } ��\D�a��@�ZE"��B㏇�HmΓ��U� ^=���y݊�D�l��i1����|���9(�p��pdN
��w��K�9����s҇���={�l|�xB�d���o���b0���n)�i��s���a7 �ދF;K�4��3ԑe/u:N�]d�]Y�c��\����W��L=`�|q��	q-�0����;uCʗ��-�u�����N"��|>B`Hg��Vw>��Wy��}eu�|���y[2��=�|�j��Zw���@S��
�� �K�<	S����{+��xk�	)1*|މ�,��X��@�ֶS\�o���C����?�Xt�ސ/��)jm�2���I�!�W,�F�ʁ���s(@�\ ��^5�z[��ѐB�Gum)o�H�s�
�7df�usf�auo �[��v.��#7��\���Ó��)w��Ρ�Ȟ4� ����e$�^*A�'[�pӕ��0L-���"#�*.��+0m�Ȃ���d&)��Pr�o�5����H�Y������y�s�J5-������є'_O^0��z��k*Td����O_��&k����~h[#�j���\�uY���_�;1�'��̺��ߣN?9���i5A޵t��u}�)v�B�n�4��w���Gq�9Mu����-��8�*#�F��ڈ�����΂��t��[7��������x����N��a��<�/����7�(��S}U�A�w�b��H\%;��X-�L7q�Ɔ�>br�;��g��,��֟���zAw�6�W�L��麈Y�`p�|n��
�WAƭʲ���Oi7� i��I����0Q�r������8�zeY;`�5�b��uc0z{y��$�#����(�"CZ&H�$�);	�(4�S�N�8�k��g�Uu;s4V���*4l��V��;�z����\��P'��#W)�
鄏v<��2� ��{�4�I!��Ub�h�悛쨕 T#��Hܣ�H�b0�L��h��ޞ
C�	Q�)�)P��ߖ�u����+&���Mzyr�;�@�AG\��%���I�bZo���$H�����L�FPS�{���bD7�N�K���I�W��A��J�H��rMh\�Y"FHЬL�g(��[����$W��(=s4\�$��my~=9�֘l��aa�[�~1x�q����7�K����ۑ�,��ka`���G`����ܪ�^?m絢��p����VY䚗)�ǲ9Cib�n�@NIY׀���2����Ǯ�A���g�A�pe(�4�v�פN���VJ����v�W}�‵�K;��P��lgI����M������qՏ�'I�9d�7]�5��y�G�
�j�݃�t�n1�})�jP{�ۡg�.�B��u�=���a�e��=�qW;V8�����'�3@��|�>9,+4��7|@�� l�ޘwf)���+{L����5o�/?�V�Y�Y�`�Y��02�@�X��aat���B�
s`�J`�4�0�{{�f�;�Y�D"g�í��i�!L���q�8����3~�4H]�&��=�­ʆc#'&��^k�eV�{\��
�{�;s�ض��r4dz��o�!�r�^o
�#9%���ӥ�ϝ;�����ݝ6�2�I2.F�E뻋��3؏�{�)`�׋$sCp�E[e}r�f:�tI�b ����v��K��neb}�@�4�������y>-�3�)��M�I�ޕ�C�@��8؉6Q尕��e�+閭�$�a���lj�z���(�Qn�p���-<�(G���̆9P/�,ׂJ��,��#������)����!����р`3Ýu@]�Lq��v\�۬Ay��$��d�(� [��tA\^����އԱ��lt�T�d!��r����Ox�������XP�?
�G�Y�P��M"�p�"�߭�/�Bt�/$E��;bi���7�n=R^O�t9_%z7�qBo���$�����؃|��W��0�f�O��C�|o/L,j����?�
C�ĥ(�ޞ�-ֈ�f����%�2��&��?=�2�t�5��-Ǧ�VsF�e��Zwt���E*+�̦�L�;þM�����,9.���"1�$~�����M�D�3
ꘅq�iË#r���C�0s��!�<���'ki�������,��.MAd�}�p
MG6v���o:
SDs�=��R�1<��Hyn�n��;�2d���E��g]/����>��:�a��Q�o��dY���f�z0u�C\J�=9��.���ν�����Q��p��ƻ	K��:�01��-$@�,fl4� u�鋏&w����H{eQ���$�m��!�� �T�t'�	<>���I4L�%by���a3Kv��@��te�k��*9��eJ�Ul�9�6�b��.*��a협A�,F@��m+>��7D��鈅� ��޸/IC;��p�����3h�.Jǃ<��*�łz8���K���zK�O#ɛZ4'��}��iCW�Gi�,b+��x���@V1YQu���g[h�8���K�wO�gs*��~>�6����<��2E)�|\�|�$g����o��q��,c!����|Z5Z�d%��!N�����E��Ѓ�K^f-������I����EVE<�1���U�Ŕo�J�����|{��3�����~.�1Ss�5��l )�����S;��38!30�����2�����B�oV{�a֧>�/?0B�z�Z]$2�̻3o���̃���Fe�~��M���Q�N��)���}Aiѣ��'^����n�����q7����*
�K�@D�U;h1Q:���}���,N1��bt��4$�9 �z�ԮCRE9����,����I��2������B31��z}s�~�����U���2�`5".���0��
�|����ả6-!bm���۩�J�ZYo�8�����`O:�h��� 7�or�]Ț[�)bYu,_�i�M"�ăh���<<R/3+!*#�[��1��)�g�X�9�V����
wB��$�
fQ*����9]�3�{�mQY�	q4��sp%�c�{<H}�r�Z�i0G>��4��#lДB��9��V���,����Iu��'$��V�L?P�YP�t�5�"��f׵j��-���_n�oz�;��\�d�����z��Z#Ah��h�����)�]	���`��i$�Y��F�X��U���ϲe�U@Z%�9D�4���=v���|��0�_����7���5n�!O�j;&_��B�۝U٦�!F�&�(���K>�E?@����{3���_�)�+D=8VH)- A�*/骖�t	[p@*M��}�!�2{[�7@ey7k��_9����_W��-�ٱ��8x�k�����*z�����SV��P�;�2O�U�m��$��&�aL�Z�` ����d���[k�L:���hp��.�	�=#vBF��e��˿oLZ�P	�7�����}.p��Q�h� ���x.���,��[|ǋq,kwQ������i!�^?k������a�8:*Q�3�da������C��ɺ�eh�'߱��ɺ&��Q����%��sSĤ-Q�p
P�%l���]F:Տ.�U�	]W�C��"����y��m�n%�!E��J�J�ф���4v�(O�����g�u�ҽoϤ>
h�{��}sʐ�R��~r�a_��d�H� �hM�:�Wh����=�c�,�����Κۄ>o���c��b�~�銤o�_�K�"�)���c��{mcD���#TS=,��t<�4.g�	�����ۦB��q]�<�1�_Z2Ϧ��vQt�������Z�s� mF"�����ژ��I��Hzr�*�ҋ  Ⱁ�+є�NK��2f�PҜ�?��o#�j�k�;�$s�:g΃�!2?�rGY�㋑T�''[N�^���	kr��s��(8�d٨F� "6}����X����R��������s-T��c�>_��)���ϫ���W�&����`��TϜ�$|�x�3�ں(�lq�`{�Bb�y1��h��� goVo�J�mk�W�7�`s�a�ZY�"_�4��c]ކdQ��l���B9��@p!���Lζ9�����ow�E�8�1��Ɩ��ۍ�03V�x�%!�M�ߎy)bF�b� �y��~zl��xR��ku�T5����a�� ����~6{���c#	�$Ի���,YB ���1�&�L�2�O�}o��"�c:���`� r�M�ZƝ�O��}Zh��Z-��)�יн��}]�]��2���m0\j�s�|�i`o!�"����)XK"A��ry��,Y LȦ�C>a:�S��zr�8��0��a��uF{0+��,e���m��<bD�'�p�]�X��g
�H��_YgS��@�;�W0���]�/�h���
�T(���h�S;e1б��d53rQ0����g�l}1#OQ$�����4U�5 ��t~4�����@�o��ń"l	�9H!���	ԧB���~��{��]����zT�m�">���Jv%Vtu��n�gg F,6�t�I���p�������P�(&���t��#�$[��"�{����;�%'t/��� ȥ����rw��9a7RA����D)����y��f�b�D�z���>�d�ƥ�`s+0����%!�0���l���`�Z�����cd���N��	�+J`��c���9��0�t�w�f��j­Do�-��=�nj��y#3ݼ}Ђ.��'+�����Y���/�W�'B���U �*�,���4����$o'��+h���ʜy~�"����u!y�v-]�ٯ�y�ɴp��'��[�!�*`?�w֥��N�T�e�v}���K�͌�}�5'�,	���(��:̙�����:���	ӷQ�$\\޶�ұ�@�}N�
%�k�H��2�պ�9mh3�u�u��Vi*-�W�_J}�W����n'*
|�k�>��,�f]�,�h�!r��5������1�W6���M"�"���p$�H�L�zd˅�UH�Om�lt�?���)�4*��Ȅ��B`����&���up�'�_i�@60��1�N�h�_�R�ڇ��w��?t�^�b�ܷ;�^��D�z�;����bJ�����f�ʳE�_���Z�t [�V��S��S�[{��>�������h�*��{h���4"��G,��V�j���:䗳Eu]�D�ܙ{��^��+V�RɊA�藚g�������=^�5���#��O�#��f��]���|���6���8Y��2���35^�k&�b�� ;q�Lf�2��;�n2>���δ����,��1�,�Q�������r�~�s;}�"�C���h�G�PP�3\g�b_:^ǫ��%;XN�8Cy�T���&`�O˻+�b{ǀ����zF���[9�S���@�?����&���jxn!�Ϗu�,�&�"�H@-�D���Y^+�!쾶���z��E���f�1^�`��C;�؅L���;�>�&��h7�:aַ��ٍ7����zOH����Y(%$�e��i3�5��XN���jȑ��h�P#��>s���Ä*�Vӓ���돻��jN׼;
]���jv��C.��hA�|��5fb� py\\��Yݳ��?��B��3:�l�)�������E���Ǟ��m �X���lM`��	x��]�h)o���ٞE�o>�>*D�N^�Ur�#&��]��Q� ����r�W�Bkm���L���ig+&��u93��<`0P`=����H�>���80�P]�|9��`@كrU}�$��ۍ��>-�R9R��^|���Z�V�5�U��7����J��T5�ȧ�p#$?�FTf��0�v�Es�x�;�Μb�A�3\�q�^�UZPP�z	v_�j�Ժ��g���~T��=P��A��(�?m�1��)�q�ɜ�騛#��|��kQ�~zF�������%!�C��z�劭p��}�d{���1Z�I�DH�k@¡�5.]r[ĐB��3���wc��� ��G����0�w *T����l�z��eb�l�<�m��B@Ի��S�-���8Sk�vGU�^�)DdS��l1U��N���J�o۾M�phs�d����%��[�JI��D ��7�_�#��o:�n�4^���y���}[�~� '<چ�)aA�����|���O&u:���Ȕ���� ~�'sp����?)������?�����&��@g�iul���{}���YO��vbg�y�����[Dt!�������:e�������-����,��F�B����b���f�d@C\A�j=���ɷ�a���z�"_x��)�5�F��9G�q�N�v�-J���O�ڃ��/f�>B�����%���ؗ(��2�W�ݓy��)*���zP��=�̙x�z
�Si�oZ��������i)��U\d5�/����f�S�m��2��=�)k!�KfH��ا�R�Om*�_������~��D����W�y �����_����'i^:�pc*���l��}�*_$jea�,AYG�4��_��V�;1v��|�:z���r[�q��Q&�@���~1�˜��nK�_�t[��C��SIw� �"�/6&<v2U��p����TUa\!�e�Y"�1�iT���g�$�hr������/��M����LXC"�Ϸ�"�|���B������z�.�ܜ�:�O\�K��b7rYJաd�ԃ��z���QL��[x�JV|�KɅ2j1��E`j����m����G����}�V��1ު̞>b���X�s�V,�	s�g*)ŷ&�?{�Qd���;��'�ڧ�H/��Z�.�zIy���&� �i<�mk�#_����'����E+����c>�8}}hf�����w�j!M�X%V��8*8��8xx���z._�ye��zi6��_[��ˍn���:	��`�>��v�2 �-�(���b���|'�����P���"�ȩ���(<l�+2�O�GW6��J8~ؔ�NS|�`M�]�w��ŉ͂��=�窉�[y��PU%p_h�m]:d���Z!6gܤ>�EZ��.�L\E�]6`#��m@Jn� ��ffEI`=�)��8Q�u�̲a5�C��0 �P*x�")�耣�Q<�{I�j�/w\���S��L<���3|�3���CZ�m���,rmO�ns|17�O��FX��՛��;Un��5�8)s"J|�=���<��qA�W�{=�����ց�Y�9������P�y���?R�cR�>];�ҤG�����p�Z��)P
x�ok�zմ�y5���$�� ������1j�	���>��������:zq�%�O��b�<ҩ~6�s0)j�C�o�a�Z{'��?� �.�Ūt$��2w���$�>�J�V�cKv���ځ�וʆ���O�E�ȳ�3�B��Ln��]�~���=��Е입��K�n�hH��og���7�}���5e���L�X��^;�$���>r��u�X0������B���'̱���Q��V�3�9RFj�nG�����ՁX�Z2x<[�����	��BڳV������@1���ԵN�aaρ����T���h���Q���<2���N�0��3�����dwm�燠y��9���hC�s@�DY_]	�oP��G��ݤ��K���'7��[{=�y�W�+�T3'?@�[ȣY��L�q���L��JgZ_�a���c�����|�7z�j�3�j8:�+�Y�:ɃyX�`��+(6.l����{�A���ۜ�v�D���C3V>�x`�v͗���$��`�s���ۿ@������ؠ��^.f��S��^7x�YH�]j!�1��G���{�Y�M��v�zǺo֧���ݭ�]�;dc��̯?�󪱀��F�=��%R�%��'H���dM/4��Y�b4��7\�F{������+���f��8���2Xm�~��/N�힚d߉2L%���n  �v�M���[�8�)/��{�18Q=}r�jL	���C�8�x�L�wbo���tcJROd��ˎ��n�蒨_��b"��Bf�JwI�U�2��Ю�z���QC�(��:Y�>�����VO�ҐJ����9N����<�V���l�,P�	�y�A��ߠj}�3$D7���q���J�q�|�W�!M?E��9T"i��מ{��^�5ϣ��j�!M79�#�� �l�U�Y~CX \�����r����ӹ�4eD�ʋFX�v��Bkܜ���G��xb�G�T��-�����.�M� ����9h4��1�d�9��V�i�*���s"ν �!�#gRK�ww<��SE�Հ���D���T�;��rqQ��|���}�c��S;Yޡ�JM����D�߲�{���#�`�s_P��ͥŪ���=�K�����=����?p�Y�&����bs&�M�M,���m3��u~䌿X����u���֡1�(�UVe�/�BU�v:�ٖ�a�R7g�>�K�@��!Xn
㯽�G
�jY�6��t��L�9@��)ȝ���$L�I
����0�U�����m���ks��HzLW�=����*w���*Ɉ��~j��$Ƥpy�,�=0RO��T�÷�kK(*&�a�iG&F�����E���R��2T��ͣIr�z�OX��X���#>��� �qn�v�H[
�Q���\,4ɦNDI�t�~���=K{!$iibt���Q��x���Z���f�ĝ@类�H8g����mЌ9�C��b�!�*/&�^A��Ϸ����-Be\(���u�T��k�v���B��C�SJ�L���NIܱ.2�Ӈ���K8 F�	�J��@�\w�=.�h���^d�6�^_S��N*qh{s�Ʉ ��\�$ԝ����('�xSD�8E��"���5�����VU�HK5�T��l����i�|�m^��41ݨ���ʚ3
	�t?ٹD]]��0�Z$�7@w�6IEv�hZ�G�"�J�87I�\ܥ�xB�Mײ$�\ܰ"&m V��;���
c](��V�1w�ڍ���/�i�^8��������3�^��.�
��t�iv�65tA�ݗ����sa�����\�'�}W:0*�9፟�_��������h�[��5�i��"��K�2�Iʊy1U�įQ�.�Nx�јH� ���g@��Nv�y�<��aQe��&�Gv�C@��M���>vd��̂�>wy(̼��p
�"ni�T������4N�����f�f� �2�$�:�F$����j�����ݤ�f�N�7>w��5)G��t�b�[���6�g��;���LRB*M�4�_�Le�O��.q.�(D�ڇ�m��(Q�0k?��Q�M���^K�)�2��nP3ơ�ē#G�ϕ���٨�j��Dy{���E(����
^���B����${���^
�1p��{���V=T�}dt�rc
���˦�M��[q��/�Q5����C�P�\��tWkW��@�u����� ��7���М�Ȳ=���B�E�2�*R��E�J},z���$$���n�ِ�����������Î��2�Û�K5]��3ŋu�����.[H�0uG�E���=H8�(�Kq�Q����g\`E��H�w�]�`�����d:j��^|w�腟5�?�k�:�,�ۍ���}'����,�݆X��������8�`�ڛB�{4
ށt�Ie3d3�������j_�3>��W�|��^C�������ݛz{r�f𐫿�G|ڃ�����H�{�Z�s��㭎���aV�!���ͽ-v%꫉��%rbyw�!�diX�Iڹet�Q��YY�|1���(�L��m�ߟ�)���俿�@壟�(V���L���A�v(�I�O���5�nn�?�k4Y�YJۛ0<��*h#���%Ϗ�� l S&d�q
y�cU��,=U�g����U~��m]���B?ӎ��ˇ�m�ީ�)d�'@郺{�ܶ/��Mr6F�
��Xkl���ed�%_?���w�(�Z��
n��H�y�5�N��P@��v��ݫ_	z�	����?�e;rb�:�ݐ��6?�i��bR�	Bd�%�k�Z<�4Zk��>q�+��V(���}�+�j�9]��ݨS�r�d��)[���Æ�#UM៳� R�A^I:�-=���F��r����8��Q��!Rgz�B��9@�&��5��.���������ni��)���[U}��^@�� �4�!��2\��-M����Y�1OyH��#޹H2�������7��v&w,�����F�P�����$�h�|K�3��m�M�|�}���YT�9�n�G�+�]J���C�q��a�����	A�/���c��?ԹNZ	]��0�p��^Ns�o�a��(q}�.�����*��(�':H55��n���q���
uc���mn� ŭ<`�#cL�x�z�Eؘ&PE��I�T��C;�e)"�n���35q~�'y'O�	��Wd�x�y���0�4�O��L>f\�	^r�^�h0T$G?�	HP���&���]�38�h��%�k�Sy6��=�����6��C`t��C�s/�X��؇aK"�2���P�&مV�^ư>��6�^ůa���W�5#:��&"E�ܬm:9j9���d\u��6�Ai����t�<Owe�~��Ne�?�"���C��y�����Ma����IK���ߺ�y�����r�M����@�����FC���<"�A=����?�W�0W��dx�T��o�oFj�νr�k��G��\(R��s�ӵ.T�bQ���=g���z,���t$�;�@��A&q�'��@	�Vtvtl�ɛ��8�U��#�NZ
3ⷾ���>������5#����p�N�D�S'���M���d�\<D\]
�����/c�},����`�c0��-&���z���s�$%�S���#�W�=�����o؍t3�������%���.FZڐ���Q�>;���vB�C�%C���𥔦{�r۔�٦���2P7��=�s���
��J�E�8���.�d���lK��ja\�M�C�C�V?M�����=] ����si�݋�5�w�;y���K�M�����i��7z�Ӆ�zT�����|&�	l��o�o��cdI����w�5��(�)�.��A������JM9*⮈X��b{8.wig*���u7e�ro�	�n��N�o�ca������=c�-Ŵ����'�M�L��2�9	~��1�$�9?3���\;\����*5�jłM� t�ҷ7�RJ8"$�/�ى~P�~�G\vf��ke�^����;L&}u�R�����	9W^��z����6I�����궛-/3;�hMA3���Es¾*���X�1�����g��2�K��c[ϲ������^��{G�(LP�T!�ɂ��RkT癒�KO�O��z� }X{-R�a�(����'�_��X�H;;<�W2h�$M�5}>W�J6+ �܎�@�I\˨b�3�ÒI�.�"�S�!�t��\���s� ����ge���wϜH��}��z�,1>)�d��"�؈�T�j�V�`K^l��l�	�6��?��OJ_��1Oֽʫ�+E�e��1�� !��TՊ`���	���;u�`�i���Ͱ���;�r&��<���(#bj��N7#a� rt���k�E�->������0�<5 �
}^J.����z�F�s��E|(���vV�r S!�By��fs�H�����-�W�𱍡�
莔VӉΛ�-+��z��� 4B+��e]�
9�}f�i�vȑ�Q�ɲg���O�\�R"w �����{��[:9��Y�v�9&��������h���A7�f��.���������|�S��t�+��F~��	*1���HNK�~�2�H������Dz� �<������{�t���^)WƩ1k�0����B�i�ߺ����`���\|�zz����zwȔY�um~7W̡�?" Ҽ�Ӫ�Q� Cn3��J?�;Ԏ��ͻ��<���o��	�/v�'TsCL���<�R�<+)M|��s�ayz*U�TT k���+Xc�^ɐ�ky��n�Gc�	����5F=��9��L�$��	���,�R��;�^QA���\�Bm����*�r�N�h5����Z	M������Dx�;m��:��3������J���Q-?��t]�TP�*�҂�s2��4���Q�����G��zgG�j�ł��$�V����yЇ��*�x���<=��v��S��av>��UuI�j�  �]ou�/�L(#��V/�ny(h*��_P���5H������V7�L�ô8��ɻ\߯�����|\Tị�\	����:NQ/���A���@F��8���Hm�tމ�:>�8�;�	�������by�V�j��A"�
I2-�"U�V�U/8Y4��p;ٻ��Y�R��!y� GS��<��z0'\;��9Y*�帴���F����B��K?�RRAa��sI!���D�gi�Y�-I�mM��w5���
�avԏ�JÆ�Fd8����H�֞_��6���Gͣ�r�K�t#����GL�M"��.E7��u׮h�����y��f��ȇ��.|G�����i02�e�6fp!�� D��T_G�Q���?q'Bjl�$�����z��|:Q�	r������D^�3!SW�.��>G���_�GHN�����/D��^^�A8Hk�~�z9�v���_�����xN�i��3�I��i��{k��%R�4���z�w[إ�d;�-�y�.��%�"B$��-�އX��R�$���GA^̥��O(o"(!��cT9��d�T�m��g;����Ѳ��k��$�ď?y��S?�<>t�A��Ю"���g�)�c���K�2Z����h�̈́!|�c����x-EL���S8�QC�c��;v`�A(���9�F�;�X�O\^ZϮX/Ȫ<c��IĿ='We��1�o	1��ߒ�"���Q�)4�9�3����sh�<U�L��U!)�aܔ�J�}s" �#ř���G5�l��vg@�X��& 	�$�%���<ߴ]� Ql�P��r��w�WF���:p��yL�|����4�x*�7r�1����FG�p5��=�uƹX���6)�zY�-K����r0�
F#�L��7����|�e�����	f��u��d�jz���4�-�N`�9q�%\O[�w��P�#���:v�m��$���f�؜ʤ,R��Z�ԈGI���/�W�֤)@f[z	T6�O��+r8���|��ꍋ�+;��	n�a.�!�W<�p
�QBM��%]ָH�y���Ӟ1uo���A�I�H�x��"�c��Lk��=q~��K,N�C��3�_�~p=���gu������������!ȇ"@_{�9[�!3�W����?�4��I�0~%m��q&miz��,9�z�?�:&1�Z�P�f��yl-�x�}�J�=<H�4�rT�U�����ѵ�@Ǝ��:�YLp��9x�T����d���c�4��.��ZɀT3��d{'��1{@s`�W�4�A���L��h�=�&7�3����͕,������;��/m�#���(�(�V���ז}x�h���N׈�����tt=R%V�9;eL��m��лE�	/;�34���e�T����A�I��	~T��<<U8=�-����N��+fxwp�ި��_�E�C'�299������j:��>�p�V�1."�q��̱�_V[�|n@��r�ũ�d�l�<ҍ�P��J�D�H+��_��6
b�n�B����9�ſEK-�<.@nx>�Ŗ@��<�Q�Dcҙ�%M-@3V�M�S����G��:����Pk�����s�����a
-;�>�}��}�{��z�a�j+h�a���a��*��45�Q=JL��c�Z�F�E���o�!�.�@�`A8PLU��M�}ey�����p���͙���kj���ի��
�l9�w�;�t���Ws�y�5��x�irN�� s'8/"�����o�7����@�y��@O߹"�x�{�Y����]�Q�I+q��������s�8�TZ��O�@1�,߱��%�)�~�hq�&�2�Y��Q@�Ȇ���٘���YX���)���c���Q���5��~���zF#�M((�V���k��Y�I�q��{�%F��c�.j��3u�@h]��$����	�@F;%����̂�>�E��m�@|�ϛ�?��h�S����d
�J��?0ZE�+`��m���H��3� ����JG��t�5G[Rm��Vt5Z������p�i�Z����W�NYH�\@E�R0f��/s�+ �&6ֹ�Д�"Q
�v��@uY�	��Y��ѫT����rx�F�8muZ+��߾R-$���ݡ����q3"��V��-�� ��%�qQg�𯃪-.e�P;d��O�˃����NS}�dy�q�3|���阳��I��x�yl�:\\w�D��8�ܟ���Z����G@��(��p�	A��O���W�}�s�Yn_�z�+�ץ�=���	7\�W��!�-A��A�, �6t����Q�M�&��g�ɡv�W[�`�إARN$��]���J����#�E�˝�'�h�rf�R�p�*�9�-ádp�q��'��3Ȧ��.����dGq9v*}���x�6�Jea��m���qt�k ��5���c��-w�%�G�"��J��Q���Χ�ҳU����a�h��g��V�lg� �I�2P���4ޠ��1\i3Y1����&d�J��^k:ޡ4I��}K���v�����qƗ��V�8�h��kz�n
ϸ��^�Ƴ�#h������;5�r�z����i`�a�|�e��ɧT�U�;/X��nf����:C�\�h~��-$2����^�tj7X�䴩�iW �����*Z�ڄu������#�4/a�ãM�0@Ͼg[��e��������8:��.���!X�9-���e8�և��4�N�����w���G�j��+�	�T��ٟ�AR���TI-�����Ax�\�Ί�a��<�`�����R� ��SF���	w���=r�,�zU$G:U�Nr\x�Lφ����ⳍ?�߫�)Dl����b+�6 i�ZDa����H����������my��U9)�͞�qE��P�;�ׁ�R�V�׶v�f�F�W�ޕ��h�)w�o8Nw};o�;�p��C���N�RM��z6�Ю�v�i�DQ���A��6@g��aWx}Z��6�V��Xe���6-�d\l�-�r��C���i��%ƁY����!�U=9�k�$���-)��_��z�B�qh����߅+���[�7�G�țyU�_T�-!��31��s��^����~k�@����쳛���iy֓�>Mb%���a��,��v��i��@���߇T�0��+8� q'����b��?Z�P�I�~!�Y"1��g��F��~�; X����m�<pb��24�-��H�	56�>����>o��0�3�.�܀�;�HS-�DQm%C��p�Ii��gi�Y[���
7�A�t�Ʃ�PʖC���a�A&e r��4lc��QGzEa�TR.=C�7�5�[Q�L^MU^��{]���šD�t�"�'I?߆�.��_��M/D8[�I��(|�����nC3W��MBZ��"T<���,߱�gj"/G�#a��^J�^�	Y!�T������G�	��56��O]�Z,D+߮q4�%���$���xo�y��[�G��m;b���E2rt��,��q��i�LQ�I8	R��]�1~���smrk J��3��%�9ĸ/-uv6C��G���ԥ�\yzt�ކ�.��nÃ�}�Ҁx7/�d6dЦ9E����~h�C��� �u&Zވ׹��!�]����T�Lǈ �^H+���=v�g���&��<"?=k�
l����}~m��ߤ:�V��>�g����`:O8&���/J|�Ƒ`;(��o�C �?��C:�çG�~���tc�����
O���6Ww<� $��[�ss�'��NpJ�gM�y!�Tq���� 40�i]��̓03�g]��6hWN���ep)�%�B28S29�B! �v�F��2�?$��@��k������TF%5Gb�#�h�	?$1�k�)E�����#0��g��Fd,��D�&�V�k�S�[�)�BJoye�6"m�[﨡µ&�~ �jibt7W�����5KM������N̹x��j�;0�A�Ia
�"��iKǟ)�I�����%���� �=��sKi�E�˝ԡ�Z����TE�����޾��S��..)����=oB��u�ı�h���t���:�ZV����d|����q���x5�R�]mU���6"C�p����.�3��J7��?����	�ǄE�9ĺ�=k�O�S��4�D�f]��-F~V���!�s��o0�ײ��.��l!�ܦ�̨0��E'� Lث�}`Y(���\|C��p:� ���Y���u�������&�q�ϰ~\(� 7
���P��t�T�,��}�)d� ���"V[�M�4T���u�dj�q�B� X]���&�Izc|��I!�ç�\a!�3Iᖥ��c��|�#P8�ǧ�\@��IǊ.oSk���Z�\Ow*����+���S<�n�/�4���2��>Kg��	+�g�|��+OM���R��n���pC������O*QD#�wb��n�_�D,�2��ȋ;�����M����>Oʥ��덍}'e]�11�-M�[�O{��W؀������$f�ʫ˨��m�EcZ�m0jEu��;����a�
q�����3D�{�:���n�,T�	�)�1&y[qa��c�<x6�{�t�i]��8�gmn����qQW�ɖ����ЎQ�����Tp��q. �*i#�D���?�>�]&l��?j��J��0�t��ZkծY�p�Z�Z<D�~)���;� �K��E�Kv��9&��ʆЂ%��<��ݓ#���r�ƣ}�KW�{�|�J'�5z����N�� �xCpKS�	��0���I����� %�!��EX���VGFk�j0:�zR��,���������E��=�iikn|�x���~��0?S��*�|!޻�2����1�ΐ�Xk����W��~c�+*��5?k|�9�-e�3h��3�T���S|��}a���_�h��5���I��9��o���	��2j�erc-UX�4\�@����ͬF�
�3�-�z�c�<�5��ReQ���\�����FL��N�����p8%m}w6�����/Bb��Z����e�4����R�4���J	O�8٠|�--[������qorC��ç�%>B/}g�4m���>�F��'� 1����{��H���mH�p�b�Q��Wo�.	j8~�F����_�.��oH�@A愑Z��/�����ޛ��p�$5��t�`�Sd�:p,Ϥ��0�{
�qh�;0�����?ŰP�����"Կҵ?>�,�45�1�!�_G0J���_�#p�����9�&���3u�o��!orx�a�G_ ��\~g�2�I�ę*�"�� ۭڋ3��L��_	+�E���n��عп���τ�~@jP->&�&ٍ?���&T��Ik��/c�23{�Ɔ��e&,�� �e�v�y�A��Ox ��݆��]8��*{W{M;
�Y8Bx2�P���u�ُ�x/�~�=�L�u��[�ʃ2�g��"Zjn�K-��a�z24�Z# 9�E�!�N\a}:$8�����/�pRi��Yut�q��btp|b�7��ø�I_�J������ّ��p����,�H/M���E}���T��b��w���1���lg�P�)4��N��GM)~�{%w��5I�6���������,���R����#��8=��z)s*�m��l�N��N�w����S�;[�j��2}��صS�S�d>z����Zj�WW)*�Ǖ���4g����wV;K�Gr{8}�s�������E�sP]4�r���dxɿ�!U�<=�M�.S8eo��8;E��K��CF��C
���)����~�Wj�4�IvD!GD�����p�
���>��D�%P��n��i���n�Kr�fL�,_bl�'� ��US?��������##�봣�y͍䅗Z�5��E��	�޸��~�*���te�xӻ���,y"۸|v���Z��^ب��E&���bVbK��-�H�N�YȐ�2�A�Jp"�0�c�Ȍ��������X��j,�AA��!�j�������ܰ�uA���z���C+����t�����& ����]L��$�M�~#�Y*c���r�@�6����Aށ���yRQ-7ļ.�pT)*b˧ym�$Z}�9��a��i9/�Wĺ6ˍM�D&<;��1F���0�t�;;8�i_��!sK��R�H�Y.GZҳ(�N�!��-�o>��.^G{�E����[����
$�*L�h6Ꞣ��L��r�PY	Q�Yr��}V�X�S �X:��ɠy��G͎1(o��p�:��+WQ �����v��,��$��W��C��TaT��ާ�{�kO=W�o�%��Y$5.)=Yf���nRh� ���ʯt՘�B�Z.�X�& �'u�y㛤#�W�5 :�"��r���&�s!ew�|k�ͨ)d'�� ��K�y��X�_�_���D�=�)�7�[zX7��ޭtv�[ �=�g4��~s��%���c�q~z\ˤI!�|gp���<{��G	!�8g�¾i@g)���k'����6ه�Wd�]�m���f�p������������5~;��Q=�׈`�,�����]�^��-�1U�2|.ξ�̷��DcC �jܴtA�Z*���v��2�b�Q��]v"��!�n��
NB�M*؝��"
�%ޣʴm����tS�x��)x�7���I?�P����I����ىF[L$o|�G��xJ��S!�Cej�<�om��D��=yD5)���9hO�_��h��21�}���j�e�#��&��|�G�)	]kGܲIS�,��e��s"���s1�M������.�6�^��웞�bҨf���n-0�^FI�A�v�H�u�[�L��︷���?A��.�{�	�'�āэ�N`1�oW�^I�V��s���;	�g&��5��*�*���Խ����	���xq�\�d��{��`1P
�ۣe�ȷj\�չ�����R�"�n/AH�Cz>�.��n��tc�>�@�$0����U Z�����bEY���*OX:Y���=��@k#�D2��� [�Ԏ���h@)&�mfl��@Mj8�͏n��Z?`�	Z��K�^��ۍw%�ͫi�vU�X��)9�����(�0 ����l�jJ6���#�d�k`��5���S���"�����Du���L�������+��P�ﮮ�%��b퓼u��I󜴚S���.�T6��4Es���u5��1Oy�9���;3�,Br�B�'Jt��i���)׳����O��o�})<���}P���k��9$������-x5;P0��V\���bsY�K�	Q'�+�/���+L6��� 	��#�����qi�c���13)��qB���c���Jؚt-3;��V�-�A�>C�����5֛`xA�>�K�E�F8��i%'Ta��Ǽ�ɉ��D+��j�[ˆ-{�s���_D�Z�z����YV~t���~|�Л)��U�-U�"��,���V)b>��WT�@g�؊j'@��SA�d��}	w��s3���K%ۜ�wc_���C~� �֯���W]ag�����>M� �����ǁ�d��!�	ڪ�1o���Xu���s/n�[����#B;?�:;r���H�{�|�*�/����IF�x����u��4�)���U��J�I�ʢ���\֘ǅ�`^x��d��N2�����uٍ��䲦�V������Hh�6j�ʊ��!�p��uw9A+�%���"]�H�tx�޸����5���5����X3�c�&yQ�߻�aMnWt-OWa�6%��$@�&�$Y�b]��f�TO���'`u�< ����%��<G�b�YĶǧ�K�y&�%i(��F���n��(2m���*ʜgt�L��n+�H��z\�",	ǸF��W��LdCh�"����J���v�����}Bz��f��Aڌ|3�43��g��%��)�ȼڹa�=q�-g��Ak$�D����+�5�.��)���(�1u����j�|�ul���)&x�v�,�Gwȵ�\W���`W�IC�bxO�{'��hD"�mxq�gEHx�{��t�l}��u�L$�TIZ��g\���;`h� �B� ڮ�p�y�T�%�,���6��̳�p��X��ӆ���ɷ@���idt���dށ�}�404y��=d��z0
�I�vǏ�t�R��`E"��/���=BK3���ꔂ�t��:�8��97���\L��tT�P/}	�wd��:��/���Ҟ��[��k2��n��,8?�s8P `�ca���B>��x�=kA��5�f�]��(.�����͊��
�"�.FE3�I�9�Quz����+RSSY����H����G���X]�[޲ۨC�N\��'��Mف0�,�'����~�nvu��Dr%��6�!��	 ��������������8�D�{���܅��E"x������灥d�R掷�1��2�]�����W���.g%���PUr���z��>�i���z���=P��%٤������@��.>cD�8X\ǫ�u�Zj�L[8�s��o��m*�	�p�O��R�rĈǲKj^�Q%����e�+IZ�;��8%@%Do����?d��^>�5<��VEumU�o<D�i��d"����X��2m��#jT��@r��_�lI���#s�c�&�
i� ��eP�h�1��j�xh<7gK�6�L��t���>����p�^�I�b�Ik��;�|���^
+l�H��^g'���k��1	�UJX��nR\��j}oT�@�ϖ�"�)�ha�]��%Oߌ�]��n��+}�jy���7�f��t����S4�V�X�����e7�4|����	�m76-~���x֍����W����,�����0� ��
�).���5|럡��ڲ�W�&� _6$|)�h�}�ϥz>������9
�-<A	wlLJ��-���4(�ɗ+��Cȗ��A��%�/�{�n_�"i�
C�ϥ\��K���R���;����p�G�w�*�"����0�e̣�����<ȡ���;��~W�s���sh�d�M�l]���/Z�@AB���؆���,,��:^����T�C&^���e�*^�e&l/��Aځ|I��3&;i����,�hH���u����P!,k���:'�i�+�����VsC���a�λ�4W)�-6[�yp{X�3Rb;�M( �^#�,���:j��[����;Q�m�'�-ZL3��y7���%��2��H�u��
�N�*�|��v8�����J��=��m#���9u�0\2F�L�)qh�q��+g3C�e[�r�@�\��ߦ�A[�����Wpyo&a{�P2�[���z�e�\��8>��M��DB��K���J�g���Q\"��֥�� �P��1�<YGh��K]6Jɱr����~�*���]�nr��[���8�����6g�?�.l�C?�.�L_�'����Tjx�c�'��&�إ���Bw�#EnC�����q�Q������c|�niӭ�3z'C�S8���!�*����i,{�U�S��+����79���o������/����N�[Ժ����b�V{�9D�t�Y��V:��$j�:�cT���q.e+�n�F��s��~V�5�����4M�XԂ�ٲ'�������礩\j$����4��@�.���q;:⒙��W�s�iǮ��G�[�GK���?}g���׍�ltdz�Zg;�[+B�H�J�t��b�r��YI����h�L�D`�:N��I�f��S�g�Hj�Rbw��Q�qo\����1"���ZĈ��z���|�yO焀H�r�l k��v���wYֿ�:���.�����ȔL00rr���Bz)Fa�.�
���ש�τo%|`�Y ���:�hbA�b����	뱛J/,P&}|��x��H��_:����2�&�
g�����,�c����\�N����ԇ��d���	/BݰC��m��Z�ʓ�4�,���pfrۛ� �>�ZF"9q�rX����8\�PdҞ
����J_�y��u�e�����}�j4J0&��P~B��K��2�4�d*�otOʩ#��6*͒���cSյH����-�t�z q���%�S_��q�v`�@xx"b�*]�m�3`�C����Y'/��·I�֎=eC�2�j�C���BL�0�D)7��i���K�.#(.y�fc�����^8�]���`%c�NPi�{�rM���E���Q&��4�܄%z $F2�+��'���Ʃy$1��i�$��g�'��N� �^o��
2��U�a�i��N3�&�_�r���`)b����T��I4�P�(K��P�&�����H!7�!�ٲ�!\�ܽ������y��L��ˮ �]�W^S�^�7��������^����O	S4	Ĥۥ��>�	�Y�Y����_��}�RW�Q�zÅ� �d�%��щ�_Y	iE�S��l�v��],�$��L��j�qp�_��(�yW�y���HO�Ŕ3&Pnϑ�U*��d�;d� 3	��<�
>�K���9�6��1@U��&$�I��7Ru̳��1S>=��^<��$cыj����j;T,��E�atz�y��q0�GŒ�I�:�Kb�}o��6[�������2�}����������<��� )㿛�ԍ�V�ܔi}6h˧nN �Mل4oo͵�^�a�u���X ��p�Q~�m��(�#1�l��gZ��#F����_�3y���5R�UDe���J�h�h��}?�ZN$&�I�+l�����&��&��§*��fq���C����?��) ����Һ�m�B�o�0w̗�G��m�} �z��؍��w�l�,:���\��!]_>� ���4�f�Y����{�w�y�,,�la��i����;�Zq��hr!O#�|��RF��'c8b�����r������#�U��m�3!;�M�X���z�Q���dL!:̆������`PU~��KN?^��&mf�Q+�xʜ�XZ��t+�l�S���T�a��w;PCb���e�C�.LφƦd�!�έ;�s�e�r��[\zq��l��2��!7N�ݗ�]_���t��������TQؕ��}��x'����:ւ��d�Oi��qu�8;jh�p��sɖ|������/��k�/S���99�{�����JC��d�F�@����u,���4�1PTA9�8Ϫ�^~��q7���O%�|p,X�=|7�'����+���'}9�.��b�YV��t7�8s��V{#m����RbX�]�����<Hՙ�9���־�zCK15y��㣭�)䊑�M�-9J<��o�Ǐy?�:�K�JqR���_����S0�,��$m`@��5?����d�q�a�qmZ[vAG%�Qa�����W%�#����
y��B�(^�����0���w���*�'��t��v�(�� 3g(��5��^��C$����r� k�����/}x8���6��)�߂��ׁ�a����v=@Q�X��XǸJ��`8��t�^kʖs���6�0H͋�A��>;�ʐ�0���u��{���
�P�}h j��ڞ�#���"��Hl��o��_��Їz�]I��������[#:mX"�3���V�Z�xsw>������OZ!@|sNt�J���V�˲�eie5َV2򁲒-R'�0@5k�n���]�(���%	�E��fd��bW���	 #����S� �(
&�H󭲟#N�"��k���g�y��H4����O��!yq���M񲓿�w1�%&��HﮧI����b�����V{�N�~z�&���uO��]+3�⭄k��[)0�C�I˽d��1�\�K����RB�o�D�8�JY �ͷQ��M�oR1����K)�Y�TdQX���j�C��������\H���j�}��,\^:�/�n��g4��U��k�w��|}\�q��zW�t��|7�LX��8���������4js��I��,���)���j�|Zhi�9���34��ȫ�t�1PF��R���X{YR�S��VMP3*��*Ϧ�Z�^����Ԑ�W����R� �����@�gc��Hu�����H��o{ԙT�}i�'���� �ZTK�g�C��O���v�*�ɯ�[H1p�qG�S|� ⚈`r/h�Uc�I��Դ��C9�Q;Мt-�0�Ma'�R���,��E�R�T7Re^���?�[���������b#=���WG�3R�5l�Ƙ1
�J��(�k�k�����1��v��Ӧ��]���:p
���<��/�4����J�&�P��!z��cZ�J)��}7��Tr����\��}��z2���i�q�N�����DQUD�)kz1X��V����Hv��Үo���E08.i���C����P�k�u��oB���A��Cc��(��T`�����
����u�(lȹ���Ū��}�����<�����B~�=��@7jr,3� ����~\0���v��@B���H9��Mh����6�L4jO=C�\�C�.9eݰS1���l�yX�2��E�9���0���B����F/�/4��%xZF���L7��9�]�4�:Z�aB�F�
��Z�� �$��b�����+��w��F%>�.`d��-F�5�3KL�]�Ĺ����a��V^�'a&�U�)��H����ӂ�̮�����%�3�m��ی�8ۚf(+�%5��޳��J�N��%Җ�$��뇌b�9���숾*��G�43�}��(���L���d��&�L~҆�����׋$�׭G�L�X�c�43k��
V~����kQ��BY�`�*)C۸�����s��X�L��n�%ŏ�C�Ҵ%���|mz�,�
U\�96��K�d5��nr��2@ۍ�$�}bI��w[�P�Rۖ�Y.%f>����L@�/�4U�&Q��@���7܂��d�0���X��)��P�� bM1���ݢ�*��3�+^��t'om��P<�&����SC����6M!P],*�N���_ɱ��Yh��n��7��B��z%���ՈL��	��8Ik�"N���+i�����N������2d\��<��~��b�¿�F�#���v��DK�@5�����	��.�p�� �����\�P��<6-eR̓�<���^j��Wc9�q$dn�\��~kHx�����o����ldI�^/�|�i��`�jR��>��a�m���WC\����<��3`aA;��"[��!��){dF�q��ٚ���O����) U�e���\�N$}��y�,�'J�������1{�%�����U�e[�QJ�Ђ�P-�+ޢ�{C��S,�62(k���^='v�*4��J�Y�����ٕ�ZGP��Y�ʭ��%�^�=|SI�9�aOi�`w5+��C$��=Bm�ߛ�Ǎ�<2/�[y�!L�\��I�LII����s�s���^n�55k`[�o�W�=�yp�M�/%�稶D����3������NO���U�Б�f'kү�7X�E'�oׇZcX1�5��O�aiȎRh�԰pk��sp�Ϋ��fH�R���M�?�?�\ihh�`§�keU�T�+�]�ׂ�Q�bF�܏��N4��&)�_�&�>��tAna\�^��@X		0d�a^�>WK�����*��H���l��	j?v�n ����6��p��O����6��� �:!=�W���w�V'���!��iL�=v�o�a�=~����1��_J&��_�w�%/�>tw
"����(�`�
�������?pℝ��C�f�0��U▴�{@�'a1��7�QQ��ה�R{֐o�𸜥��a<�ϲ�^x&�����Q�K�ͷ��gm�x�9�|O60��u�L�Ql	�����g�#D��g������*иw���Ֆ��Hry\��2\4�A�φ�@	�V��������Y��k��wS>�����:*���#}�c��=/�����s�ډlr�Au&o�*���2FAI)
���v�S���ʨ�[�8^�L��G���~���`��W.�999VAs�J��S�����e�=�f��"�iO�c�f�o���u�~I�k��y�Þ6�P�Ӎc����p�q�c����f��Μ��/�1��f� �L?7�\b9�˄����b������ω9��l"C[d#�m��ej4�9D?��3Gƅ�Z�
Ό]g������xy�����?"?��e�sI~�F��H)�)�D w+$�b���<@3���n"%����l����f�G2Q�Z.���0u�☟��d݂T�����@͜�@0%<,�I�Ģkt}簶�6��q�������?DzK�(�,ATf��$�;C2�4�m*++�����c��o-�Ɇ�aw�-N��p��%�'��-���X��JU��@8�EQHq�yd��CY��T�U�N����u��})<?,8Z!�[!�o�~?�����l���-�7��i7����R&2��&R3@��ڶ��o�-�6a�_]���#�O� K��p��H�uT��V�Y�A**|��)����N���;���4��Jp�;� #���aF3�