��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0���C	�i��E����`Zm� L�,ac�C1�0�[�Al�ی(��U�5�N��sB��{w��u<�L4�T����yD�YL<�d<���ਮX�g����������!��*v/{�"���!�1�'ݚ����������E���n�����Qئ�-|\Rnv�.�-���e,Sq�x,��Ie�����(��1P@��	a"ב���e�����
^�
A�O��H�}���x��]���ԇa*��M���ɛ��r�Dije��^G ɚ�cpqhu�t���fO���"[�Ϝ�tW�����ֽ�Vrf4;��J��s��f�ċ��� + x6B�P+�$U���dZ戯l�'�T���]��M��髸�D�
�����x�8)J�,��4�L���)��H�����,Uy���H��-���e�6�H7��ÿro]m�WX*y�A.\R�6	�S���Ȟ�d���������8+�5�.��c!$S�2���N4|�ih�p��Jd)�U2e��E.���eEƄ�� ����A7�so�*�9��C�Q����8��n�QrH��M@c
Rk����P[��xN�����r~�3���q�k�&f��o��u<�;��h�9��iӥ�#L��0�<�^2��P�'i0S3�:�rg��}j<|�w�ㄙ�ꪥc�H3]I�د�9�z�:�����wMk&s�럗E`v�G
�8	C	��]���:�q����ƍ�/���w,'�;���h�U$�����|�!�3O��0���|��%ooM�+��s�7��0�>�R2ә3T��!��t��{��E��(�^Dͽ#p�vC��H��i���|v�1�f���y�adU�W�|��m�	�)o����plT&�H�?��æ2�����ZEܙ�?���yx���sk]:���Y����b���JuԒ!ζΑ�qI>]n�����;�Ι˟����c=6K�fr���Ku��$K��*������y$_ȩ%K)^��a~AՄ�H�2�"��eEB��X�L�*�f�oB�
�W�5�`�&̃=���x���`i��Y�|���,�x�L�î���ˤa5IwLM����m&Pq�?&yK��Y)RBm2��`�l���;�k��i�`�R��^rS�k�'�M@�F�da?ץZS�N�3Y���,��0 6`-�P(����J�Bm�t�U��'d����E���F�u$x<�̜���)8(B���&OP���A�n�����#�r��$�#�#���3�*�p��8�nd�XNi�v�������X(i�����55���-�}� G]?Sݷ�:��D�(�\kgy��W�8�z���㹞z���Ĳ��w��S�Xz~�%R\M�k�ؕ�B�⺔�?�Ϭo�*�c���
�6S���\V� z�-G�G[m����!��&��V-?�ߚ����`��Dʖ`r�~��F����`PX��!ӗ��D���M[����u��Ub�OI�,�q�j�_Ǣ` \._k%������kj���K5pr�ϗ�&8����'F��S��t�ӵ&�U?K�<f�䊩��^D^b���;�[z]��f� S���� ��Z����ҿt��ɇ������8�Yw/�E��ם-�PƜ�g�Խf�LD\��^��Ƭ��)���z��Ŷ�x��8�oߓG��8�,��Y��� <yQa\C�.Y\F��L�~�J�(�1���&���vO������m�!9Th��n�aEz�}(���&�w.@�+v�.	ȕ��[^1t��p��1�B�c;~]�+�|`��׭J��,���s�"�yG2�϶����e��{��e�0̎=f��'�ׯ^�L0��h)�	B ��߿D0�,kl����l�F�X��N�z��ME��t���I�K��bI��?�(���Us��#���T6K�g�h��'l�BS¬y���":��΀���C�Uxu�Va���X|{l]�|ȡ��g�`���y�~u�+oP�װN,� ]�u�
\�Ɉ���	��yə���Ǣ�.]�椣>/�*�./l��2�aט��b,�,��Q0:�[̀�'eZ��4����:n&�Co�ᒡ�.��6��u���@��|��nw��ڵo�/o���V; �5L����o;���*)u�/�-P?'�|�@4����M4�f�I����,	s]p9Y�ul��Γ��Y����q$L���� 01�B\�hR���mpP3n�����}"�ym��n��U�-��UV�?�I��C�UkY��}r�S���|=��*w�)S��SS��͌h5A�N�Xr��Bw���w>/���t�� S2�ͧm7��\�+�wF?:���WٹCE�n���q�<��qyoل������=����wKG�5,�so:���G	I�$a�fc��vg��G`	F��4��`�㓴����JZ���� r�%�B,v�)���& ����y6��D�hy�����f{Z�{N��і�>t�>��ya�^J�@8zӔ`*�5��k)��.5�݄Y�\����=�#4G3u61�!�%�<�mo4�0����*o�&L��Q��~WB \����x�nĵ�vIÓ1��7��}�_���c�t�Ge���6Tw��~$[�O�j�	��qȕs�	�D�d�����1^�3�>FC�o������2��u�~ڏQS��_8g���j!B�x�5��{��԰�n1�Y�f�bv���U&���$	�VU!���0�j6CP��� x���f@�\m�u��I�$&��B��.�ԯ.Gd������<�����"���߬��GF�%�~?Ğ�)Lqk)��h�V�8yte���3!n����Z2�.We����=q�=)�K��Ŧwʖc�����&�C�k��\�k�<�b��s���ȵR��0Qq��!�~և=�9[���&���) ��pp���M3๑��Ǹ�N?wE��<!��5�X����-���^�=e��7��ϑ���w��l�V�%J킨g�V)i #����� .Ƃ�&�c������i8�lm���+�#��鉡���&C�	��!�j*ufճ&�E �$@��AIH*�mh��)�<�8eHI���o4QMeh�[�0�]ѿ䵦��s����L
�:C�yȧ1��k�ä$��y��z1����_�V1k_~k��x%F�W��
���!93��K�*xAvܶ���*κ���n����
"��;� W�D�.�9@�ݲ���2Wj��В@�{^��M(��Gq�ʬ2����e�X�f�gmw����"n�?�����p��v��H=7M�=�����؋V�?���B/?J\O6a,�u���N��Z���/�4���l٬��$� �`9&�?����/����R�����WT���MVb
��.���Y)���E
�X���_���
����Ez�O��p����Ȕس��T)a0 �&�>I��h
�TZ]�f굕�C,AsN^��|��$UI��e^d0��`_;Z�f�u4J��?�*-:s�G�>z�]�����p�$�6��"��tY�Y��`�y�ǭ�a~���U5a߿�!�;_ªJ�quNl��GN���ӭ���¯yU�J�0r�{^z.�j$zI|��H2�<G�8�%�TD���}���Ҹ��U��kR��=�UR��׵9q��>x ��]�z����)U����5Z�F�a8��r*�ט��8(��>;�.���ZŌ�%�������e57����鋦�u��o���'�\5�����݈�p�f�B�>���%����ԸwY]$�%c���.ш��0���[4�r�:d�����Lj;t��?� P�!��{�d��j%����G�3���'�����s���ي�f���!���-�N,N/3�t� ����x�k&4>���]�ز�B�@Vkl}���Sj�'[�"]Ѣ��B���-��fRŷ�Ā���8�ñr�C�f�s�F�B���GJ|�&��"#d#p��c]���	�Fkm#�E���[O�t�J9&u��Z�&A���=`u��u��P�[)\�8�/�G���S�u����\��#zs(\/��^���R�U�|d���>�i���*-�c�h.���j�$���l��Y-D�|b��Z#�_!�,�M�7i���0����n�>b<�r��O���\멏��r$1>��]܃���R$*y}%O�����lN�;�'�	v|y�f�z��Y�J�o׳���~�Mދ�e��K�1#�5  �<���:��t��=�-��|1S���&U��>��r��]AF���*
LC�v��������f����f2��fB����GE�q6�\���~Zz-7�N:�G�sh_��v��i��l��o���좖��\똍������nhO4�=����[P8{P�J��k�i��u
'w���ԍ���A�+0�=R`w���s�J�H{-��-��*���R��O]����P>M9Q�Z�`�?�T1�/�Dly��_�4mfa���ݶww��_�)r~�?x�t+�Y�f�+�Ff���IhXy���Vv?�o�����8��/��`6�j�Kd=  z�R���2u��X��y_��nU����OT��� ����M|h�a0"z��������$ xc�M%�*uNl�2���@n�����[W�p���%H���{ܒn�d�%qR���<UJW�6�u2�U�
��_'s	ݒ��%�?I�YA�d��u��:�~��sL$����3Q��c�i��������?��XFt� ����83�K�� +MH���W�C&�'��q�8����Qp�pSs@���5_y����G&e�� 4���m�oq��P^s#?Z���yd��חgt��.9Jmd�XYϥ>�~L%ԙ䚐0T�0T��U��A
9ժ���L�BJ�"���һ�����Nʻ��7���;`D��B�V�=�ʨT�;x�[eˉI60�����vGPȓ�2���?�$4��8��u���,���̍&���z}c�38��f�)O���7����Ks������i�&�A��+#�5�ܸX_a	��ڇ��9X���j�p��7#�?�� �c�:��"�%(��1
H��$g�v���3�:e��
�^��Q2�=PW�� �V�d�C�2V�$G�]f����^�*�&e]�5Ҫ��X�R	)on*����KkfJ��`3uIzc���-L;LN�?�v}��h��{e�*7�B� �L�?>Q��(�����j����|֯sQq��n��m�?���)y�o�r:��	��	4q�ġ�Ag��B����c�G>+mz0����%<zX�'a�=l�?u��'��v�OTS��1��1����wZ�،�&�����=��(yhY�T�P�ad�g@�������9Ȋ�g}iF�"���� FЏ�cW�ˑ̠J��)���� ���t��ӭ���d6S����j��8S�}ܷj�c�fbK��	�Tm;�Y̖.�E���B��q,�i��!GO")�jQ��/���V,�(;%�+��S��� /�\dv��cnb�i�"E7�u���χ�B�T� ⌀��fW�֖+q�q�x�������9H?ށ�.��4�����rHb�L�.��5�{���i����H�y��\� F���ޜ���9+�:�?�7�<s�Ea���B���p����������}��G�e���Te�X�����Q��ID����n7���?<N<���eWAÄ��P�%]��}�'�$]���m�����n�@�
?Q�|-x�� SsT�0.i~7S,�#��ۼS�V>���=&���(�H� �e�2(�Oe�el8F����.�p�_fv�H���I�2��s�J�l:�It��������.A���×̊�0��o��w}ԛ)��	�� a6�9�Ĺ�g��6�=`.���s�x�c������E�Z>{t=тR�:��F��ʉuY�5�!�t7������������gdǯk�`d�(2a�s��D�[F:�Y�V��o��.+�Io|X�t)���"�{1�PH�I;�s*ǃP )���2�bx�T?���{j)�N;�EU��d���	�d�(Ƚ$.��N�X�_��xjR�|�}��-��}5�c����^ر}�b��Dh���i]�/�07*�rf���No�!UX>d�r�R�E7�d��Pr�JO�4iި�O`/i�H"F�4X�۩b�������c�y<8xDT\лDIep8N����,���@��lV>%�F��
[��@�d�Y�(!+�1&h����Ι8k��Ebt�7��o:���Uʺ���Q�󦘜�3�аѩ��vm?Q8��9�:��V5A�����]�Z ���C�ѯح�_���E����%h���#��]~��_1��g��aP�!�,��w����"X��b�V�k�2OU�����=
� Q�Gˇ(�9��7�V�s�{2����O7��6�L����=@'ż�ge��i��v6m�d?��NI�_S��j\�����2�.�Q�f,���@�T} f D�{J_a�[�����5Y.� �
\	�k�&}&�X	�ɲI?�cx�څ$m���i��v]�-�=}����8�`>m2���x��e�4���#G���s��(��}�*���N#����\���hW�<� i�)j����ʝ	�����%��)�}���u�D���-����#�l'l� }�+s�l�cB��V�s�t�D�;�4�d�p�z�����s�iX�����T �&~T�d��nDeEj��hD�d�"��@�£�����b܀8R�O�y����&��P����0}�`�#��&�q���C����-�t5�K�.sY�Qa�NT.���a*ic.de-c�,�l�7�+��\��xח�%N��UU��3}����
vDE.n�����/����q�w7ĩ���ܼ���xȞ�x�U