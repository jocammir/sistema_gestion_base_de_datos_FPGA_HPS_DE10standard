��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0����_���3e���ӌ,n�vLUW*L�f��`�����;����yj�|
����A2��a�"�]7ή�;�7�x����)[�|dm��8�B�@N�4�z{�j����8�Jў��s��*�%z_����$WZٗ�pQ!l:߳4Ob�H�7K%_g�z�g���(����D�P������V�R�#�Ʋ r`i��vR{D"���~�]�Z�Röl���CS ���r^�Z��r=��oJ�l+V��{���)t�x�@.�P4&V�
6 >"�K�� |@l��S������Y���@H�4$,�Nj���-�`�koR-��!a+ug0�t�Q�L�&(1�T���A}NjV���$�u?��[�>�5�d5��p�����;j����c}�] ��@��� pC��������v��DDYl���iyH��p)���eiTvH4I.��"�����x.�G*A�s���,ڲ�Tk2��j��_M�O2u�LD�C�4 �G@6\m(��*8>�6C���+_Lx�C�y����#�<p�c�htkP m���Q�<�BTP�!@��]ªF4����� L�r9���9&V�B�:N�̛z�ss��J�//Sx�~�s�S�v�?�W�4{��w�'����~jo��ό4���S�L����]7rm�� ˊ&�CD�ޢ��{�H���D ` �ێ6�I����`��
4G(Tӆ�(t�/+���X��uy�^-X^ ə�㗴�S���R�Fk�&h�_<l{o�JNz>��V��ںhY#B�q�K�D����eF�B�Ӵ�
�$���Ƨ� 
d"d R'�/!�@5��ͼ�[����'����Kl\�qQ1R6���&2�ħ����4��*�mƳ��p�!�dm���{�����T��v�` ۷I�W�9|�z�#���#�"��������,mUܺЧ?�������K�2�1�gqlhO%u�F�3|	��l���O��E��(G[�]c�
�R���=�9}��F�i~�}ƪ�FǍ�u(z'�fwx۵t���妙s*�f\����{
�s�a�����6��	F��`�K�ň
o0�2����w�S\�7Q�n)�������ht��C��F��{�|���>�P�9�n@�8z\ѿ���⠤�z�>�� �^��>a�+��S����W:	B�#k���>�z6H/�
����*��Se�N�N�kl�F�z�������6���Kyi[��W�t�p���Ԉ���j�����f���`�v�2!��	�)��DN�	@�j�U-Ģ<��+C4� ����0��y|eT��ͱ�:�Ij:l��D��2[�����#(��K�̧�� <�~`v��ɟ4?�(���ܝT�X��h��Ͳ��\��$"H�8���fjq;�z�4=�%W�_�����F%L���K��۷r��<���Q�o�_/Z�Slځ{�dJs���]���{���D�����]�p�I>Ae��x9�M�z��uiE� ��{�G7����/F�:b�������\�����¿��ջY�d���fZ���#�]Vs�}e7�-�i����~����>)��טEY��&�r����x�T�Ֆu���y�$\/�k�D�ߋ��W��
EZ�����o��ťn�g�������`;~e����*�A_��J-��i	��tU��F}Խ;����P��`��~y�4����*yz��ޟ�����v���R�k]Lb���r{$�2V�y9�3�co���8�[i�R,��ɭW~��_�en�ݓF�Z��=�S��T�&/�lx���Y������&9?�"Dߝ3��c#g׬�1q7&A[Y1x-Tn'���ƶ (�p�����6%� ��cQ:IR�7��n y������V�J)�����X�pSܰ;,������P�����^�0��#p��Y�$�?����)A3�L�heR��<��L�_G�%�@�/�_d��Չ=FONof[�Ҥ��^;��R۞��A��E�Rr��v!Δ����?����:5�ܶc����Q%�Ë�ֵj��Q�M�FQL8.v��F6�2P@�K����y�m�6�7.��p��=��P�k����
=��Y���@4�P��׌�~6����]���XK��	ߞ�r��9��q�$�?Rdr�oH�䚩Y@�2��<i���/��'^�C���w
��˽NR9�g�X=J�XL+\[��L��8����;0��,/)��ԩ��,��^��K�B�����F�M�-,��͉�^P�J�o:�)ׯ1��~':&�@z�FA5H����pI��IA�K�uh1�)�r�]5����~~�(�k#;yC�1��q'�d�8����,�+�h)̲���H�DB���������e�Q�h_�z�����3�+��Ěڮ�	��Bb��)E=ξh��`��b�K=<[3'o!�.��X*�=����&%VC5u8^N���'�O�A�pi3%滜�4�ܒs�]I�mD[�I�p�ňi���E�W��߁N88[�n�ޕ^&�Gϴ�iC2���
����y�vx0>G`r��ɂg���v�zf��c$�+E�~v\t6)[P�,u��S`E_�s�eL����rȊ�=�����j��wA�)nQ;�zm��n~���Z�o3_��2�ໍ�L���PNw�԰���1ҵ�B17K��Ace��JTn��I5�W��n���'���y|}���Ș�Z��6��+-���d�_m?����7����0���I}�Ts���כ�7�X�(�mY���I��@B��ő��H6҅h����a��Q��gX����jV� ����KS�G��hO)�ε���xk�E���B�W��S^�#�eb�)��fQQ�=��i^�Q e�3��,|*T��������7�c�_����]�̃�v)�q�&0�o����D[�`���g3�h�J"�<�WM�.�j`��Xr7N}�I�h^�!�on#z� � w0K������~�S+g���yػ����Qz�,�P�-e�+W��I\��t���ƭ� ��e�% ��u,j@�[�ќ���`�3ʀ�H	�bת�Ҫ��a�26yl���<U/���o�2�Q�����c�*D�:hDk�������R����Mg����;b,�������>�_h��[e�(VR\�<�AP�a���.��?驖��4�����:��*A�R����_u���}�0���L���a[X�
����2�Y�����n�����1z����>��d�4f���k���}P�_�t~TKg7Rw���_��� [pWEq����k:C��I�|�F�v;i��p��JG3�JQ}���l�0�[Lz�+�sHV
T����C�<,\���C��]�|�3�	��ُE��k�	�"���u:�M��I�������9������EK�I�s���#���'��nʄ?�{&-!C�o!�����n�\IG!w�$.,Z8ن��*M�-�����y9=[)�o�"�C��h���'����ʼOUIcf9��6wEv�h�^oІp%P�"0Om�p#! ;X��b3�<PK�ȸHOA`��tBX��d���!a���4���h1*(�l-���U-΢���v���X���Q�ZE�+d�ꏦϲ�<�4�J�����	\<��x({�ic�Z��� �`)5�e��R�\��z�lM���Tn��~��.�r�+���F���>�	6������
��{G(a�?�g$���1|p@:6��B�K�2j��ny'c�}4>UIg10��'�'�^;��ڝ�[�"����C�����r�*��R�s��a�d��$����`n(&����g�R<�0�'����	|z'����m7��={x9l�D,:hj^伞�,Z-,��8�N��7�Ƚzq�n�ʓ_�SV��e<���kzK�q���Z���� Q��y,J��?�=����^w�QLH�JΊ��, �u�b�L�-発.o���ѩ �B�v���0.ڍ�=4.�a��v
ɬj�'�8I�q0omGዒ!W:���0�ˋ��JH�t��c��69*u]ǷU�I�y�jGp�(08�ؑ�%�`'�4��&^ꀋ��z0�G�����F�(=��yB��������"�,8|� ��g��b��k�B_���:��E��V[�G�~�m��*�z&��?�b怇^��y1�xD�IxW�zC�;>��B�b%i�o�*6˦2�d"����?C�
��\F�>�J���9t���7z���^1n�Af�)$�DYXO���*4�	�5w��%V����#1� �S)���qa���=�9a�欌r)�V�m���k�b��9�Jѩ���ɳ������F����wq�l� Ao����޿';=�>��Ե������Z��
�M��ԉ$ʚG3� 7��E���o�ְ�L]A�hz�x��5:�TS���.��$�/J���K�-�	��v�f�C�eZԜ��<d:T	Ȃ�ﲰ]��X������r����	!��I��!�Z>3�<�ǃG_ɔ�-�L��<CI`w�����x��o���5w �?�G\ŎC������_���Ű�r8z|�Kʻ���3NV�ך{Q<b�%���p�Z�/G�Q�O)�|�E[4��%(cԊ�.q�bP0�	 �:2A�k�^?a�&E����7g�v^�|G3W��8�_ѐ�V�mn˖�ޏ�Y0�%�,��j����2YAWq���,���/�(��x@�KA�f�i�y�	d�-��6LD�9� �#�կ�"v!�!g��j�23�h)��mL�[KF����'V�j�!�k�I# _T�O��fq2oD����ښ��4�I��@vw���{F�h�$����^`*�Ǡ�|����W���r0���-}�2���=9�oa���y��O&��W֢�=��L~�߹���!#d�`S��fm��C {J.no�m�6_�����"t��M�0P�>V���������j�FZS��lz�����
.R&%5W?1�ڞ!����D�A0t�S��x��I�Ku�J�z��i��2����zxa��8i��n_��3��Q��]:�o��%�ɘ'�"�Z�z���2Iu,Q�:���M�۸U��2����ъ)6���Zz& �?��\]Ц�$*F��|�a�2�ɈE�K}�P ����[��B�d���ib������21�����A$=�wP��`��'��nE�pSY֗���l�F�E���W�π%��y	�qnv�� ��Ժx�`�[�E|��˗*;6_�URsR�$J��ڃ��>tB]L�6�D�0�P.�躼p�ОRZ�-��v���������P�u�^�<Č?Q��=0�i���--Bx'����!��0�'B����2f=��op=�g[8�on6��iKI�P�|�i@�6D�Yg�0.���L�Je�#�`�:2��G��D�!x+�`E ����Ͻ�c�r��������PG�mOf��C��%;սl��{N��0Ĵ���al/�@��ѭ��׵7wT�0�w���_�9Z�dpb��-@;���=������=�G��f���٪��o���w4b��~��wD��[��Ds��V��.@��vB�Z���/��?��=B �@��3.�[Q�Ƣ5�%$��ϗiN�q���]���؞Id������ѿ��v�l-3�N<!�z�4>�H��3��j�R���>��4��؃��h�;xő�h$��(�x�[���ĈC��	Voq*/j�j����?dO��(H�����s�;Z��3e��\&��Qj��n��`_̣���!���F*����f�\�Һzzٛ���6�FQ��\���W�r��?署��ԧo��#<L��Y�{-
0�t퀒����kL���Jy�9�n���+o��h���E<_�'6
E�z����(�SN��ѳe��k�:r��x�,��)�X�&<[��=�0�<��Ä{�����:���'�
JJh���7WE�Н|C�����6�����>�,���i�W�^��H����?Hj�0KY����5�"�N�1�u�� �*�
��з.&��Tϖ=f�B0�f�@��v����r��RU����:��z?	�e�~����V�{<�[�ܝv@���ƿ�L����պWnӁ�k�o���=��7��jW��9!j�r�<�f��65N����!n�U���t!nI�t{���]`��I�ho_�y�sh��������;su�ѭm�+g�l��
7_MÌ4�o���9��mH����;����}|�gny2ߢ��Ҿg�0D�c�j��ր8�s�r{Ĉ7ɥ�0�+��b<W�tB�5�{���	�@���0Tޢ!ʕ��E��2T��1��h0q�d` ������~�؁�S���ߎJ$X�����6��}.f���t�T"���{ۚ|�)K�i�G�r���$i~s@BR�Y�o�5��������]�K%���>m����ku��>�Hlg�&fLAT��������!?�������nC��+�/�����cᾑ�ݾ�Đ�x�>q�ڿI'�H$���zu6�X����"h(�0J\�	��R�D��-m�o���#�g��d��ʂ�{�g�� ��4���(jGٙ�IdA�$)� �&"����tk���"If0�>c��]r�LZ�#��5�E����?�"��Kɀ�.Ѩ�t2�a������D6 ��9r��l�8�5GSE�����%�n�L]�iE��6�U�"9��}0�7�ߢ��W�C����I�Π�����J:�D� �]=�p�/�8@DrL�b��9u��ɲ��(�z��ue�'�@�܉����d"�;��ڒ�ɝ�Ճ;O�	{�^Ny2f4@������\�������C� �
��B���6i��V�.H-��^��0� ��Y˪��3Ԡ��<��u��,"h�T�\������XG�I���4eϑ��0�	��G?~(�� 8Ԉ�0��\r9 Q��])����ٗ���[�D�{k����m�m���i3��C��T�����x�o���:��_���4d2#�h�#�������DB��y�vj{�q���$o��?��'�6�!6H�bv�=��V�BY���D�S�"���-��i��T	�D@̌�0!~E7��}��4�O	1	h'�%@�4$z��� �R�����;�˾�?��VEA�B����1f�ǷΌvRöz�C|����a�Ys��+����@tf�>u��o�xy�3�F����2�ʚ��~,zX,��ץ���-2�5��jP��,�D�" E�oaE̜f����yMCV�Vʁ_+���0U��Q�i�%k���������]��X�_��Im�X��{�'7l�p&�S�q�h
�^�>�@���~J���5�ۻ�+W��}��"���q�qo�HQ*�����Q���e�S�L���>�{Ȗ!G�`<�ۑd��{X5��*�2�e�����Xj����i�T&���@}�ID�Q��{b���Wv*t�ҏz�-1�r�Y�[����?���+��{<��S�7��a?7S.� �]�:������V�=C�a�#�"��K�dZV&_�J����-W#�+qA��w�a�4p�n(n}K{�����oQO{BrƐ9s0nt�xƔ���A���H�YS�`�d�%�lH[�ݨ���?1�f��X4i�=:�k�#M� U>���q�����Њ�+E�ل<!Z;�4�/c�-��[�x\k-�}^���E�r~�99���D�d��"�=e���dD�Х/@>��?n6Y{� ã����Z7�`v��Q�ˌ��s�-��k��<U+sIJQ��Ǽ�a���:��F��Ά�M-5��o�Jy�53�
=�8n\L��؀�X��ڏ�ݓ�7E9O��]�X�
�-�k�%ˊ�&��w�ut�j���_ո�O��h u�9{͂,8�k�׌Bs��0�¸�>���+�w*\���O>�����3��}�1-���֪讙�y_/��O���f`2|�pN�>D8ėx�	;����췓����ץp�>�<�YiZ�v��W�g70��|y��}&Z
�Sْ�O�u�JI�4��QN�S�b�8�xL��x�Y�,��sê%�mN�RGq�y�6>�Լ쌂�����;*{���z��g.8hZ�IU�D'!��l���#��|���n��z��=�\Ė{±�a�Z�j3����$&��=�K�{2�01��!��,�E�q�zd)�HЦ��hFR�yY���l$ �{Ifv�=�䖸�WP�4��i	ɡ�C�h���ܸ)Ƅ6�_��fC%��?���Ѻ��Ų x�*L�f�a��o�*�!���+��ˊ��߹Gn�����@�"��\s"���t�W{�7*�O����Q�\���pl4y
�r�lȴz�K67F�03�t����Gs
|��=�픞��Љ^�o��g�l���v4Dlg?��/�'f�����ULI�2�ƒb�,V{���'B*>:�v�.�e�xF�`1�S��n�q��)�!����Y9�$\!��t�/GB�� F�pf���d��Ȕ��՜�p,��^�URn�yLy�_���M� D��~�ŵ}��e3	������)���kw�K:|��H���[$s0��q��i���Ժ,8<~�:7w��6$�93��vp�ǯ���C��Y�e\-�<���%�f)Q�6�x\�����/ ��\ML:SJ�2���Xe��!V%B�C�"	<��2� b�Aܑ-�W�AHR��O��Cg���I�7P�uȒ?�ȃ�Do�7�:�ǆ���:7��">�7"��\o8��t��F�J�$O�J��/Q��2]��>)����+���ǌl�?�?hIj$��֧U����Yj,�N����?k��H�n�#Z�y�GJ��"W1F�e� �Z>޻d�k-술��@����?>&���L[V�ТR��33�-��Fe�.��܉��j|\�� ��g��#�h��_��=̻����)wB�6#a+[0�窉���H"�^���!AƬ�o�_?uVW�Y]�[u�o-����ڼ���"���뭘���^[6[����O�ۥ��(�_b�M從R̫Y���?f,�LC�:���g�?�\ťq�F�2|su������B�w��ז�za2g{�b� i�n|p�����SWm�*��?p��J�l9�^��� ��N2�Ȭ��/;ǰ��g���O��Q��x�rԖ��B@I��>8�&��ueb!�`� ���;k��\T���� ��<�,��"}v�#�zotje:Q=h���(�(�1a���K�a,������������U:�%�oY�y>g��אk#�q�
����bTp�V�
#l�1��:��5��#��|�偓���h�2��F�)�ڙ���L8ͨtR��,�5���@^kG��F2���ٺ�I�S�D���: J8	���O��)�pAB��kl��}��v)��xi�s�[D{�v��0Q�L���S4w��\]�@m�����v��xh�������9��Jfx���V�w�T��QI�'���|9�<-�-���\0y��x3�S�*�U�����MRn�Y���kj|��@(�Gܩ�!ޗC��k�8���i��%���J�}2Y\�c�R�elEǾ��$�g;�l��;p���Ο77������.9Ꞵ`V�q(]�튈�D��G�U3���v�����A8�ƽ����ם�)��O�Ǉ����`�9��
lAo~��R�I*~G����[���I�m�6�=�\���#  ��I��3,�F]�7N�����\*R�����݆�l�&�[�bG��#7;_�R�R�y�Q����/}���rn{I��-lq�ҭY�#du˱7��Z�Y�X���:w�1*d���v"��3�Hɷ�)��H�B�|3 �� ��v0Lh����S�d$�,S-Ӕ��t����3=�&���AWY	Rb	�j�W�#;/4����"��q�<�l�ܩǥa�M��_�����V��Ҍ���k�	�i}��� đ Y�ݲ6�h`����c0ϼ�*=J �^��U��@��&Cf���/��*����%�8.�&���Gx�&�t
=�����Q�x�m���R��"$۾O�)���^n��#�� F�M�r�Bd�:�2Kk'y��Mb��ҙAhH��]�ID��#7f�S�����V�rhG��_L��s�D?hL��L1Y.��X^i.���z��]�k�{x�hB _���Ar�v0���H�
4�B�Rz�D��0f��~���uZf�m�$.�ܥ�����q��}Ј��ͮ�:ua�� ɍ~��G�[岑e�ˊ�a�R�����������Y4#%=�8������q�Ь=kG�n��K¥g�z���z�B-Āը�^���}_�)L�����i̸�� L�TU���f#��>���(,a~�ke�N�vB<�(��i|m.N���݈<O�:e�c�$�wɼ9�N�{&>�g�?)�=�6�p��W���[���������̾��/��POv<�Y��]��'��y��;�p$�e���aq%���]o�Ϳ�����C�غ�nHG���ۏt���X��cΨ�h��b&�M[#��	2R���֛^S�L݆5�R�b�S��t�z<��m�y��v[F?����si����G�6���yL�R
h��f�"��%�ҵ��x}4��%�8�)��`��d�O�&��t���|"�R`w�ezC����}���9�^�u�TI8_~WB0�� f�8G�75��	����\�.��D
>��%����{��9S*�D1 X����ȐI�$W:��o�{Žw(++�]��Ј%�C`�x�����j^6�"�z�i������"z��l%@�ސ�Kb�U4FACh�Tt�����_rg��B��+�rl)f�ﳶ�ڔ�H��`w��Ft��m�F��9RV	bx�Њ�,1�@�UPV�y(C��V������(Um���H�v���8�R�W	�ix����14�>)�	 3[ �1Y�zy3��0�R���,� ��F/���$��0�?��|k����'T���b��;��8e�_�����7�4��u9�<?��lH.yWR2�q�1 �9Z�3�u�Ȳ08��3�۫1'�q�Usu�_��"�k$����S�ޜ���Q�wG�L�X��4oU'/&ThV�/>v84� �q|� ߡ\�4זH�1</{�FA)t��wQvC�:�G0+R��D#K��W�����X�J8y7cj#`�U+*BM�M~�h��Tab � ����)G^5�4��� ��5�Jrm�9L�Ttm儖��9\$)��B���J�����d��J.@\8�v����wEY���;3m�ϡI��*�����Wk;���0�5�;�e��'�m!�x�:>0!o���+���h�Oha�ِb2(!�Ł��x��[z?Zum���@|ػ��e�_�݌F'���S�t���V�/9?�Uq�2���W#��.eg��h:�c[��כB�Q�!BM�`t�l1:�֞g|
�Ԉf���Ⱦ�;�mʾ^^J�Q��a>s��?;g�5�Z�M.�o&?K��vrA��}t/�������(�_W����S��Z����(77�@7��{"I=S[�Z4�	���[���k��S=9�-z���}۶���^t7�V�vD�R>"������P��s����[^� ��n�e�`��	P=�
��:���Ò�m7s�'�_�&�#��	X�T�#�ԧz��� �����d�T'�߽�i�����8=��1������E#ur�7?�����l���ui:t�&>����CP:5����Lә�j�o��ʃ���\��{��r��^}4��o�2� �Sa���B�����̷+�N�b�୉���'/�����0aX�F���j�[J��57 ��(\^����0ϋ3���P��J[����1j��AM3��:����t Z�����U_�4����g�+a�	L0�ϵP���,Y9��X/�m�'i����9�h��k�ͽ1z��n0��Z����f�<��
<P	��N���$��D�_5F�(ʃ:K�f�3�$$KB�Z�H�?T~���k2zӗ*.������do�f���VZ� $�CR|��C�9��=E�c�p��Īp�}���=Ձ��F���S%��׌-�+�,��7r{k��.fI;�i�援�b��Ss0��9h��_xim�&�bo��#%�4+Ǽj1-�p��9G*���vK6�ͼ\2)�:�A��t-�<������l�c"�W	*���C U����i�_�֞.�� D�]�����3�R�uK"^F��@�sy�����6��?����8���v��Ǘ�=]�#���)Ul�[G��_;w��d���7�ZeAD^s,��D��L#@�ǋG����������c|-br�����ͷ�ڿכ�l�T��uk��b������m�L�3��H�+s�>T��W���F�ԵA`c�HKw�&V�!����5 �Z�;�^2U�},�z�S
b���C���;�
��.DʙU繻T�U��r�\�G�%�V�ڵ���I�a��'��@Ѿއ��*(\�8�H}��A$�E*v��񽸪��
��7�:M����Y�И���3v��\�f�}/�DZc�ʊ~X`NE��w=�]<`tÑ��>=�"�k���	3ċ��/YV�MA�_�ޙ�A(Q	*�5��`J,�n9��W��p�n�Z��wQ��8U����_1#M�6 *��q��E1mv%�:Hh�ڄ쌶_|0V�#B�7wz��8�����ހXQ �de��n����W�߫-�i��� ��uo��GUaOs��������J���)%���Pyu�]���s%�\��L��v"���C�W�p�20� �W�H:����;��:�c��3�m^�u��E<&6Sxܢw�Z�����Z�����q��I�`�fV����%��ԓ�K)�LI9���Rm��!�SD�;ɄwyZ�wm	����
���=�q�+�����Lm��`��Hb<�}�}������+�z�љ�0/��C &���m�_����gb�{�mЗ�ki+^�}R��'�и5�p=u�{$�X倽�	P0y�m�����ܨ#�+�ގtN����滆�+��isaa��F|��0��!#�6�VdТ�x���,Un��38�pMż.���ź;w���?��j�+��b��t<Ϣb�>��� 7&�S�i,�+6��O4�1��1��`��Vt�78�C�-Уz�c����i�H�r���D�;�)rs��&l�Wa<>�I�,�t��t.�9����'�f#!bBq{�==��ߣ�`3��Y5_X�i!�8A xp�s�XI�����2ZH�S�7��l�)�~`U� ��L�D������|�%�S%���#��o⎚p���h���E���\<�����g����\������o��`c~h$�y� W+6z'���$rBĎӮ�T�n{��;~axjX6���3����޷�Y,8�&F@ߥ��Y�!`���5��A��
$����p�|Z�Ƽ���W۹W>U�Ms	��MƝ�e	q�˖��5�i��Xٷ�U�)�C�������.���[m9[B�N��z3�s�8gג�0E��O��
F�'�q�|Əy|�94Y2�D����I+v�����(5�E<�lԼē�3<�F�p��e9����K�˓Q��`B�#�� ��q�������6�P�m��G�M��1
 Ƭ���v[՜��q�3�:O+�?a���14�<F���r"?���~,��C�2Nz�j��ȳ���!�ov��RQY=���1���	��3"�j㜚"2�K�h��̈́M��T�u�~H.r��/�Y����h��Ed`�v�s}=�Z>N�X�{�S�o�����	��(�o����i�R�9K}��#��s��z�pL#t�r@�m��hz���] T�|�Vs��M�R�,-?��˶�zc�+\#f�?d�|�%|ޅ�픾��<��UȖ�L�P[H�+�������k�BS�Ӱ�51a�!d�5�/�U߂��Ł�z1�Aה��M�$z;6��;R.��M�I����jѽ��WW�u��_P�[�ӒƐ�mzq���>L>�
*�a�؊�S���)	����s����u��44�({�P���Dv���&�7��_�Y�������E�p��h���?2��zZ��[�ɕ{H�Gf�"WMU�Ρ2�7���f����{�/<ʹiҔr]?���YS�����K�'��w�d޼�t�^Y'���k2�x��_Q�_� �i�H2�^T	I�sHJ3�;��4�OiY^N'�[`�K�������^����GI"�4t�s��W�X$V��&�'�'d�Mu�MQU���;9�oތ��w@�3��x��\���]��;�헟>�4�#���ŏ\���.,ɢ
>�z������W(y��4��u^(JI{��'�#X0pp��
k(SX/��P[4{���
�����+g�U;�6����}xm�.u�0�a̡A_���m�����x�����N��V'�M�X����4�j&L)&��OW7��Ý�S��Q�"@$���IԢ�mo�C�6���fD�`�~E��J�:FX\�@�O�(�g�=V=��oW����j�xZ^G~-��f��1+@B��X�?që�����
���?�`p�F���tk��͆#J�˼R� o�Kix�DZ���K
��_t+Z�(�)[�--�������Q�#�����"�RC0��OL�Z[��$3Lh~wm�`ﳋ������,~���jCݥ�9��KN���䞢ً��vA��o#�Az��Z�`�B�*FZɵ��0���~�8��S�!�jy���g��0�U��Y°LMiM@_XH݌�~7��{���O	����at��fJ���I>�El:MW��9�'����}��o�Q Iq>2@���
Fh���2=�O=V�uO���=cI�����?� ���W�#�I�����(V�?sJq �G�o.�B�ܾX��1k�tX�j�{���Y�"�Y���_'�.}�Tq8y�D���yA�ln�8�r:u �Q�ۥ��A��CV�pa�#�V%v�ub|l�'�y�Z�nS�3��%	
��gͣ�Ѧ�N�����ʏ�@��&-2m�8A�U�.�7��*���hʢ��i��ʥ�TN���a��g�>�_�h�5��kq������Å��n�-�;�g�<�꾱!�N�$(��ƕHkGTp�t�S�H�i�[���Alj�z��_-2�A�)E�~�S��:��	�0\}��b��q���"-���ᾌ���'V=����k��
x�WI��y��?�_�g���:�Rp3��AY���Iӥ]pg׿�F ���B�d�j�"����N�e�5}�?� K�/�۾�̍U7ۨ���9�R��mK�`p�=-�|Y���-�w%�u����\K�Z�>Fcs޷�4_�ƬV5�߷)M�����^�k�L��3�H���n��Ȑ��	+�a��/j�|�dN�f!�|����ϛ�V������<���d-��T���#����j�19�LI/���.�����';�����&,��ؚ��g!�s��]d��M�����V��v���PW��:D�U��Qؓ���y$$
�5�$(^Q|v7y7'L�]P���)�'\�H�,�z/*��|��^��8}qwxI%2y�!��$j��b��o��	)�D�R{e�w5Z3NI�d\��@'�4�!��"��/���e�'��5�,����h�R�o1��$*!>��n��o>����|�6���+a����(X�!9��E��H�b@-3�Q�������hB[� Ku���������ǕyB�1�U�$�o;�qF�"Z�"�(�F�s��Ƞ���{�6�3�O�-ʟ�w
3��!��:�$1D4��б&�%���H�m�"�~�S��o��-*e!���(t��<1��W��W�����f[w��_!�h��:cYhW��`����\���S9�h�-/��B��Q]�֤P&s���MS+l�y��[��C�^��@����n�ćǔ=�|�U@�v��>��09��e)pJ��bb7~x���Y�N���:����_<�/��Br�g�������Y{5CX�ץ�M���7�btN�f:�m�r��1����,��D^�ĜQIiN�;b�����<���x�%Z����@��`-u�*s�����F�i�[��\`-�^*@j��Eɲ���ż%�$���s�I��<J'�{��菜MU+�'�l���T�����^$�@�R${����y��Ǿ��!ӑK1q����E�E:�a}#SyF)���3�2���R���C�za��p8�g�E8F�W}��/!�&��{��	���{H	��/@��VT�.{�y��Mw������p��S!����I����l�.�FU���2,��ڿ��xv�H
��@0���7aˆg��Y{-v/�i���u.ۜS�D�L�r��,E���;g?��Q��ڃy�0,S;ʩ�K{�L�Xx��亇���A��=�l�%��.���!v��Z�ܲ�*ч)[|� s����TB��Z����Ƶ�� |Y��|�
t��e�C�5���u����m6D�M,DqE����cj�h�u/m=��c�y�[t��Բp�2.��$j�=X#��q�Ƕ��Vjj"Y����B:p���_i�n	Ό8e (��_�����qh�k���(Z6��j����ڝ-#YC=C�HE��	����=��9`�U�u�{!��lwqW�5��e2��7��Ä=�1��Js�
�
P`�S4c�+�t_J6��i�]n��g�\��2r�CJqRtp�'��kcSd�߭H����dC'Ŝ[5�Z�1&�P P��"����#�s�>����0�t��L�Y�=�rK꫕��HB|0���?��?57��Y>3�䀖&/]���F7�񦯗������`}�ۚ�\�a&���dV����8k2o_��PAw_�JJ~�+Z��sh��h������DIw�cڤ�4w��PC=�$lco���բ��M	LHN4zs��dL��h�9 ��ʗ��D�&j �����W�/�K��'x���!rJ���3*GM`�|�ۯ�� �jD¿�wά 4�R�.�<K-^�=��F����D-a�4�T�N����õS�P@)
Hg���@Vka��C����A�\f,Y�͑�_~�|6פ^Y��'���SN���y�(�����ۦ1=�>���z���ֽNk6�^�R����#D��d�Q����S�- �0���O��D���_]^3=Nyy��t�tL�]���E�0���I�f��.�|���z��Y������"�s�7·�p�z/��[��gC�
E�o��^�aU�ot�q��Efě�J�YK_�o�bXz���
ad*�t���%w5�XA�WJ��:����sL����W4���\�ge7�H��O��J��2`-�2�D-U�$�mw l��J9U���K�g���+2�TsL�������ߌZ�.�Ϲ�m����6�����*q�kW2nC����B�^s�o�k�&�O�d8>E�)ػn~�	N�� ���W>�m�uF6|�oo�;yu��ȓ�\i�I��J�2��yx>:>���-\�]6��Tn�����O9����L�!�ͣю{����[�������#�j����h��<�h��R�iSn��މm��<3\��;D���@B&�yz+�JQ��<I˭X�Y�=�-��BUzL@� �aM�q��p����f�&�I��>K3A�p,�N9H��5�&���||�%5e)81,;6�N�c}B�O�;�f�x15i�;D:GЍG�_�)���t�u�=
��.X�����w��S�k~> ��o'�����F?.k`T��!W@���,�ͼ���>L°�2'�U�Ѱ72��e ��u���3�t����[=��$1O&+�t'���9ÏS�����C�e�����h�ӫ4���$��?y)��s-=]#؃����h�A���X�g8��^]�j��Rat��b�dV��e�m�m{�"ց���t��:/y��.f*]�tp�I������HE/Kd�8��P{4��	X<��NW�lMU������m��n��=����v�r��
��r�\	���v�p"�l�����2��Z:�@�-N��n�X���3y�߬*nc=����k�r��\jO���:J�}f~ڢ�ʃPX�~��F�db�K�J\TS�v�Z�,��������ܵ�b���g4{O�9��< +�_6�6��^N�r` �^c���qp�+�mG�T��ʸ&;����\wz�P:�f5|���M���g�������o^�#lt�p�q�Y�I�+��m���F$^0l�@�;L��l5�,W�b�M�{��S!C��];��@�B^W�4��^���UޭD>�`��'��?=��h�[�l�;J��e�G�U����Hs��C��#�Urb�fV�:��&h/��L`�7gn�h[~�%��T��2'��t��s�Ƚ��L ��>�:�B6�8�7��e�c*K���ވ�*V�1%��XZF�q�0ȓ<�Ό�%��ۿ���\�a��������KPZ����a�OY����K�D��,o�����^?͗>d��Kƨ"���/'B->��)�/O};����#�Fw1@�W�9�h�>��0nj��A����� `��5���[�k.��Zm�"0�nV��������0l%p�`ǝ��;a�oNk�"]
"G�B�cf���~�N�⚛<�_îQ��V�[�����x���&�!1�q �DsMҳ���0�|�Wq�$�Q6[o�93��|�]Z�R�����c=����Ok�]�8cD��F �")8�>�|i8Q�'Z9��|�N���k<����p���{�zו"#���8|��Z{�zľ}�vXQ�Jb�� N�Y
x��g���iz�����|w��}�sR��o>w�8�I�'GM�x�VvP�6��6�Gg�h��{�5�n��._/W~\q��ӴRr2���9�7��X�����a�
�݋�(%�eW��z�]�<ϗ�Kg��{�K�y�p^������EL`�:����wV���0��?�C�<>=�4*�I�B�u�#b%P������(Y������L��,�y�Y�6���E�GݯdJ���YW˕1�G-��y����1w��[!$KO�2�˦XW�#�}0�������w�2���򬪥�W�Sš�����q�ӿ�����:�g�?^p�0��I���F���ő�j$"EE8�N�COX��ǌ�,E�����Y��"'� �$�W��0��@"*C�&���k�9�/eR1��N��P0���M$L �Yٹn�F��b/�N�{c��o��D��*cO[�q�Y ���U�S�`�j\�Pb���R���3�X��8`�h
��Ts-�Ot�L���k�����?��f�|�)�|# 1������)w΃=��m�,�o&��Q�Y�΃��s��~��{k �oـ����H(�Z>�'Ij�{�|kҵ����^9�������8z�K���.!�n7�ljB0����u�7D���X-�K��=^���3A�����Hꖚ�[I������$R5F��|`����h�b�{�S�-W��u�(�R�پ���(��`�fM'1&Aϊ	�� �-�ZI`)�Am���Ī�'? �*�q-��`jr�ҋsB%S��O��x]��G8���nJ� ���\ӼZI�EE��mYG�{D��QI/=�˛����b�3Q�!6��Wlw�i�� ��?ë.!�R\H�ɒ0`��<O����|��mw�������ϋ�r2�����N8����w`�,9M�T�˲��EmC!*�r4`�x4\��cr��Ư�������/��Z~i|ª�G��ȑ��.d�U�WB�����o���x	��c�I*!�*�Q�caXz˗�������jW7ܠ���%�� �|�]��Z�c�=$%�'��nץ�5�}�B��Q�[��m:�-�ӜG�djT�fFTX��%/��{��O*|�w���@�>���Í�Q���{>v���h�i��L�;:U��X,����;���'s�s�! З�%���ޮ�7a!,JL�W�Pa�a��P�sp��U:y2]b�q�Y��Đ���"@���L�|�ٱ�x���K ���Q�e<�+B��+W�WZη�a�`�0���6ptj`�U{��a�����n�S�PV�4��8PŶ��YO��#KH��=�V�����1n͆[jk��b
����r=�TfdL&*�t�d�!B.lJԏ3�(*�Y���$���ד��~w�7M�4^
�Q�p������Y��\�|GQ�"�D����:īk�����ƙ(�au ��,����wt�F\:AN0�#x|N@آ _X��kڌ�s	���8��ЊT`ٲb��1d�wͤ��9e{~tT����ւ������u=E8��G�쳠�Y����~q~��%wJ������ٛ\���K%����y��u5HS�o�ѷG`�� ԥ&���=����X@����'�O-�9��� �]3ۻJd��Sd��`/x*�m�/�/Iɜ����3���9����W̻�rÏ8��:Ҥ$�q��h{ܓX�4վ<��ܭ �nZ�FV%���ŋ��Κ'v��,˜���"�s6}�^�!y��{�A/d��C�^%V �P���|��F����悼�:�Y3M�dNP$n�W��J��yȵ��*�|X«��9����97��鐪/�;��20��˚[�S
��*�k�j@�ѩ4w��44v?��&��b��K��IȦt�ǆ�����Q�"kG[%`�(SW�}3��W���4 ��y(����Ǳ`�I���~�7�y6r�B��88�TM�C�ō5�v�d��{[�.w�1�"&��2W|��&v��@d��@����1�AZ�m�p�w�FT�	.�^�jp3��K���y' ��k��Q�$G���d����f�nF���%�6w�'zY�#	2�(�?�u:�Z���M�u�t�φ����>�㸧0�/p�3�X�[�31� �<Zg���Q�ꟶ'i9 ��#��Nh_%&X^��
����C"��H������l�S���ШW��l�M�K��dBU�8q�������H:�^0�2���#+DֺL�kF�d�zN_J�����l��- �+�gU�����`t�=[����.����k�{��V�7��QpR��d�%VFc�-:�����n�//@������_��wK�XcէG_#A�Ӵ���Yh6�f�'LǇ�L�X��p����j���A($��ށ�
�h���o�`f��A�r�h�>����M�cGo9��L�H��N���!G���+K eB �V����Z��d�83 ��۹bM�s���3|ۀ�Qb!ʹH���e��ߑp���QH�)��t?g��(���xU/j����ֆ���Y���E�w�61�E�_l+o�*2tr&Lڼ�R�~�:�ņ{&�;�l�R�m����_�bhqD ;��=��9����#n^��f�^hc��>�kT���I"`5C �+�|W���Bi���_  (�CDd*A��a��Akh�[��:ÁE7h�[Ȕa�- [�.��_�!s+գM./�p�TV�e�����*�1^q[��f�W 1�+e�b;L����o���ʈ̔�4։�Jk� q���i�V��A�n���'���e�t�B�4�1Ǩ��0T��G#^[�!�)���J�dqn>C�X�c	l���R�n/�Ղ���+�sյW�R�AIb4b���(&�Ċ�	�s�#�2}�b��L�Խ��G揤���&�o�rn˱E :0���s����q"�M�e��H�m=�2���_X���凮z�"�MP�i�ؐ������1�q�.����RI?C�g�8ǟ|Q$�w]`�D�f+�ƒ�z��3:�i'��Av������t�\є���0�*��x�ܲ}ì� J�����sy�Zr8�/�ش�R�>ڏͺO�$��hȶ?>l�]��n���e��F��jW[Bޔ��3�����~�����ټ�<~H,��m8���'6rI�@�a;�ֱi �����?�e\ܺʸ~�!~o��h-�&�1u�l0{�J1l��vā�S<��C��>����=����tV��Q��|� >�NeVxK�Wk�.��7�_�- 2Jbi($��G����}�.���!��� ��Z`���4�Aphm>ndc�ĸ �Ҁ��5�^��8Z�v�G��ՁU�s��X�>���)^1~�(����J-�t���ه<�{��	�D����}�~�ù��ܳ7C���4^ATD��P{�A�w�e��C���/�ǚ�?���|�{N��2zZ$�!~��_vGI�5����E�[@[�����Q`A�<ʋ7�A�
rPģ���p OEZd�]j��e�	|�fT�6�C*�1�y��5�/4�l���5�,q�`��4 ��V$Nh��=��8,�ϧ��؅	�A�1��}<�|+���`�E��҂$�����'�@fi=���1���"��)���ҵM�3���O�(Y#R�Ձh�h�t]B�Ʒ��Om�������n|5}s\��B������8J�S�:�l��=#���_GPn:CJ]@�$k�?�d����F��G��Zo0��b�i�C5`�<T���Z��/~�C��>QP�o9�%�^�T"�܈*.�4����#h!��x����
G���_vJTvY+��+Y��yܜR<̙��CE� ֮ ɷ� <��bl�[d||9bs��d�I�-�F`���Cͺ�e�>�8�%'_��QQ��d1�@��� �o60���ط`��t#�6��5$�
׭M5)�I�R녇�{�;��و�W���f��vl�e���8�m%ʞ|#h��V�aX�$��������w�������A�"I6�Do���/��N��_^$|�e���H<�3v�.r�O�@<n�uf���s��b�?)��g�b/��yH�e�����y�r���%�	��v.<��⫁M�(Oy����[�b����Yρ?��`N�VE���t��x>�fpK��*8|�D-qD�<F�f�o.U�DVظw^�p#����˒�4���1�5�tj�I�r�_/]�����?�E&�; ��_V�����U����@�2ew�v����5���r|�
1�_KED�>yL�Q,]��َޕ:l�Aƺ�"r�0��Q %a�c���c S6��2�3��V������K�~5(��CE	v	�j�ߟ�\�i�.�j�Dm�g���"�P�t:�՟iE#�Ω��1櫹�VIg!iN�5���a�M����;b4j	;Z��e
(��MX��`%;����B�����e!\K�&}}ğ�BPO�usr�����-$�Z�b��Ğ/y�(��[C�R�U"��
�8��8�3�>5N�YBɃA��`��5�)����*��쬬s�	������ʚ����0^�X.
Z����~|Y�hL������\bE����_@tP�s�xs�h�b9�#u�3����i��^��7w;�i6���;׌���>\]C<�I�cv�v˙����cR�>D|��I�s�J(Q��+Z.������%��D/|z<� �yh=���L'|> ��I)�w���z@�$6F��Q$ �s������5^����u�5��a�-
Uo����1�j�����Ds���S�B�ä� �����2tRkDQ��l�֦o���Zg�В��u��Q��J���.p
�ٗ:�G8V�~ =5W u�$2�h��27�|&(X)�]3�=� ���w3`ʯ���j(/��f��WҮ��*̈́0�_y��b
���\��԰�R[fq�>��ZEз�khEKɓ��|~���Q�(�巊i_��8�0�\VQۚp]ɜ\����&�
�1ԕ�i�bj2�F�\k'�Z�LZ�H䭨��Tq�a0-�I����X�zH�S�X��ݐ�q*3�/^���&���%0kY�>HV�Z� �{sQqz5���g��[��%.�r!�'��4�	�k�%e�^�9zM�/��p#�4JEE�1A��߿SMo7V�a�;��3ȇWD>`Hu�%$�.YU��7rA��Ϳq�	t����ƫ	���f��J���;���`��T��b�����w�^5K�&�I��uޞ�8��<�/�a�YK��+Ĉ˘��{wӈ�K*
��f�̰Z!�����юcY��9�؈�72.5�^跢 �ܭ|i�Xzv�J������$���6���${ͳ�S��?�R�(��Ug��ڨqe8��������]+��w����a�4m�ȜWox��d����(���C4���;��g�'C a��<&�@ Z�ud�J)�>v�.��]`�	�l��ڳ��A��2N���``�,ֶ�a����?��7���������H�7ő��Uu��y-�Fɻt��\O�6V�m��7ҵw%�����j���v1��R�^�&�`���f�#!�ϻ�D�b-�5��Ǩ���2F�Z֞�(1.��D{�G'��^Xcc<���&�W���>�������QTs�k��yP���f-�[��*�J���;A�(�uv?�ճa�X�0�S�*�>�\覕�,���Sz �: \:���vĚ�^a�T�Dhfz�R��|q9?���ٷ0�5ď20-/��ss2oc���+�O��
���8�4� o�����{QB�>1P�=\�E\R�I?�
=X���_O���ܖ3]���]�(��Z�7O��a�_��I(7�g<���sLف��q�n�7$L}�{�$��K<$���	{#�c���%������;�b8�8�~ll�:�_s��η�#���6�ꌮ���u2U9KQ��K-���M����� 3i��� �0�2�AB�-�x0���^Nk�������Ya2��{��3�d7�ф�m8i�I@�fĄ�Wo���L&�V }8�n%� Wl$C�ѲFv���v��C��֍��1�!��Ͳ���-{H�R.$|��g�ܷ� ���)��շR��j����|ѹ�F�-��o�X�����S"V�.��r�1!�� U0۾��i2l��~Ή���4�w#�=L��z�K5�Fz׍R!������L��A&j�je~q�Sh��a�	�����TX%�x2��$��!�s���}��cES��,v[je��j|�>8�1���wb�?�+`	�r�+��c�gyb�#�Då�������R\�}�k[��њ�:�yZ_���`��t���f9g�=��&'��I$�u?� �G`��B�r{B�ՠL�}͔����k@�F�S�{���w�%f�� �^u�>�lZh�0Fb�
vF*�2~��$�U��o����^U�K���$v�H���ۆyK�7p�\��Me(�s���j!� c
�b|�z��)��Jt�$��m8s�I+$a4ߨ�pXe��0�Q��<T}�~ q�uG�D��Fܒ<Cv�Ε����dR<����t_t=I��ߣ�p��Tn/1n,q*Ӑ�UޘϓL����^�O������5�G�����9��P���-4h+�S��*U�F�G����6��>d�ر3���!jv�5��w�L:�����h�@�͟aAɮ�Y�RŇA�|�}*��tBu�8�%
m��Q�ǌ���_)p&��+��|�yn��w35���dً�p�o��D�3��_�O$ˉ��ps�3'`�.��� "�gD��/��z�f���I�~(~q�-���a��/n�u�@�OX�w��E��#��`Y�����{�g��segu*
C������4"��W�=�R��h�5r� !�>���z[�w���[��L��Ц�*x���ά�;�r���q�n�,���o�^)p�WU���Eg�T�Z�A'�=���k8�l�>Ϭ�d����\��\�笝�4@�X1�w�5$��'��'e9�ӻ	 ]BvȹMI��bv�ꠞ٘�4���PC=C^F�Zʄ�ݪ-��y�*�a���������j3��Fg�=wԈ�W��7�J6`|�v����N��E�1e���n����粆�A�����9s�![����{�\z���}c��H2 ��� ���4��&׿�؜*�nwAE(��w���.��Kb����j��v#�����|k'�) i�6���t�r)�y�y+�~��
����h��ёTF��]��[���������ɓ�VI�G�������oI�������|iӼ&��+�͔ �����,��W� I�.��ib>!␋����C��3���Fty.lk�e�i4�#E
���Ӄu��rD�w|��[^���&X���5x�S@x�ߧΗ�5�A�yc�!"�C��I1]�s�y�G �2��4nG�͂gY�>���0�Z�b
�؛��c�y�*�|����X�x����f\ ���WL��n0�m���@�<WX}�<5�<4ş1�}$7#�8�"'�CŦ�h�DF�����BO$�پ�[�k�讧�����YX ���t>�>(g�L�-'j�~�b��]�1���Q�?em`��]�lsI�yz?�ȟp��G«�o�q��K�ܷ�WVo!.B��M��e�]�V�I�^�����2'9rJ� �1�4QX��ܐwE���nj5K�oԝ��O��L"���2��+�@����m�n�u��:<�(�G�=�� j"4F�nW߈�>'ʔc'9z�o���T�+㭾�����X�nP��5s=aGi3�Y��k͙�BO�^�T>�c���G��3-|��I��m���06�c{#�-�,�ŇK������=bQE��`b@�ČTk��Pn�Ř�1k[W{�*%i��Z���G"'6g�jYC_<��E�X� ߨ���1�t��7�D���v\ �R�!��l~��@�{��.N�lZp�U���b4z��:T�r9i5��e�)�dzx�k�xX�__��R�:��SN��Ȱ�y��͓^]-M���Gd�� �<m�Ws������aS6!Q��T�[����c�Y@�*/x7=o1n�S�ߐ	��_ɔ0��� �oD�$-h��mń7�Ĭ�h�WT�༊��Ȍ&8u�D�5��s~����aᕓ+�L��*W���/�N�?�g��H�P�Fg�g���+|"H�^��l�wm�X�?�P��bM0�� �S	�z�X!���#�a��\t����D�#�kr��`�ɀ�0<��D*�4��O�XB/���:�r�3/����ö���0qe�*ӥf��Ʉ&�Qai��4������l	�wl��FDB�Sg�he����L�7�� �1Y<EKpz Ό���\=5c�̄�XQ�X݀�K��������`u��+½qm���myM�"䦜�_)����à+�ߤ�I.�1j�f:&��.��&k��������h��|��] ]�B0h����2�]���J�ȹ��!8�pj#>�T������wq��ܘ_&��xC��j��u���ܼ����,x).�-�-�Q�8��ư�{sT� t׉�*�R<(����<,�")k���HY��b!c��|B` M��T��I���s8-V����������D̛�A��4Xz��/a�e,)����(�$��ݓt��/"����/�N��֤�Ş��/���C5I�����R�{��J/�f��],I$J��%>P�t�� ����oy��F����j�qs��oho[��
[���R.#+�v�����R<e:�:=�ZN�y�!J�h[ޒG��y+'��]�+��*�jL}�"~jtǜ.�b&��<Z$�bf����<b�:ѧ���y0�;mQ�n���0�"���������l�:��<5����Gz=�;98�q��D�:�E�_?
���a�
��땃�mH�٨�
�AoP������.e䯣�k�BS.���U&p�5N��ߣ���*X����S�=��a�0P�^i�����*KH1������hA>�>Ze��ln��n4Ǵ��J��{��Br`���@f�o#��:����yP���B����Q�����j32�DR\�G<)���L�I$�-b�y�Y*��a z{�IoX�ʭep�C3$�o�vF��0?Y����\�I8V���d��ě0Y����4w�KR��#-᪟Ϭ�L��y�?*����]��Tڮ��Ǭ��]#���Z�S}��<?�Q4,`��B)�ªG�#�D��T��7�V5m�&� �;���ѫD��m��|b{[��|�9uյǥ@}�-��2�1����i~�	;Vc����̏�wl0&Zϖ0R��:̆!ի�=�gH�|�K\U�ɵ�<
9s?�U�w�[�6�A���0��^š��'�&J�����|��9eB��(�W��m/�O%�L�~�V&�d����¡ucO�׾��\�	B �d�:���O���f_�e�☙o���з�X=��|�d�<�����d	�̲��,EX�@'���y�8�`�,���5��7p)��{�{�� 25�筃НxQ:�����.H�p��Q��|Y�'��~�4a$Ҳ���6��jI ��(Ȱ3ܗD����H������������@���P��Bd���J�BP<c���~9&�-�f{�3�IP����RÑ�?Ɲ�|}j���΢@A�xJo>]-�I���B�\���Ŀ�D���=������eM[�.ӀÖM�o�͖�NRq���	�T�|ڙ�D�dq��$7'
�j��p��R�}*��#�E��uo��m�˒o��M!E�jX���&x�.B,�j,��/��ņ;�3}�f�4���ɜl�_oD�H�r�>���)f���5�#����>}o)���Fu�Ο	AQDB%����l���<5�(W
{M�#��w�?��*̀\�6*"�Q�Hfq�A��ʌ�:]Qf�0��&�&׾LI�ƌ_"�d�$��뮎Jp�,Jj�W�d���qv9mYaa��}!1Ӿ�q��1BFJf>�E><y�^�=B>��d��80���F���g�#���}M� ;�.��*]�N,���M�w�9Y��/Z]�A{��$f�����/�K�]t
�Q������O�[@�<#�����<�7�V_rw��(M�W�����M)_��S���T6l:��V����XH�����!���)��c�T��6�-�i��k�|�[M����jP[c��%�N/9(�=o��^��W ͹�.B�K'"t�z�2�ZiSb�^0J �]�ԑ�91�npA�2�(�;��&[�W�nqj�+FH2t��lu�x7dy��@eD�EJ3�Ջ�0�z�|l�� |3��,����`)H�&-B)b|I�����⛈�q5�Yhk�I���\�����2���mg�3���K��`��?�O�1��5c�li�ص���ߧK��:��ê�΄؀�l_�c�~�����崽�����o�3�/O�m�Rr��@�a2�
��GP�ܵ��=���o)�$�h���������b̐~�e�ƭ���㥢M����ӭ�:�o�)���%�ޗ3���LI��[�H��3	xA?���(TOB��%�}$@in�Tـ�
���x>��@�MB�V�M^ا�q��a�f�����a�<М��٩	�X�X)��bd+6k8A���)Ӳ?�έʭ��#�K�=7y�CB��ӟ3�އ���c�A�8��$If�������
UP��~Pv��>����O!ײ����L�r&��e]-,�	�@1_� 4�g�2�R��!&�
�g�)���rf��"�j�/Z�#������#$���T�>8C�%n-7����HN�ݛ`F����D6wDO���q�g�n~ʈ�U�i=�逫3^�������\`�۩�.%�5.�c[g��< ��<��RlHא���w=r�;>6����C�`�_,��L�[������}[�GӈC/�`m�)O�ak���s.(1{�2v���j�H��K��쮑&��È�Ѻ(�Z4Q�^	�޾�����/��2���p�p�d����קj���/je�+UqV��<�=�[�2�ڑ%x�@[^�/[Qt�U�_F�Iדq�sT��zm�@/VS��}C�ݸ`e����F�����tP��tY�$�o���Cz4�z�0���jj�����nI�������I�0�ӵ>�4WR�Uh�=��v5��(�H�� ���&X�L�3���X&4�@����i]
= ����it�bg���g?���߃��B��:o�#�������f�N�tǫ#y���=��P��&;�~�:�a���Y?�	I^v��M� �h@ꁩU��<qK (�=���ؚ�z�/
���){�eZ�i7���Y���"Q�.ybz��!V����5߿{q���ܘ�~F�C�ෛԪ�����d������4�t����m7��2w���آ���ޤ�v���>%���ˀ��W!PJ��Eb�P�$d~��_-K���T?� ���z���JɎ�b湁n�����>Z���pg�?1�(iQt~�KO/�'ŉ9�<�@q��>MQ��9�0�ѭ��K�����DO��0"�D���@^}JT ��l'ak�鷷���g E���ND��mx�:|�[���urQ��n������J����!dY����~,Xj��RP��2�__�%�_�,}Xv�!HS忿^�9�+����y�P�K��A�,�a��m�9����$�B�v��[�hȕ���@ћH��R�Ά�B"���z�M$�@Vr��;�4�Jh1�Al��t��I��s�y=L��Ie�&���,��sXGM}��\�,O��L�J5�d�chi� z;{��<�����}e�)ؽ��>\�d�<k��._�ˎ&� ĂUDu ���]M��Ӫ��_�`����<�.a����	�~�i"c�|�:=���4��Q�~c�gW�@e���n�ycDp��������YV�eJ��L��qЎa4n&��"�!s9O���:�i�O������?(����~}���`�Y�������,�G��'�Nb��g0�uY$�[��e?/�tl���!e�dsU�8�c�Lx!O�VUAuGx�r�H2�O�޺�6y��+r
���;��w�3�C��QLnߵ<E���@�T�u�\,�������K�"��h�i?���p&*��� ��e�$ ;�7�u�y/�l��F�ɶ����P��5�$���LPǝ��Ez9z�L��.���(����`��-���e��Mm[ض|����`v9�j\p�zV����H�,;�s�[�ԓq(B;I�i[Jmh~��MF��V��dC��p-�ʟ�$x��W�s���K'@�oHǟ�z���X��T�@����6�w٤z�:WK']7F����ԡ��5�hWK\5�yIU+K��6�FB��F'����AC�N`�l(eQ�ά�{->o7��Zb~ ҿ����͒b��#�3��<Ä�
��/"�+:����EB�O?a��KK�`p�e� iVΑ�I��9��$ƴ�΋gzN���m�'P1�i`]�H�?MdX^9Y�y�2�I�ֳ%I�����nP1�A>�����s��q�©�+��
T����%kVJU���4i�j��呻�z}6�F%������b2��qE�}т�x���=����uD:�Ei��j��Y��9�A{+Wi�"��:����h{���aJp��M��K�+��J��H��Jg��j��y���ږ�G0RF[��|��rA\��y�!�׷��z��@���Y5�m(���T�����6��$�I6]��H�m�Sfe�1X�W�|bڇvM{����@5ot��m���k�b`~��F"��P�����9��ƾH#�ym)׊z.�#�M|�:L��g�z����̓w�&별�j�+����	hw� Xq����A.����s,��1c�=|���"H��Z�M�˖��^Qk��N۽�t�}�]R��9����Y3���vz%� �dD���q��Z�fR��g]_v����d�L�CQF?�N,�-(�_���Dhk?����n�Xø������r#�h�5Zg�f̦:r�W�=��QS�˴i��Q'���H����� D��F�˿�ȋ���'��p��~c].�M&,�/��o�&����(#&����x�\��];}x�^(��I q�H�Ԕ֩Bl�0���A�3C��Q�8�=�瓾{�K���_OM�f/�__���1:��:V����Sc��s����)g��F��:�c�p�f�J�85o&��?W@�׌K��`1)�SQ�T�hbXu&�s''�0%嚙q
��7�ZiV�QŤ��.e.[�on����"A�EĐB�		�R�_׍���a��Z��">����_3;��';k)�}")2��͎�U�U��>c���V򔉈wy��b�x�2�>�tQ����J ������p���͠��d4�䄔UXPs7��R��\�	��4��toՒoO��#}c)��	x��q���B72��K�tWK���yq���xL���7���3c���]ekd�.A�>�cX7��m�� ݂=�i�)_�� ����@�)�U��镂HkƇ�B��F/%ZeZ�4ȸ���MC*���Ul�B۫C��|���1ӡ��XƳ	���(오Ȋ.@.�{����!aZG�]�>���n�8]U��&�|:[/#�:���
sd����8�Cy[A˽"�C� �p7�ќ�������`(�Z�L����7�N�p�FwF0�1�^_������;�Y��Y)�.T*A��J���?�fM�fT�`K��_Y1�
S" ��-wh�{�e=�o-[+�MS�E$K�@�f�Њι ��(��4����MS��9QdB&�v����L��%��[J;�#2�hy=3�k�?����7�=��[o��vx�*�e� }�p�2���&a�49l���uD�Ã����+��ud=x��j"�?n��9��Pm�1~͹�m�,���$�ElL�{g�%��k�� �B�ceL.��݆�,W'�ɯ��(!0��^���ל��eC�s"�~S�ҧ?�E�B�@*����=�_@���#�C����hwAԯFg0ϭ�,���C��.�#�[d/s:	Ée�
v'u@�S2�$>���<�ή�%x���B\>���`3s$��F�E�-�|�PW��$U`���I)�A��j��t�W���<�c�=ڟl�gV�3��	�xj.���Z��`����f�+���(�@�G��F�q�QC	'�(�UL�P���r��R1��gՋ����6��sJǊ$w�(%��v�U�;�K����p����`T)�k%2���Vp\x왐N�h�_(h=��� ���gZ��$5W��)�U��R���ۇЮ�5�{w\�l���7����{��ޔF����"�%���S#�f�r
�iV���N��S���tK�;e9���D�Xw�; �wL⮥v�jBqeU�C�CU9��K��Ho����RB}�=���>꫖��?�`�Mg�_ ع�a�?�3��E�A������0�^�V�NT��/�p?��P6�+�돃�	E㞂0|-��RVb���`o�,u�}h��`���̕b#�u� ��)����N��b|���b	{7�	�''��a^��ي���8�Xo�����nW\}�'�<�nU�5��6c��J��.�`'���a�F��|^CA�0�]�Ȥ���?�-[�����+�B�Y����n*�DQc~�<�<U�P~�(�-�p3�0P�e��D����;�g��>�㐽��B@V���>z�'�i�W˜�'�7�RgƷ�L�)�B�X�y.�Db��v��._���&DE�Oi�G�:%�@�w�iqP-�x9ԦJȒ]p�0lԢ3]IǥM�0A�JB�5��=@��2�uB��c�7�Yl!+���f�,c{7݃�vQ�0�i���|�Y�|��Y���m^�?K˗�y�*z)& �����Y�Y��Vvn����9o��;>��=7��C���ID]T����,@�b}��{��E!i�n�;�	ZÃ�R�^��%iԈ:��Y[�����ݰ�߉ �Pu�f�{��X2�C"AlK&�d�p|�U�l,H�1��P�Xgxf��!6�1"G���������jU,X��V�a Y�*�iZX�B����S�P�-���|(X����0�o:�����Kn��vXA�h���kS�;wD�>�c$�_��黸�(�D���j��k��PϽc�g -x�ؤ.��d����g�כ6�8�B�i4�OVô�ɘ��'�!��!��(����eC��$�Q>�
� H̛@+�W}��D�R�v;{��(`t�"���dm�����L��}�T��t5�f:���C�}�,R>���ז�PH`�y�H��Ų�C�E;�`ߺ��jC���LeC����:�f���1 q����� �g[;�##�Zɸv�]#���h+.iՒ���G��2�Ó .?%�
	��X�U,O[ǬT&���9�����j�F�#ӵ}i�~��^3=�G��Ϸ��"�����?��FnŹ�ͰWn
<~��}�Hj��-Ɋ��դ)�ƪ���ӘH7|�Ҹ���i�d\��)/�F�{ ���`��jQ?N��nt2,s��"�����ӛ�s����7��H�����Ia2��I�j
�u�$�U-ԓ~{��=�*���k;��͜�d�X�d����p�d��M�??Pc.G��>��E�{�˱��؉��+g��;�5ǢF��o�G"~[MСD�͌���S�,�}���{����B8��OE���o��;&2F���/T�� =�<AhT�Po��}�ņ_�+}YK'2 �Ѳ��3�̇���W�ӊ�֑�´�i*;����$QV�DF@瀀7g�.|K��W�s�n��/����`���`�����[�Z��tB�v�#�o����	�;�.�ݳ6Pn�`�U	
;s��C���8���g����ylܶx� ��ՍR�c��(�$��Y� ��Yvm<0nO���Y^�Tx�0�I��j��}�-�s�DF���RG��nI3~�4ݎ'��b�	mӶHTOǪ���m~��d8��.ʂF|.��؋�ș6A�B{�g	���;n�H:�V��<�\����w�H�4X�WكI�.��J�X�l��!�V��ΣY�=�z$����mE$}��5���r�fI�ń{�q�]����@���Q9NV�r>H�d#黧�V��H��ų��nN�}��#��,<U��c�}���g{݋��=0���sR��_zOꑔ��"]��4"�U]��~��ꤡ���;��,G&f0�1��$�&I5�Q#!�⇘<��_x�(�@��[n�c ����n��څZd�������Cx=�U�>V����l/
B�ڥ̓��ݽ��J���u�6��XP��ֹ64;q�4kK�k���h�̗#,%���rS���ȍ��A���4Ҙԙ��'�7��K��yB��W�`��w��Z�H�z7q*���Vw�e�o.���69�I:C�puK@���.ف+KH�?5j*w�l��{,2�K�Hh8el�-O�(W.RFx!�� ��vf��ɋJ�#��	�]0�GVT�����8ٲ��nO}Y~hU3676XQCэV����C/:�Mb,��!F�I�!{�d'�L37��{����+&ͣ�`n��jy
ڮ��N{ٻl��9U�>[��|�����٠q��\ջ>���"�K��0�"5J�\� �ᩖ���K֬���JHu��t�
�dt��H�zܫ���H�]�I��-p�G��*(��a���myq@����9E*fu�-e2�x�I�$ܸ���\dm>+��Mz	OL�clZ��4���o
'���[HM�bo�9��'�5NQ>8�Z��^�0aq>��Ճv�����T��;�ϑ����
� ��� OԘϧ�����J�̨�ANҤV��u�Rه��H���9�򟊻݃���B�n6�j��'�@<.�[�ba
�Ĭd �ﺀ����/���G���m�x�5'Q|@N�����r�T<<}*�����"_dtHQr�'�'�wĽ�ٴ#}�@S�tl�,�	�\�|)%�.��.� �,.d��L�A�K����8�澩�?�M��u�C�@�P�s���A.�*<a�49��p�KO����,@}��Ξ�P�m�@���d^�yvV���4�!�X�7�|_\��f׳$�ZX�W,]�{�M֗$�ph��(.GP��b\�
UHG&`?�9�w�����i�;�����7��ܻv�%�AM&�Â?��#YM��#&��^�O�9���e2�!�X\�xMV9^��Xr��x<�/�p��-|}p��fkBW��l���XMƉt\Y1n���J������J�y�C�����NR7��S�k=�����W��t���]��ynS�r��Z}��VE.���i���_�*���0� �!��4Vx`p�h�Y�;%��x:m�C'�xJ�YϹ���Y$�%L>y�5V�@=b��4LJ�Yϟd�����k�f�-�|�����������*j��lE0����yE�B��� �h�
쩴0����P}E�B����|UТ8(de*^P���A��tgP�(R�$b�=�?(Fޛ.�F����.L�x�^Q
�$���a�9��xI=�P����[�,�r�ԓ�k�
'-Q͂���2݀)M���p%|����,[jCm9�ʦ�~0��qqk&:��ѫzXp�0l1��J��<\�CD+<�Ǜ.�!%�4DԴyϛc<�-���!9z¿7����̢��Cr<KNT��qW�d/x$��D��/J�􁁄���>��P�ܥ.�-єq��w:�*�`='0m���A����`n^�_�$��jz�\3`D����٬wWǄ�V�*�@N&M?�m=�UK�͕i�jn���p����$ ��ޯgI6t�δC��E$���n����1R�\�x�B��N�_m[��ƹ�u�yA��[���B���[�+}gD��=ܘ�|��Ӹ�&�]�G:���g�aae#�g��L�����`h
�zCK_��G��a~��	�6t0]�m�e�gCP����������3?��A�w[����/J]X~�uū�b�Ӆ'�2y0�tp��-nC�-�6��"�BWF��`��/�|*8՛���'oGkc)�b�`���X���L������u�{T����u$��߻�cx�FG� �mB��*�YpLO�4���Q�II���JUH�%֎!���XNӞ�L�n�f�����:T/�t�75�F�ZS��Es�^�ڃ{�V{`���H�оW��暈98(������:�Ev^��ᒄ1 &i��u^�ٕ����3����bMS&:v��+�Fr�C�ǵ�_Z�%w0Vt���m��4����G���i�� �R�e�MwF���g#�|���J��A�K$��(Dϱ?�<�4Y���-� k�L���u��)��v_p�x�eP��R�s}���U��i�>�h�m�2��+�߈�6��Z�H˪ �b�:�#'��-4�tẰ�+��.�ůD��W��Q��`��U�IdZ�]��r[ ��㶬X�F(�`�F���`�|�S����\�"$y�h��LC�$ez��Ry���`��\)��3́F�<̈ m��y&P�眠��Ը�\M���!I>�E
�����Xd�N�+cFBzG	������m5t'Q��0S�6U�u&��P�ô��lh���?����y���'�퀭0եߨ	#���?�#�9/��{�؜5�M��A[����Czv��;�3�@#*kd��/ ����u�-��m�Ck�lp���#�X�����}38�^�;��j0�)m�tHMH�h�z�Cy57����[��V�bY��ٚ��\A5����5��V'��f|��k�T��7�]Њ��F�K{�蓽�����Ҕ�	�A��p�ޕ��W@���k�X.�/��M�>���p)��L߿^ho��U�rC���D���7p�q�P��R������S�<o�TG�rH:/o��o�M�R
�<�e�a�
��g,�I$��K�:&���kK�/��[�=�^Ʒ=��_ ��hG?�J��AhoGfR�J��7@�!�z�|�������W=�o֤6��|@R̉�-MO*W�:�:k+a"[r��O-?�E���7�0�ެ�Y.Ӗ���6�Ur{É�!C!4�H��݅���j�Q�=۹nu���9?zn[����-�����Ξ���ũ:��ک���T��Tt�p�?��ⶪ$�����̓��|�TEW�����]D�zv�#c���owz~0�a�:Cܰ�l� �2{���n!�`G�rrub�,��y�y�9�%7C��u��gk�S�H�Y��y	 �P���ZlT�d�8�09��.%��vI�pF��<�J�����{F���?��ӎ`��3Q�}�~5@s�l��ʔĩ�7bt��~�_�w�R�2��d�[���"�Ҧ:��+ujF��x�rN�0�r��������d�+<ܕ	��i�R���=�@2��9Ig�م�-��:�:��8����FQ��{so��ol9������ơnݽ�Ҭ@��R�K�3xK���
�Wi�8=��p�'���P��j��&,]AB'�Ml��,#�w��u8XM����d��)Fa�SjfB��~�M��̼�e�O
�D�N�`P	��f\4��7.2���o`t9Bj�1ڏ-�*͙�;�N�U���W�z�)t��G�sǱo:ߒpT!��`\�+�G��C�U?7`�wE��d~���{���J���س�d���;>g�Z���u�E��m6;բXӝi4�\
~um��􌌞U$j�Ɗ�,1�K�=�aUi��TfYϱ�r&�6��W��b�x�:S��udb��P�&0H�4==��<����0�:���no��a�v�x��{�5�6��G<��H7mǵ'6,RM�sF�|����jq��5����a+<pZnc'�:B
t��U���!�d�%)��XZg&�d ~���4�.�n�lߦM2
D����.�c����(Ԏ�4h��<rsC]���t���(?�]�5���߇�ty7-o_t�[��0#}�����9���Qδc��Z^>07���̐t�+����0�B/�G�<�y�D���v�������uwEa/֡TE�T\�+J�o�V���M��UUe~\��R]�����o��_�n7 ��Ǽ?�$W���j�q	4^�a��rk�l��i�߅��n3竦&����9���B�z���Fv��U;�J�(���Da��_�''� p]�J*�_d;��΅/�&G�b3y�e����N������VD7[��&��ᐖqPƤ�=Ej�)2D�a��Ѝ�c�mftg<� ?|�OCĖ��S�u�'�;{Z]�G�CT�^M�:)����Ɛ
:�1/6��uQ�`�r��8�hk��p:��M����q8����s����xaR����Ȓ"�c�%�:�
���-����Y�ӈ�l�����d(<w^�8�[MD,8�g�W�����f�솳?w�v<����-T�/��
n�l�~�,�;)��;1���(
��S��J��Z6�ԴTNq6X#u�ƾ��4Ė�҉Ð��r.���'�0#YøJ<�z���/� "��+�F�I]�����}���[h�U8Z���&�K=29�i����Y�	��s#B��<uL54f.��~kr/-j*�hIsꗪP�0�KJƘ�%jN���KW�$�m�G�lM�*y��=�Z��^(1��凉g}Ϻ`���l0L|T
l���!2�/�A6>2��8�c���ʗɫ�?u�����Da+��:A��>�k��=W�i��s>.��7����_�:��*}��r���W
O}���uARwmYN�]�i��aG�ȇ0Sz?��`
�`�L�u��P�	$U�S�ƞ�Ӌ�����Ǐ�x���pٜ^q����4�_��m{��b�ݛ��l �)x'?!��5�評 b�ܲO���CM���SU��≅�Iu$-9q���I�B<sv�E�5ibʶRemj��nn�E�]*S7�k§�nu<�����d������J���`��h���7�D��$��{0'w��21X�?b#\?���d-A
���*��`~�����Z�ׄ���B����p�J��}0�U� ~��w1�Y�F&��+N��=Jc�.{\"�#�-B �̢?�\c|�����	�����=�- )tƿ\|�H��%��V$Jq�G쟑UL�_ʘ��u��
��Ϗ�Yʊp�3$\$3kCi!� lGE`�3�����u�c�O���`K��hJ��ɭߤ)e��҇mN�H���������n��"��~?'�S�c�~���o��r����a�#^�p���:��.�'iu�����l�c�X_��7q�A���r�v�0ƈ��8��n�CMv}>���@S�f}Һ(�v�4�V� �8Id�U4R��x��_�T	[��DC�z"_-X�]u��c�.A�[�~�����H����C�rV��g�_g���j�W��D��N_�c���-���؎1��^�7�N�����z�Z���#S�#�֠e(�m�W211�)��#���U\."�(	��i��2X�����(OQE�u��	6�g��!�P`a����(��,<}Ҡ�ˍm��3�K�/!���^�I����p������[7���o)vaƱ�O����3$���&NI^�G��_`�ޞbh�����/�������M�R��TxQ,k��F�2�b���]g�PvM��]�}�Հ���8���)!��1<��@n]X�b))�[�'�4����j�&a#���WwD��N���R�%C�1���l�9�n $�������:7����欀���'$�M�� ���v�k�ZA�K Ӿ߯�.3����0�ɞ2�_�o�H>&]>�Hn�]�0���q��\K
o,s�Bj(�į�{��q��t�!��~� �7�9��;}�@�&o"-|�hV�CQ���g5j��W����b�=��<V,aC�~4�J6�ʬ��B�m-`�N���(}��H�W�C��[C]~���{ep=�Ưi	��v��Х�����QT��^`d��Zj�ڎ�T��Pv9���C	L>���z��Ia���T;��#m���8p�IgD��)1	N& ��53[�%e�7x;�l���;�s�p�<����ߐps��pP��:"�������w�C�����4Q8\�4���i�I�du]�)/X�~u9Q���
�����Ryǻ��
���!��á{5�
�}��l��`�K�sxH0���O����9��Z��:��E�}�o��۹�'[Xn]�C
���h�ZzH��c������i}l��"�5�R��< c1b�EJK��ܒ�%�<k`k�j��jڶ ��y	Ĉ�Q�p��Hy��Ey��fG:B}SM�`x��g�8��♟R�7�T]h
�f��FX˹�ϲ�[����n��� �Ae Y�3\�c�j�l\�Qi�7���eq���p� �mZT>����R�� �0us~�ݩjb$�3w�`�n%G�Ք�u z��k���X4��1]���$��䟅�k�9�B�(�����8�ғzy�_ j���%��ܶ�����+hS�=�8]��w�ћ�_dxi�g��E䗔�g?�?<���u�?�=�o*��ғ�f��VJ���������[���K��~��	 *?Q�*��L�U����1Wv�[�k��҃�dĔ���=��ǈ�2(;��1��Qe=�d��f������^M�3�U�f�a��v��y�	�d�n!��hqح@a�u�$]�m����R-:^B*�'��\zT���.�����4gKxS �]���/Nxц�����g�AZ\�uZ�udH�%�Ap0սoJ�y�*Y�u�Q��Ӆ�����x��#�IqUӉ�Z8Q���y-`?�E޼�����:�L ����,T&�Ztnut�K����f&Ѿr�n����������#�I�PP���j���y@�-��S�؂�yF���`�s{G����eJ�t˼Z�/�e��L���M�1������&�����  �#�CnM�o��(���8b���Ӝ6���7e�q<&�y���V�^��=�)Ŀ��[X�1,�9u�ޟ�g���2����V9�u��������E7kD���_<*Y�?��'�哇�&?V�m+�������ܣ�8��@H�:�NE^��O�I�4DQL�*WKK8�1��(�������IBh{��e1�2����(����^�Ir��w"߃z���)�ም�P��N�U��ҏ�Z�d�R������`a�X=�z�I͖�,��g�$����ka�6���b��T�[�E��'��|H�D6�w��w�g���blҪn���EM� :KOL�(y�c��xBj鷺�%P�jf���{��2᱘,V���+��|�4S춪i�+�$��u��*r|6�=���ЯV�R���Y {�Aǃ�JD�gE��Ƚ*a�7`���$S@xd;^a	�����w��Kv>���^)"��$\�
=���bt��ƍJ/�n��Ē�3P��5�H�ݳ;g���K���EOD.��Z�a��dh����{
� �`���d��s�Xx>�(A9���*����{�&�J-ѹ�����+�v��[�N��!4�xyo/v��]����IW�z�O`FS=#8�y�
��b�p$�z��N=.��9d� z<3���S�� �����Q��!H�� ?��_[a�)@D�	�L13�d���f ʔ7��|If�0�$��d���Y�jT4�ћ�����ɹ��$V�v�:���E����K4HD�oI�fV#����BΦ�	�*�g�8Qh��:Mg����cS��dv�A� �	���Ҟ�,�!��=l�Q��}rG����>��W	o�V����e�2������J��;��:�����vƭ0f g+�~��������ԧ!�5��G�T)	R\>���q�AM��0���K�x\T���]Ή�?:Ͷc�X��	���ؘ/�Mz� %��Y����K$z&���觪�/R�J���	��� g!!��OX�I��>[j���ҝ@�-okZ�aJ,m�l!�>
o���ÝU~05gmg!Q��5��O���ğ����#�<�2	�,��W�[~Fj���%}���dA�
�݆/X0�ϝ� cW��
�Ӽ�s���\t�Q���ki(�qT��7�'��%G���)�Qp�`��� �y��܉L������w!���V3�0Q�ޠ�D��Q�T
��i������R�&��M/��VAL����^f<�ɥ�Ǜ?�@R�:w$�݄g��Y��t?�+��{=Jgg^R�|�A�L�=T�oS���0��8{i�[G^�&k�P�''!d����d_���Ħc0k�F8)Ԛ9����[�bAU���X�� ��g�]�)�N��=T&
?���6��=ޮR
�q_�WZ��8�T�wp6N�P�2
,�?�;|[ F�����-�[�@>O@�HDdG�2>.[�@���Jq���D�v����e�$Q8hރ��ws�w�韏�=#�[F�����I�r],�b�A���$[v��~ʬ��Zآ�sS�T��5��oC̝xu��D��8M S �ޖ2vyn��7]���w���k���>0g�ڀg����]���#N��߿	�RHsU�.�_�43/��4�h�x�-��DYTgl׸}�2�y�|�JƝH���o
cJ�~\B�Ǔp�&�l��6S�a	�UT���i���;�m:�R��t:�p��Fz�Y�%�#3��3�R(a �3Q�L�����@p�D�WF�B�}ڭ�+!b��0�D'���wR��):��b$���o�91ֺ&˸���i}).�>ьX!�0�&�Jb�q	��Mf�ƣU	���<�Dw���C"���-�d�?��t�m�Z�Aiu>������N��S7�V|R�S�.`�RV�0f��'((��S5��'Z���u����4��w�oA��vFC�`�"���9��5��Ov�>���bI�YΫOh@TD�ƵLҪ��~V��Qh�o�g��U�>���X�8�u��F����M�3HY�
�H�+E�;��cպ��8��i�)�N����e����55�-��t���ffۯ�N�m�7�u�q�;�ZQ�N��'�����r^F͕��d��8`|�¶j=o��	�  �; Y�g������&p�R�|�1���Pl�h8��SRf"���|���i��_S��τ�W���sH��Ք���C%[}7�3D�����[�7��E*�KPۗ,�m����D�E�v��eh�!�L�5��wn�i]������Im�����->���~!�˨x7um�b���k3�L^�:iJ�f���u�~i@4�K�$�{}�X��M��+� ¬0�@�Q'�,�{��ի��Z.e'�?Q���[�Y��@%���3u����]�),����B#���TY`.	����7�����}j����q�.���6<K�%��[�k���Q�����w�����x	�>xv�z�5�M�3寔���:Zt�n���~
TZ�]ҥe�5v�(���.7�C��]���=z��FB6�yC�C�+U"�]30���RKU�'Ul6�g��
��ԣϑ���ý��I��YN �
�2Wk1%�Rr"�ğ�W=wQ��v���D6����c�ת�����p�V�|����P{���t\�	��ݐ�Ϛ﹋�Ȟ�7OF]�,I�|��lk�$��s'��d,�޺���_��:�R~�V�I�ūLP�<�+$��CF���B]���<�k�s2�d.�֥�j�RTo���.l�-�2r���z��"č���;Q�%�+>�I�'Rx���}��@�l03H�J`Qc*~�BL�]}���>�2X������9�P~���YG#3��U�=W��*� �dJ����H	g����bZK��P�Ö]調^��*�����˙ by�~ҭx
��D�S�	���l�1��&a�wy�z�
�s)��+�C��`�c�
~+w-j�����K�TKc�cߛ9Q����C_]��c�����Hx�[�P0�=������yAaȇ̯��Ms�N>���Dqdw��1��#�n9GS��>������Ty5`���'w�;�g�/1��Xݤ����UO�Ы��)p��E��
k�+N��� ��t�$�)���?��ޡJ���2��t釥/��x����}|b���	��NWz��km0����m"W�顏.!]�E���{B�L�i11�d�QP��x¹��Y"fԣyZ�?�Õ|�i��r��C"*�S$ �S���@P���\��r�ח{.�QF������Fӥ����(�̕>�&IM��x�j�f���]z)�����Y)?�h�:wb��V`3��R[���Hw{Q����R�8���Ƀr�,�����MS���R�i��c)����Q9@��"�l2�G�	���9Xo�6�Gri�1����NoP�L��J�-�V�2�6��i�ķ��w�!0�7�>��X�����p���AϹ��G	�?�n'��wkh�N5� 
�3���)�����6�ٯ��8�g�G�_2g�Z�ssr�i�'\�L�BtTBEWe.�7����l~�r�s䯷z�NK�Gx����[S!Ya9��藮k���9<�Ȣ��������hX����c$_�x�/!.(,?������%�%	�Qed(��no����x�^/��H����X�����m���9u���ҝ=�n�U��i/>(�$����D��`���B�ic��&�g�^����3�z�t��Mؔ]ŕTF-�8;}^V���8f �*�@ܹ�z4�������)>�2�Ba��Dh��_dv��v�82���:;)X�xRn��}p�>���,�y�Ǆ�,_�]��eRF(���|�f�l��DgQ�}$k^�R��9�n3���"428�N����잳�*�(��Vu��]fS�}.�m��0��sV�E..a̡ߥ_�,����c�/k��5���1��n[�� RsLԚ��9TwbM�ū�����ɺ��\#D����ne܊n}��p*��G��w�G�Q�"ں`���l���S;���	d�tC���y�x��z���%i���H�M�d��d0�LKe��hp��p���>�Bh�����?��qo��*E��c7��n�P��8�Ŗ� �P���6�ڊp�XV�,�4S�p����}�,'�*��C�,� �t��&$��LYy�XQCH��&��T;�y��_ݭ�dˤ�/�y,�9�E#�R���l�A��l���օ<��@�i��U��b͊� 7)6��.��S�,T��~Wx����"��7�r�k^l<q$Je�G�k~G��U��yء. ���)�����i&�A�R������P�1�}l�TEC?P �ؿ0sHE`"��m\�^���B���ϵ��+��E�
yaK�c|��l}�k�����/����:5���ؐ7]��s.�V��	>�J{��l����3@%߮��R�s��R�&���T�
b���)RpI�)�ŞJ�v,��rnt&z���4M��dJsmiz�r�>0r=�(c�p2.p�VLWD�%�z�W��aМhnٮ�,Kiɤw\�B���G�a�HF�PQ���7ܯ��k�(ȁG
���1�b�'ū���6�8�'!�@��R�. �9�p4ȵ���AKy�g&�D��T��V-(�R�Hm]��l(!)���o�L���v8��&�� =2 [��&C��S0��AVY�u�^��p��UM��ݮҦ��P1��z��=����H6Ɵ����u�L{�=͙�������'�Bh�h�#+Gb����K�`�=�����-qN�rX&�mP��XI��Vxdz�����􈯳p!@>��/?R��������XI23�e�T�i�W��7�L���ڨ��!
�;3��:���me<�&>RQ�?�_2��"���	L��i���$� ��Ŋ�����o4��8�
o�'k|�(=	K (e��(��-/r�(���B��*K���m
1Ʃ|��}��V���Cla��6Ss�W��Ս�
0���k�/O Z�C��Z��0ŚƐym������l�A�F�Ey�n�Y*���2�ٽ�4�����<!C�	Z��1�v����Dk���$�;pLQ�z�G�i�9s(��x3�H	o`x��U$�j���s��6����?���S�k�d&������n.Ch���N`�ߚX�h_�xe&����n즆%�Դ��W���P�ǟ��}�ʲ����X9�~�l�~ʷ,U����am��i��22�.�]���F�Q����k�{-�o��?0}w`Ǧ�>���v�
�w�]���S��&���LoZqy���h�?��3�hў��:g�Y�������ŀ�:IC��A����獀����D��A�ͳ�+5i�9��u���Z�J���b��4��	�'({�6��{ƻ�Cl�/�w������a`<W|,�}��@�`�Ij�u!75B�eG�ݪ8�If�o��b�Jdw�{��������|E�K��A��ئ����K���h�X�����iҹqq����xwJ ��3���� e�{Ŗb��T$\wQ�{�����R��"z��ȅ��=��u&���m΂!���N2��@+.J�?�n ��B�%������G�E��OP��b��n#��G?et�>������3��s����+,�L��������Ŋ��(�[��П���>^�M1u%[�i��zZe�Aży햐���ϐ��:��
C�Y���>t{K1��8��k�dt782Yt�=�yh��fgf\�=%)�s;�H�:�U��)y��� �']H�l��.;��/'� �)�����kEe�UP�$��t�;��%�B˹���O\�G�P?q6
�;`^�b$�c9>b'�ǟ2Fŵ�H���y3��) ��=E�S���1�<��A���d��`"&X�g�[���+K�\��������	�Z�/0�ە�l�qpZiE�|�Q���$��+w��0O*p	��Q�a��ΠldV�ގ\�s$�P�����[�X�`,Y�hHBB~����̇��s+�F���}1����7�X�y�,yt�H˅ejD��5�#�0����%�����!8�b�m�oW�%6���c����3.�Hi�i�sᩪ�@�S	ї��j��"@Xw?7�c��c�#P��x9I�ٻ��CC�H�_��Ҳ'r�h�[�UQ��u[���G�-Jg�^9%�H�4 _�0�u�ן��H����4�A~�ʤ��gK�21G?QJ_ӏ�	 _+�1i��@��A�w��|�:Q�`��Tq�����~BY�q�iI����
���ߠ�;J���I�2̞݃��F#���[ڻ+6�i����COno�gǱ��_�����uŸD�#TA�$fm�Y�+��	'�}c�	7���/�a/�U{�{���+H��ð��*�T�l�t����-S����ޱ��.EJ�L�<�j�Uy/^�Z��S�Ÿ�ӗ aȃY��?�:b�k4<��߅���L�ǋVr#��X����Β߂G�nlakγʅ��9Dp�L5aZ�Ra����y��rv6F梇���]:ez4�0�5L�'s\��.���+�a�2�a4�eP>*�p��K�)��е�;��k���ƿi�Z��ր�"fm 	@̵��%qR>�EF�^YS��VO�!�_ykv� 7�M��C�9�2��j��ɴw>�?#��RXA 7���YO	,?)���%�}�"����S�MR�0��D�A�u!����1���Z�o�����=p��Bb�"$�3c(�>����@�^�Gsٖ��/2<��Ĭ�����7� �=�y矰*]��2�ż��?��
֟�8E��{Ӛ���3RC�_��v��]��$ꐼ��=M�PZ7�P�8���}�Y#Rp_���׳&�=3rg/������o]��G^���l�7�=}�NgxR�Y[8wv��qhW�W���oOF��Ș=��^3�G���v��!2�� I<V�d�����Hk��PT�VW�$��]�2VC�J<RD-֛�9�H��t`�Ae��#��CO׾
}�j!�����Y�4$������z+��7�ٸI�� $d]�_E6�9&�Qn���� ip����Z��c"��z%�+d T��ſ`H2�����$��!z*�&��"�|�����H�������ǃ�d]A]�$X~��4xiEYp���(��\TC��K��:��Ʋ�����t��M�v���[_�F�5�_Z?��/����M���4��*�.0���#�3B�.��L��8̗�(�y�e��9�������u+8om��ڞ�^mN��X�i��z�w��w+�����Y��/���v�1��Њ$r���G��N��Tc�M����^%T�߬{)�Y*Y5G��$�AFX�����Ԧ\V�ҵ/��<����)㝩���?ڀ�*	��m����
y�_��l�>�N��3=uծ�J����3�$�g��g�3�VǑ0o�ʹuʸź���$'� �$�%����EH�7OL�4>�ߕ�-�{z�r�6�]9�-pj
ܝ��H�4X�ڰО�Oز�f�$2�0m��~է�����������#/�Y��[^�����P�~�q���];&�<�0v�D���k��7V#H������YP�/�\j|'}ֵ�q�vr��M�m�$�
��oH��4M:T�W�4U�p�;�@���JyD���� �2בÍ1�nQp\��~I~G�b�m� ež�9EaZ (�I�v3U1韇��Wb��d>� �ЄD�_�N\[��������jaU�l����V�����V������-��u��zǠ��m{�ϸ�X���?a�5� ko�]�$�z�����,�N���)��g0
�Q�pU�,���z��Շs��P1�d䏔W�a߲Xބ\�ۚ>,���Д8���✖�rc���=D�� i���1��&��D�6�Q[i��oz��37d��{����ǭ���Q�4���Z���y�Ԋ8�ﮁ�%U$i����u1�f�z�. QŊ�����S���TZd�/�E���G��ܸ5��QQC�0�դ��ύ�d����`ù<j+2��,/�l�[qڰ�bf
e�0&�(_ߔt[r(�W=�y����M$���TC�䀓;��A�=�8w�C�i���s �*�z�vJ]T�[S5aE�l�`��?c,
�R+8>0U��s70L��A�|!�����(�c37�SuČ��5�O}�a�0sUBk�y������]�0�B�r%b�d��3\\G+����I��:��G)�`���K�'�Evꨞ�e�c�+yW�����m/��F������
k�XW@��o�QDPa��L�w��q���&1�y�@,�x�{�����\"?�e*�C�	�r��0��O�c��(��.�[x�P��(��u(X��2���P���?��dK��`�L����c' ������:be֩����x�BeY�n
CCO��kl�:�(N��Sg�Zs¦2k߅��)�Ǝ���S����n�D�IaX}h�l�>���2εg�!�|S�n�o�,���T���80On��V��U�lF�A�Sp�'����e"}
��܏x%�D���3g�g��Lj��lƟ���G�ݰ�<,]z�f�GhR�Dԅ��"��:6�\a�k'�H A�^�F����0�3�%{���ӏ[y�P�gn]�
��	�XQ��PMq � �D��7g@+��2p��r�qT�i345�r�)ڏ:o�Fp��J��W@anV�~s7�*��N4`k�r�.���f;�)���� ����\ڏ��[�1���R�l���x�oL��a ^��ua���&���3�ц��@���,��������\0��o��7�
���� �u@~�X��Ȁ��JG&�:D�+,�BN>�꯴BrT�	�B{�J8��h��fy��(�u��u��!����`4�R�V��L�g�Zcߟ彿��G8�������m�A�P�T��C3P�^�œ�6l���V�wbMlkX�鬚8��=]b��qr�^���R��S�c�-y�'�wH17��̬�M��s�@�i��1�64�u�rGR
�����;K)dxF�|�l3ie����~�N����񻝤�g� Շ�i*�Z��M��j�JL�)�R�4��}�ǹ�۵j��dT%_���J��R?�±yJ�c3��0�)G�4Qc�[^	E��_	�$=�f�49ˑ	�=��FAb�W
�AG5`I���t�y\��gW돗օX�ϛ<zg��߃�l��U}�e`g�*�T�)�yP7��Jt�/g�59�㶋v}DĄ4�s�tT֍q��E?ىW?��h���"��`��+ Y=�K��1$���4u⇜��Ѷ23H�h0XT�ϼ�s�����=��b�<�a:x���ѹ�_�=��p�lç,W�6���y�l���l�ͷb�.'�;2o�HT2">aV�Q���ڸI<��NĘ�	�?�i�-�!�B� /:u�6I��C�}��p���
�݆�ݗ�t��
a��F$A>GQ�)��2k��ͻ��`?v����#(�)z� D&��D�(	�q�'��5�����F71�G.XE�P�!@��Y�n+���� L��B��M��$�H+���H�-����%�*լN鯖zqT�jb�m0J֖��w�����0b���Hj�Ns\���V��D�]֢G����&�g�wn�v�m�E�Q+tW?:�+�� ��A��X	�"9!֢)�11W�ᵶ��'r�B���(��jPD&��W^v&=���b2�7_�4�}�"!�T��O9*�%nptŰ֏��ǦP����*y����!�E��-G����9��qV�q�$<��&���n�wZ��KU��=����0�I'��LUʙ�I��D4��mڗ�b
���B��<���@/�;�ΗS9ק	~U
bR��W�͹��Dc�U�1Pq��2�����7c�!Q��p�^ �?���6��W۹�bGn�H��f�UuK��CΣ/��)6W_�$�xZk7�K7j�8?x���V�����ء�o�T�5��r�BF�-���j��,�i���{�n���4����yw�Mu*�mc�?!��q�F?��F���<����FX���gm���9 8�[u"���t�m�2��dk#@i⽚��[��>�Ba@
�#OG֢��}�84��*����)�6<=c��u��Jr�_궯N0#�gP&�`i����e+o����{h�D�$�l-���Uq"����6�[}h?��<�MR�7*(zD Q���Q�i2���Î*�f����z������<ɔ�Mӫ	�הk�#-(6<m�g�P�.�&�/�	Vi�S��)���t�����Vv�ɔhnG-ׅ�L�=!3V�p�5�¢!m��8��Pp~����!�F��f�&4�eI<ݟ��JEp���ahf�W�������#o�P��6�̟(C���c=K/i_h�P}���,='�	���;��R��Hg�5�5'�"�X��k�:Sj�f"��D��M6�����'r9\mu��-l�ژ�k�x�����?�3��I"6&!L8b9o����ZH#�ayY'>��c@���!Y(�v_�W5G���f6;������$ �k��5��2)F���Pw�4��E�B��ر>�m]~�B�yT珬G{�D'Mم���g��1d���]�]����x��7����!���2�I3����9��I eP���C�y�Ao��j����s��
�d-�'W"�x��Pz���˥�I^�����$>�,�Q�;�h?@,7�d	,�A�C��N�G�ѐJ�	Gd��u��h���_ �D��Wb��r/R%���-�x��ls/���H�|Z��Hxʿ�q��"�d�񨸙hn����g_�=x�%�ɑ#~qbY���!�)5UT�zZ��ĕ��v<�j(M+�o��0% ����4`�"���ܬ���������i�4@��9��Xw⡸g�����:��#bl�sѬ��l�H�|A�&
1�;��]�_���3����`����}�,eRm�ץ�ٿC���F�"�����p�wп^l�����Џ��H �����Xhy��Y�Ls�s�U�����GZ���7���I\�����o�U�����>AF�[q��< ���m%p𘪝o��5�Ok���|�4E�m���H�D������'{6*�� ݼ[� �hc��j9�K��A��&���v�����?�c��!�u��Wj�=m�*)2�
��9� SM3�#wh�u�Qk1j,�D��;2�g%���&1"Ǯ�\�����8��w�X���+Q�]���%wv��0^����:�<Q>x���`���TF�3K��z�>�)����Ʈe�f���`@ �G��f��Lo�$���<�J%%�A��-��ߑs>�hf(�
�0�Naq�!��^+m��3ܷ��`猥6��)FI�	?b-�$(P����\(/ħt���=K$\/+�A�v�
�kڡ_\�-��ó�N*J�\L��XSP!�)VIcucw��Y[qHѮ�dH��5�'�ҳ��f�.Ĺ/�Zg�He,h���t������c���ͯ��֕�y�e@�l<��%u��mQ��̚��\�q8�?�K�[5d[o��Z�~�s�/c�����^8���ʹF��g,U}�e|]��9"���!��䆟p�Ǿ^-��B���ac�����F�Y͖���tXdoGj�cH�h$���"Z������lm���WM��@��H6;Tq8��7k7Fc�"|�Ϻ����4~��D:#�[�U'�r��h:��~���w�gŠ�ۤuQ��lÃX��sl���OTc���*r����gށR��S�sVX*K�I#s�x�QUn#��`����I�+Vw��}��Q$���<g"d���O} �i��Le��S���"�Y��K��Qґ��U�ޑ�&��$�&�^�t��V��z"�� KD�Г��� m�/�[:��jtD$���Q�.b����<*I�������ʪ�} ����ɷd�� !�0�������Q�r��dR=	<�A��b:��A�J����o��o,ɕ�	��7-���.��u��yZ�&�(n�� Ky��v����T�ǈ��RK3���X1�U�ɲ�:/{���ő'�8{���3�&��,��V��Y����ߞU</�tDdb����̣p_�e�)��Wr�DR��p�4��߆�"�D7_� �-ID1���W�iB����\@^S�C`Lu�g:�k͒��:]���#�$��h��G묍w����2�X�(�p�{�:M��yұ���N$#��a#�~�N{��>w�j�0`9�:ͷ��ѧ�+�~�����rȍ7��� �= �y��qEк��<�3�ў:�:��QE.�g	�N�LU�@�Vt�-G��u7�H�3j�֎������L�B�xwT9з��U�ȶ"i�i��_.cӏn`|$�0��YS���]��I�84�%	kC"_;k�I����B@��b��hf��W*)S/P��ǟY�����(���!s}��H�B�"�Kq������5xY��q|92�;:g��{��W�@x:=��L�p�Y�ҟJ����7\��"��+Q���f.j$<��/�%����K�ͭ8i!�oP�y�\v�g�7��0ޤ;oiuc�	C���teQF��cS�Zl���EY{S�&|�l�	w�H~�dF)��V�/,*(�H!�[k*Μj�"���N=�V�/d�^��b�L$]��B�_n��~!(�Z;�e!�b���0h|x�'s����gδhXCy��4������~�.-G���'mc-t��C���<�舖_���w� ���^��n7e��#�0�B�s�@���ˊܱJ�c��|�}@L���F��JXc�	V�X��5� AZB4K�~x�f��*�����wl8�����7����t���)��FD����]t������ٝ8��(��b��]u9�����[�aB�~/X���
�y=�k���U�B�����ԗ��t�\��wE��w��!�kD�`w
��aa�NgL�<���GU�Y�����u?�Q�U�V���M=e�.�Oy	=_��1��Ɋ�ݪ�dzK��ׯA�y����/����@s�ሑ(_���H�ݒ�Q���/�뺉�D�̈́R��~�����s����nM����a����%��Ҭ�K�ƽd�\s�����>�ɜ};����U6)@��	��*s�eK�ށ���FL��h�:<�!h�t�lLN2*�<H! D��Ƃ���!���������g�-(O6���{�����4�;�Mm����#N�b�s��䜚eމ��v�R��b137�5�NO���ޑ`�g"rie�u?����c�tH|��B6oi:WC��Q�r�Z�c`y�8C�%b����d���ٗ�`ϖI������������W��!l<��ݱ ���Q���;��8���	2�Imv��4/w�^�&�=��~�����E�En�82��YJ���V���J���J����
�����0;\�τԥ����͚�E6����.�+Y@`S�1��}�x���mʧ��ew�a����-`�Q�z�W!]��J�)��G@�$�l)u?VPk@ѐawg{Fܓ;��5i� �n��H��(��?�k�:��і	�_�s���Αܾ.N	v��ڠ;s/�~�؝�3
3�h"��=�(e�F%�r�g��E�,�f��~K��+���i��z��9�Dg��Cy��dһ�4=�T|�	����y���\��%�:��]��S�H�Ւ�u=9u!>���/���m|8�jJ�C)����\��`�A'������#LrC���9
�_Ґ��1i?����bۆi��s&������?��x�&���I��i����0�ܴ���(��L�|��^c�����g����F��;���z"t#�W[�㐫`��l^#���=Qk|���7"*��GI���	��Æ�j�@��h����"s�O/UT~�N`��9���:���Uhm)GKg�(����{"x%���.L�;ĸ<#u�FJ�:O���?{�k��]�?2�+l`@��|������f�����nk�~��}��V$�8��Q��� *���S��)�9��q�"����to���c](}�[��/�Td\�4'�������9#�-�hѶ��1�b �E`�t��JHq��O�E�o����	�g�Z�ז L��������$���+^,�9�0�nܺv�E|��ؔoɷ�A�_5=IE��6�Q���ހ]d+���!'�l����8כ�+�����yn��fj0]�����`�
D<�S�Z��s����#�a�M��.EʀX�G+�H��uL��p#��;#�וp ��Hٺ��_���>�YxY��ow��D!��-��"٨_��{R�׀���>��+�ك�p�P�6���oJ���m��E����N�R��Y���^��1�u3D���}s���o2�z~{-�����@�ee7bA���Ow��t�z�Hm�d7���e��У��0�]TE~����X`A-�i��BG��i"��#\^5%,��IWvL͗�{��qØ�A�v����L���A��c��d���e(��3ޱ������K�L�rW��@��t���#�G,R8~h=�4�7��[�{���I�e_���/�{�z�N�ipW�Ȑ�ڟ]78d��߲I:Qx�"�ڬ/t�T�uT�8����=3��s��X�	e��<O4L�=�t�����9������R�f��eCa;LV��&=��2�ݟe�[ӡU�,ߘ=�w�JE�������G�L�YA\@݃{��f0$8qe� ˸����Lû�~X�O�C����S?rd\�갈�Ap�g*�1T	{ �0�K�A-�i��\�ik���FWP�"�#_�<lA��R�D������8a8�j{�m�CR�ń.ڋ�aV�|�S���U�:��I�	���ڍ%?�>4}/�ޕۢ�}�4E9�%lYe�i�
���H�m�?��P]q�;i������j���eX���ٕ�/Y�o��O`�g�}74i#"\����m'0Q?�yT�xl:��9��:��&T����j���_�!6kO@]�՛q�aT��U�6��;���n6�����q�I�m���h��,�����<���	OI��`��(��AU�sG3M������k'���/��L��Luh5��ـ�펴��Ic{��h���ȶ3u�3cCkvuS��~���JB$�U\M�o[���ޥGO\Be�UN�ҡZ��w�y��<tљ��K�����с��$9�bޔ}T"�`z�O�a֬�:�%$E�5Yd�y������:9a�����Ƈ��'	����=[�5��`7����>qs��}Z�"b{��0\��ϫ��<]7�A/�Hβ�M���L��yVM9+r`��h"��?�c�/��58P�h�DA�'�۲�V�{�z����Q��G
���ɯ�
\B;�$$u��ҦC�#_J�³s�l�E>���'�eދV���=X^n %�[LS�d����?{�n�X����ӓ�> �ȶ����Z���ї���)7#��N�m[g�X�)�
�Զ�!!dw�pMO� ��`|��9�r&���K�AJ�'��XNoL�B�9)��P��^M��5z�����l�3hB�3� �N)^b��G��n����Cε��4���	��~y�h�̵)()LMr9�qjP��ؽ �P�-D����Ω"��P��C|6O��-���ݭ��S�ץ�а��a�N\���3kdvW����'���|��@�E�=VA�ʲ!f�C����t�Z��I�y��,G��X�_*U���8ڛ���ҁǔ���ez�"���U!���:\-ܶ���~��C��H���f2O(a����oG /���,�^���2�M==	����_kJf۾���r
��D��`8�����'K0��q9�Dr��4������*��Ta;N����Ja�+��$a�
�\p������Y����.�4��ca/n���ar��B��:�`b�⅄s1�K1#���Ď4N�����#6k���],�v�����A��8襽�#�Fr�,ɦ���-�qy���Wë"�W��m�d�83:=������ ['�@����W�@P�X]0�W$��Wt����y��l!�1���"_��"�6e�Vvw��Y����: ��:�dߒ��!	/@O����BzV&7���mH�P/�a��6cK���.b1A����E3�Od���L0�zO�g<ٹ?���J@�j6d_�|�A�eF8�Qސ?��gC�5J�NEG>cZ$�@�ֆB�����R~��J�2g���K�0iC����x���+2l���W���Y�eX���b}Gi�(s���x]�<.)mO9|ْ�73�'�C7��{���lL��SW���>2p���Z�Si�t��I�ɣ2��� 3��R�a�U=����uN4�X���7�qQ����;i��TX�D?G�����4��˜�a����+�2���uy��t��N�iħ|���2l�Z�N$)k��#O�P�p�L��k���{$"�/����޼~A�~�t�Ӟ���i���'((YO��>A^�z�T8?@���/�B 6�"�p�y(=�V����V&  �<���"��ţU'��긧`�
�ߗV=�� 8�sAS��i��pG� ��iZ#�*�+�Xq�G+j��^pj&����u�؋�;?Ԩc����G��?d� ����=���"i9�"���)��-�ë�ǩ>2��{�@ܗ��&I`.�!j����DuVe,jx�C]�����4H+�����`�gV�'�Z�b��d)�@�G��?�>Oõ���Y6:K-S좰��[4ȨZ{q$�z��X�]~�	�fؤm�����.�Y��͓�y�@���5e�$/?[v�k��#@�@�A�n���!W��h�����OY8�K�Q�-��q��t.^?[ޙj���%���hMiE�\:5��$q?6[O�4+��S�ˀ��Α�{G��%'�2B�zJ�-��i�^\�>���ub�3����kN�FQ&25B�vg"��L��������,y��Lc\��0��W�k�!vɂ��" Ef��W���64��]�ZS�a�A��S�?�>��DSm���p�o�h7����1x\~��EN�t�b�ۋy�-�5,*-��	l/�d*�Y�$ �C��\_�-Q�?�]�0�ˆc��m����EN`�R�:;氦k�����6$��I�wa�%Q��\[XP4�P���Vkm ƕ}.�<;'%)������鯒e�y�o:qTT�w����|�g��C
aC5[5+����m2l&R��"�u�J�-�*2�װ ��k*��4!�"m�hꥵ�>1��M�d_��g����(��TQ�nĆ��f��U�"�߰�����m�n#���s�Pȭ�jV�����o:/��-���|�#xz�zPpN4��a�����v5�.����XE��ڂ��n��p�mۦ�����B��r(v
B��o��O��,y��m���p��1,��P�gZI.����̦u;�ɮV;�K�����a0���ր����ӳ~���	V�K�I}�mѲ����R[���6� �H�!��@�ݡ�Ǚ�v���N0���ј9���W��4�3i��i����	�J��>o�	h�\E`R��-P&$���a���;�����;��ǿ�Q|���/R˻�߸U�9`����|'�������N��Y�8�b�M"�KH���Chb�a�b�xhқo����W�VFU�t��k��X��#d�y�ɹ���+{c9T#R��%��hE����� �j���[X��wr�)�����2Z�g$�E�E�Y�7Q(Ř�B$|G��~�C9{�T�qG3���05�=Ǥ�8��p�^����^��y(��e����S��ʾ���a��B��t�q�zȆ����7��g_��p������q���S��=VB,Z�q�gV�y�9�MʫP��;���L���X�:m�;FT,����z\�o�w54*O��G5�f��BW�B��Hz���Lz�u���D�������ñԽ�zO}Ά5L��� �Y��3
EVe�,\o��8�zX�H?�Hn�0e&rR����r$n'�~��%���!�f�W:���v�ru�J��>m?aÏ����5��_w6sb�9cn���7� �����D���Zw+���V�	yԩ����Aހ%�1�? ,��LR�ú:������຅�Ը+��J��Zw�b�A4��&é��8�i�p�d�
JP�Q]�4u�EʙP[���~�$��dvV��[�\,��K��Ϛ��0B�|�eDb�7&�{_�P,������k�NSoP�sy�w_����'�Tv�zm�C�՜�$�^�'��Z��R�lI�0�o�{�����%��s53:3	�VuzF����ѹ<�ax�1������"7߿@��� P��,��Ce)�-�W�3�X�\���>��Z t�*y��r�]�,�����B µ%��`7QPE�����yj+b�h�L��Kf8�� � |�=�����}!�i:\����=���7����=w�ߓ���!{-&�#��Ms�NӨw���.��8J$�/-�8d�&�!�j�q�3�e�2T�n��VSiW�>�ݡ�Cn��T�ү�k)1ɢ6�>�f�Q5^GC唈�A�<����2
|�1�b��!0��>�aJ��J���`E-����ېm��k�ݚƳL@Hͫ?���mFD��W�L��{l�2x��蟅�$Z-.&<SQ�k0��GI�l�9�7�����5����䳮��"m�8�T��������G�l���[�U8�=P����J+Ӛ"h1�{̢�CM��-Y>��!6ц_5B�z~�c��ʁU�E�^��܅���c�"B-�!��5�59������\,[��31���	�-E������zJ��e�g�4�b�N>$�:�	὇]6�O��Z�	�ֈ�&EnEsi��s0(���Չnb���8�|B6�)�h��,Q%��|��_����(Rqlf�뫾T��Ų�TK�������	w3?����D�8~�WX�E珈<0��&��
�k��������N_������.�x@�k'�+|~NZf�y(8�nk�>u��P�9Ba�{� V��gr����jn������<�Za�sYyZ����c�Ď���?��"�5� �bDIxKpbk�\�7V��¯�޲�{��͓�o8�r3_�^��U�&��{�X%ж�c����+�1�*����ô�O}��sN]�7�t>���8�dr8���/���m�U,T̄7�#}�����i��:ʹ�r��[�EĴ��r~�4$	�B(�@�~�6$	@�U�F��8q'�Β�-1t�4�R�@m�7�^yn6�]y ����Z8��"��[}�G�a���dB��X��.�Ð�`�z�