��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0���C	�i��EZ7�=���=;�x/%`�Y������j�Q�T�f��u����:pIC%��w�ٴ�H��:�7獱v��_2������b��� �����Am�7㰯Z�M��P����j�>���tq�v�¹Q����פ2 jp�;�,�'����P$��qW�rL�PP^�T>�j������ڿ����l����I�˪��J!\��@��l�f"Pj��W��[�z&d�����P�=ڸd�l}D2B�ȓ/��W�=U�7�LNI?rw*�i�0��]T$����r�Q>�m��O����E���M�>~Q�9o����Ea�4�ͱ��cZ ���{hia�B�*uHf�8cx[
Eʞ�s� WK����=��jx��rvD\Ң����X��|ǲPv�"����x�a�wҭ���#��z䷣�#MdO$���&l6���ߤ5T���$>���n���5㋚An��+��lO@��r�	g�~��w<� R ��
@���MJ4�K���TS�/�4I&N�~�9���26_�����_cPW�Ŗ8xrw#��{���bYDw�cw	����G�N@e�B�6&_����b�)���سB�h8��#cΤHk�) �N��({q����_�Nf�KM��?z9W=:��S,������!;�E�p��l1�q�@�.��x5��'S"�6J+��9������.��nD`*��ٞ���k�G���c��i/Dl�C��P	C�O�M#���u��xIC��Yͼ���� j��ц����S���0�����!h���`0P+-�)N�T�S���f��=�	���� @�/�C8	�gL�}�`׌g�i���������j��^���uE�o����"��
xI3X7�
^Eꨚ��Q���F���+�A
�%ʄ�dQ�mU�<PF�о��a=$
���҅2%�,ټ�h�����[���^n�����w����R&f�G*A�g�w	a�4�?wSǇ��F�[0>6/i��w��k4n8�S�(I�X3���X"��I�i���٬�`����A�n��KX�Qjr#h�ɬ?�"��R�@B��3����m&yH^f�z�g.�B~8$/��cS_��Q
eG�δ���v�eb�&�=��v��^���;�y_gY��o���F��x�d���DtN�U>.s��@��$"����Y���-R�v�ܛ-�&�"�ay�����mUDi{�Q�g���+2k�}�9���4��z����&����a���\#��m�o�m]6k!̈��>�~�E2o=1�ݹ�	@̅Y.�*D�<��mA�A���a@���z�뮪�u-:Q�7c���]�s&0�5-O��E!�����VR�Gr��	����[�5���s3A�y6W����w�R��?���R��3oxӘ��ౌ:� ��꤁*�I�"�&�ƅ�~(fD�R5o�X�!�|I-[C	���=֫���7��z�W�`�)g(h!���gX�\�?SF|�;'d�HT���W�S�	��kVí?���
V�����<ׇ��´�2}�YG�����aYj�J��Afnf�!&g����;�5����]m�!(�8���[!q�:���5ʯ=�WhAA�d0���ݞP���u3��4�{Q} j�Oyzn�r�e��T4/��F�t�"ݼ]�$w����K6��^�[�ܜLFT� у��,�����Y#�`d�:���d��G(H(���Z�Y؃��R����&���v�܈����;�=�3��{�-<��IҞ�@z��RkQ|x�T�L4�Ò�V��o��'K�8���}�I������z�O�{kOԾ��U��+#�H����)]��d�K�*Mi����T��ƛfd
��/+�x�҈�.n_|�����	@�?r��A�%�`���2%�
�y��֮��9��M���q��
D��_Fy�\W[�Ի�*/'��/VN�C���1��Ȭ�ԭ�x���Z�jr F�S�4�]���x���)�	#H�D���ܨr����W�W@�~�?�@�1�Z��X�j�����b"p�Q�,O�}��~vΟ��2Uߑ}\������u�[�o���i���\��l�͈)�
;HhO�c���{�B,ם�o���<F���P��Gc�F��n������ZTC�T'��/�GItk��H�^�>r�K�����D%��~#�r�_��je�1�������0dJ̡ը8W����Q~��J����6�qPCA���2�.���f�RO,�j�� }����I�@&&��z+��_��FA9ش֤�(|�J	���J*���i���}C�4�i���p�?%�b#A(�p���Y�YJ}"q��{��/92|�'O�^D=G��fGMf��-����F��my�aT<�ެ���Z��0u!��z�4+l��X�^��j�����,|�l@-b=ʕE���F6M�P�_n���G/?r��� R�X���σ0�+=�x�
۹+�&�w��GC�4��r�	�v
t�ԕi�¨��K�W}^��ܳ�_�-ǜ|�Y'q6�����c9t���T�lGB���4K�m�k�^7�0_���e�5!}T��5l��|����W2h%6i�/�0�)
�<�~�$&+��!��!��[��Č�"���0�Bq�_���h��
3��2y���fKZ;�Bٰ|����&.�qg��"~g�y�cG."�e�	(i4C�K^�f=�X�^Q�P]0I��m.�]i����`�!������:������R��@����&^GO�k��ޢ+�������g�;����=yZ�S%\/���{�����b��y��"#YH�^oo���<5�p}i2�H�I:�*����ζ��Hܻ�|y/��ڶ���.#4�ZKNA��c��l[�F���.��h|+-�A���(�L��r��z��动����?���n�k�����]���g�RFW���a�V�n��ÅdI~�t��W}I�ܒ%Y�n���8#�}<�/�%����<��U�y�����F)�(����j�C �~1�S�`ᯝyyyC�yHQ�$�`�#�0�̀��8[�s~��@徱�����>�q�6����ydm�!`��G@B̳��]p�S���u��)�R��q��9�<b������`!���V�4ԦV�������h��G�1~,R,y"!N�k�R���J� B���d�`� PN�?��RL#�( ��GD�(�.*�t�r�����l��t!�<��Y��z8���z�)k�z7�=$2�9\K0Y���Ϙ6�4A$~���\\��'�Yą��z;�
��Ӊі��,��.vҥz}�7���O��Q�T[�:A#��Uޕ�^�z�t��� 9�J̢��Ӽ�$Z3D0�_!��%�nv�EV[��/]7����� ��]��
_�3+�k@ܙ�.D+I4f�S2asQ%p^	��L?i
eYf�R{i-��^v���3�a�h�@k��� ���f}��ƸK�{�Z�.�8ᗖ�Q:�2��J�>��M1cȠ��
}ʿH�sS�FQ�PR�_(��H�}܁�~����'�E n�oS+�d���՚/β5�~��e]�cm^.����w��C��ٹ�Od��^L6W&�|[[��#�������;�{��8��S��@i<���u��ѫk13���W�&����,v%�@�F�m'�Ԟ�T;c�h�Θ��uR�c�ĵEG����{&w0(=��Fh 7��'w��l�x�xį0�m�'�+@�
�@����+��v�dכ#�R=�W����B��:�.��6�]9��D1b`Ni���:�<.�р��
���S�<�r�$m]*������D�K3�N@÷�d7�!{�x��aֿ����W�Tb��T���ɢ�k��-nP�La��$�A��f>�5�h[��@4��O
Z!�B�7�h��������h5
S�1+���+�Y����̟�W�='�����oQo{jAv��$����E��y�7m�!y���)�?j>�s0�zq*/��B�ql�ll+2nC�\t03�KA?BB�����}^#�}h��V~g(
�क���m��,�I�v��>���
����W�����O�@�?�\�:k\\IH𶩭x^}B;�ށ��$�aDWW�w���+�(�&�"q�7Ő;���N奺�sa�1�,;���(_x��#l����W{HM���%���L �����Xcc�.�P?�5y*�.�K��f��7ږ�GNߪV-�O\rQu��w��y8XԘ�s��x9N8����q����=�c�|�ݸ��o�kӺ,٩�ְy�x,`aV��j-�G\t���_8�����O�Aj��e"���C�	�(���O�㑍bzwܲ9�F��Z�AGU,��V
�h^&��Qt�i���%��9�i3��CXk�\.�;�X����Ⰻ.�7��TJ���n�1�'�1@L�)�9�,u���#��!l��W��R�V�ɞ���� )�Dpt��O.*S����%���Bj�x�f���=��$��UC!�ϼ��
A����}>?��@�[zV��Yq���<��(7�T	�Mz`x��t�9D��9|
'�dx�릉����WJ��%2N���!(I�EO3$�L�ֲT��[w�sV���Q���jt/�?��*a��ٯ��
��>	�/r���ɪy
Y� O��r��{�M �6?�Z��=M,�Ў"f�]���� ��?�;��^�4t�������l��t�X�ȷ����Vڗg�aV��ҵ��L��؏#����>veT6�-h�c�;|g�H��'ɳ@�ũa�X&�S��*>oK�[�V��䀈l���m팥6��e7���!�R�_|`�I�s3�Q���K~}�R����4=���L���hIa���u�Q��SCU4rq��f}����@?����!ݟ��;2�m/�E���Bɶ �C+���2P~`�O����6�SL���d7t'����l�vM�m�֭�q&{�ω`D-BKbɰ��(}|̏��2����7لP�*mN�w�V���&�CטQ��7�����l�����=�=����*Y;��� ����X���s�<�]��M �� ���袂'k ��l�Z0�5`�ӎ!xJ��3Y�q�t���Y$QK�]?BP=�D�5�v��""���V��i��ʣ]k��(���H�+�W��3i���V�s��v�3p\h��y��C<�Ö��`�Q�f+>
|K��@Đy�Y'�w�J;��~��Rp~*/6?����f�^p���%��PԊ���M�fb��#O��� dɝ��U2����6�Jl���YbZ�դ��䭌2u�#�����nh��i�:U���+��L��O�5����bhμ��HW������i��8]5��L#��SBu�/�jd��j���Z�P��Q�mx�A�?.�S��*g���ٌ	#'�00���g'26�[��k<:��]7@DK���Gb��Ԩ�v�i+{�n����jV�����"i�aC��ቃ���Ŧ�t�����uv��g��O�&�4����&�R�{�w�R��5$&�{���Xxb+'�Lj��46\6�����©�s򔁎��t�H�U�罛�$��
T��/�#�[���a���k����f��͕(����=d�JΎ�y?��PI�@^3AY�5���O���#y=ԅT�m���q�U��ˀ*��oK�S�r�#�i��E�9��<�nL�;��!��G?�����\�נN@$��^g����0�J�x��Ui�N��ȼO����iIS�4��t4�[>x_����e�n�
� ��c��������[T�Ҏ0z�ԁJ�H��6����Xǹ�e߆�aݴp>��Eu��&�(
ZF�^�7OR�9���>��XEα���
RoUs�� �
	+<ir��TA5s�}Y�������*.�YHi�MN*׮���V�t���_7�)�%a��OT���'�xF�R�j���fd�;u��Q����cx���d�ޒE���s���fq������p]�[!%X�t}��8�e���.�m�|������+A�}��[��⦘<r0��f�l�ӺG�R�BL�*ۛ�y �V���Me��w���{=��
�$�e|	�,�ʾ��ϳ�����^S6�Rԏ��]��\�%�e����8<Sҍ�T�+��_�%�ȱ������:g���������o��$�z>�]���0�Q[�x@S��ԉ9��e�Ud��L���K2�oԭ�V@B]����tr�^�-`(i�\�ܨX1���7��*���e�\���s����3o���
A���$`��y/�>d�¤]F+�Z�W�J���C��S����8�\��H<�vG5C�4�K�P}�(�H��5m1B>�=��D��W�x�5w�vGҭ��=���$\�2����t_��b'H9j݃8�i%h��?pe��,c�x; =/���hkW�')����a�P�� �x������ r8Qd�$�w��'A��Y ���$=>�L@��{��@��⠛
ɜ���O]&��3!Y��-9��br�ic��WR=�نk�
l��*����s�$�g�Q�3?�Ց�}���ڮ����5��6�|�7�`����3E�`��%�i�R�^n���?��
�
��>�g���ǽ!ՙ~I���ܞ��XyX�ӶC��@	�&�����=;� �rt;v�>�.2-�|aQ5@�De�~@V��\��V=�دHiڹ�*�p������"�r���Q��5�#�@�z��99ȅ��d�8U�c�m�N�	��wA�Ƌ�1�a�
X��y�O1��H:�V��R�S}Uˤ�4w2�1���S����j�7:�����0?��HJ?o�v��f�yk�,R0`�u)%����)[bb�̞� !�����?���I���(�a�)��+M�c�(x�bQ��hR�5�{Ѐ _?E 1+�|q�`�r������u0	ʍV���lܓg'���s��v_�R�0V�u+C�	�������R�Y�q�F�_�^��y,Y�rz�ߺND��_z�'E4
�"gx>}g�DW�&B��1�`E˽�U/2�j#^n�j��IÓ�R?���i��d����^�mL��Ob-n}$g���'�i��3Z��Y��״���N,�[GCh�1�@=O8mYQI��gۃ&���ڲC �қ���+����aeƧ"�����唗�$�j���Ic&T��2u$�ɏ�ج��q�e])b8u��|E�ٵY.A����9;E�'���]Mὑ��e��V��V�k���5���V�Z<��ć���0���6pf?w�E��k�v<l��A�I�a( WLy�f"}K�wē��e풋��@_e#κ-k���c�Vv2�ʷc$�j�g����QK����s�m#�ϵ�xdB�~,v%p��7!z_��ZQ/�q�E؍k,z*Lv�x��CSi���^��9�4��ݯ+� K��N����/Z�xE� �����s���T^�,_Zg^�l�6t�W�I�X�����S ����P��M����s��,��?mp�F����|�}��{�ʹ}�B���y��30�b����}����>*|X�����C�&�D�XM�~�á8�W]�ȩ��P@����Ce�Ǚ�;�I�^}���-cb���~�TŅ 빧&+]����-��^�@a(��@шn��.��>s�BB�,v5�V��$��P���RP)F��bȲ�,�^�`Vsr/��X`X�Sխ�1���ǳ��*�����@H%�W�_�� �l�1yDy� >��O5��^��b��O�$MV�
���-�6Z�t�|�� �^־B�� ���̙��z���C����Y���h��!tM	�����-o���.���^�]��ʋl�櫅7���T�� Td���t�x���>F{��FQ�ԣ{�J2s-J�k��*p6P�fTT��Jg�A�
�n��l���]�*C�=�%����?�`���1(����M�cq<c���n�΁�k��M�k�۰,�Ȋ�έ6oq�*�.m�Қ���9*C��R���Ap~�t��ޠ|	]נ��|�3�H��&��6��Ga��"p�rh�j� ��1�́�|���b�³*��z�P0]�Y\)����7qcֲ��� ��>h��B�6&"��C���,�P�#迅�WvB�u���`�����y6�K>{\9a[v>%7��37~��Uq�:Oqd��:����{�4�X����@�ۯ]���l�eS|�=�M��NѷQ���P��<�����u#�/5J�˄�[�p�M��O�wR�g.�|�������&��v�?r�����D%��� �@�>�h����q�#���ŧ��Q6nA�R��w��ע��}�I�� ����! �CT�clA��,y��%�q��X��1�	��I���e�^�'0,����0������M����cR�Q�gK�N����$w- �Im$b���7����`K,��x�,c�AlIaϣ
t
h����YB,J��[��EP=��׌�.гg�dE�01�W�Hr��׵�������
~�����[;��L�Y�:��@'�S@�vIb��/v1�6@���?_�S[t��j����("��I݊C#-���7�gJ�}�u=ۡ�"�WpO-D|庛��%v(�6ۿY�%��t�́�\�LSۙX������8�懷�:�-���j�DƎ� �(� ���k�7^i�^���n�)���~�y���^o|��z����^Nb|���!�~W���A�pw��^����r'��	��7&��V)�w���<v�g����O���qK��h���N�}�U#�D*c����Ȇb ar����^0ZIl��A�M�ډ��]a�:��>Tmm�[���6]''�pk���Po�vԍ}3j��z+�Mj�����q�NV�m:��
�qO�eno2���o�?x�ϙG�`.c	��ٚ#D/�h�K��չ���ס<r�A��H�&Y�>x}=����&ݗ��`�v��k6����A�g�_��F�$3�|��K��Å�M묑��"����}s$ˀ����VŭL{�F�u*�.��S������e�ػ�K��5�+�Ls��r��dUj�!���^]�a;�-#ͣ1S��S�ڻ_�R��x�/1�� �W6o����}sz��FM��@ �/�"��eȝ��D�T���+d@����Q��Y<r
�8�to����+{���QйWŦ�_�{ލ��.8u��I���P&�
�c*l��Ag�%N�/>vS!��J�c$~�i�BKw0PD�r��F��栐��j^d<r�=�w3�{��������j��/�	��,3B�7�L�<?U���=m��iA�(���Z��ۀ�0�F��۪&g�I��iT�tV��
]xsDj�Z����ݯ�a�n�C.��sYz�EJ��T��,���Nq'����v�������mǡ��T���W��%�K�G��,������o3ʦ��?�_ Q�> f[�c�vR�k愝�D����xF�Md`aju�JH�6���E��3�	���پ�
�4߫�����\^4xw04��;�m�z���w=�����1Hȓv����*�,H��/��n�Ȃ�<ͣ��>a��'�@N�DN%{�or V
 �an�\|���[��a��;_�s]�I�-K��i#ɘ��h����K�wQRo�1�%����~�j��dab��<����#�F>����g6�_����g���y���G����(�n��\���/*(��W���dAʉ#GP�i4V��,7�I�'F���8A��1	��g�F^6�HNGGw�k(�Yp!8��� ']��E�@����J���NQ��[�F�~�W�]�͋D]�5@�xw�g�?��hm��!+��T����K4�՞o�XjAō`8�'8D+֭?�sX1P$ˀ��f�,)R