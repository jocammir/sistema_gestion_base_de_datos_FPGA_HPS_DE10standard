��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�*�\�ZF����`���c�"\��/����1�Z�"��<Y�6���JG�ܼw5�Y�.s�%wz�S;Y��,���]�����L��͙v�<H]IB��]:�5dy[��P����O@����6Ա6Gx�=A0�z)���,ڴq�s��y�
`�^0�7���w�$�2�r4e�I�R� ������r���勉/aY��f{�\7�L߬�!3F�z�8��6���Jm5�o�Ttm������ї{Y�U��oN�{ʐ�-�<���[���������L9O���ߟ&k��
��vf�;Pj"e�ԧ�-��j�P�op"]�_9l[.���)�_J&A�H�%,'+N�f���*���N��䠞����>�@ƨ�A5�E�}��4�����}����D�A�ehYOh�}��K
�"�!�wDL����@�Pg�lV<���#���@h��8�|�0:M[*#7x�`�P
Ypf��=1���s��|5W����U��W�/���]2Zމ��i� lt=��5�#S�ZN(JJSN�1� ���+N�UI��$2[J�4O,S<ƗN���56;���IEҭ�Q묓`�Oix@�%&sjJ\�q6:�
TJ�e���n�`�
Py�	�'�!���X2Q�%��O����L�8����vT�� )�K��U���]�2 3�����)�W���g�=��%*)�)�-���ZY�ȼ�!�'��/P����L��{���do�Q����1#1&M���p��)���D&�;��/�S��B���������֠?�ѕ��Rˢ���$�R����O����EF�1����oM˭��*�{��,��˕�y3�P�Ϙ�OV*���o-2(	}#^,2&���V�P[����;z���%��+&�!���W�4mWv����@�-)}$�����F#�6+?uJ�]�ȭ�� �2ӼR�2>�P�t����-�����х���ٱI�MY���]�%vi���@7�GBw��p0-��xBԛ��Q������.�H�+��a�j"��B�$��l�M)3H��qbR�4M�Q��E8��x�����-L��R��u 1����TjN�{UǞr1A�|�z�Kqkv�w�}2�4��aV[�l(#9{KS/�L���򜹌�`���]QQ��g���5e��tL�T�*���䄒?� 9ܑnf(�2ʗe+��v�'|�zE��Z��)͜:D��ML"��H�2��~{=��ֱ�kО�=�d��X%�
i���ZQ��A3rz�`|���i:�Y�eJ��6�+@����r�$�<�Fd���#y���	��"U������z��|��+*�O��K��J��Q�j��%�b%+y��a��3��MZ�6���U~'��� ��>M�F�m���hI�[(�)�$Z���(�N����#S��߸ǭ���A��D�b��u�KB�kԮz�ccɴ�9���dNz�[/����$P�	3���7w4(MzN�fQ,[BE(����.EF��N��9���B� �{X��_.ɨoϳ���䤌y5C� �IO�6n����Jq��(>>L���`�y����Oʈ������mX�U�v GM̊Y��)�J��<�ߟ�3��.���l�U�LΖ0^l�)��?���-�87������/���I-'p@ޒ��a��&~"�7�RA=�p]�Y'S��Ɉd�h��+֊��q�[E��v?�y��0����J��@�,@�� ��]��v�'c7y��S�q2ivn;��&^"I����wwr���'2u�_2&g�X����lh
��1z�/�&qoV��((��puVk#l�"��;Е���╪Ԏ�_C*�����{W�Q�����9U����������d=�g�?3�t�Oi@�����	���˝o-����hc�}�@��L#E����Q��2Ű`�6�MC��v�ͳ�v��ʕt����lS
i	K4ht[��f0:Jz���k��LF+�V|f7��afh�`��~�r�q+���sԪ�cHbx�
�������H����s�U��	�1-ק'w���P`��|dm���ɔ�- jK�����E9x �}{��9r���B�J�V�R���/O�DK���%OM?[�.��Z�UlE-�Ye0 ��6�ؐ��9�0����'y�W(������=���ߔ���+#Bq+3���;b'o���e�ȡD��:S󧻕Ѝ�)�ꨘۯH��':�(��g�ⰿ|�@��U��c����10FƯ�S�ﻦ�=��[���H=�-/�|_��Ag��c��;w+��͇'u�\G�8��08�`RKKШF��w+�S�(a}�슍�b�=�"%������VXt�A�d��#C"�������,��o˕�St��b�(*� ��$B!��=�A_��@�*~Y��xƯ@e�����t<��[�A��jiDb�\�����L��JhU�$��ƹ)�f���lWw^{�9`���,h�e������H���׭ʘ��G�6�y��[������|��J/�{�Qh����j!�<FB��%*��nl��A�eP���%.��^�c���]�qM����)i��P�>�ϪV�������֋ͱ�YWj�Gbt�J|�pccYp/'���(�e�̒� [�g�����d���G��E*���\�Ur~ ^����o�A���ܦ�]���."#$��m����x�zOcWC���i\/�AP!*���`���K@��RX��z�N8[;�,�N@�Y ��"m�s{d��"�F��*5���o�+Ɖi���Y��|m.��ȀH����9C���}��{cn��܀5�a�E���_�gLi:<!��1]
f[��#�{���Gp��x&0�kb���G��|��-��&���a|:�B����zz
4,P���F6��ZR?�V�y/Z��J�$˖%|����I뎚eծKT�݋�Ъ®���+Ă���#��&i��ibe����Fb�˹l�^�{���Ҋ�k�>�\g4��g|�j*��v/ц����MeD2C�Ë}= �B��f�o�P����pX�0�~���q�ú���W�٪��Cc�;>�w��Jq l�˓�gsB����q�mF�$_�9#�k���?��@����ӕ������^�U�f ��6�J[F�:C��.I���	cχ���\�^�<rJ��x̹"��x��@�b��֮�@���7Sh]��,ވ>݀�(��KS��Y6�����&8�ٷCP-=�u�|*���,o��:��=��
#��.+����� ֟��%�Ut����vp���)BC����c���);:7�a1g�P�狺{(����~VR&��4P(ns� *����+����_.�SX]�[���[hf���[r �2H����f��)%�[Y���)jn��@����,��JB��p^i��dp������B�h	s�>9��ĮH}�g���f9��hZ@<�Ub7k�U���̵bxc�wc��p~Le�ԿlG3�Р/{��V��[s_o��K���탻J�rkm��86�6�ž_:X� Þ5P
Z�Rk����i>�|]��"-e�u��-ng+���b`����q�����v��I�N��T�·�S<�8�H�f�a�o���#�+��Yt6���
%|!y9J��Y��|a��c30���#/���mk�P��XwlW�:s$��K�m	�KF����/(�Z0\Wڑ��(���<S�bKR$���U����`1��
�pSg���cٜ~���Lŭ�u0i��xi���M��E1=D;��LT"�Nꯡ�_A�H�ޣ/�G!��j�u�u���	rm���5,>.S�)��Xg�s>��g��,H�U���f����#	�6�7�|\ώ��������}�ؓep���F2�4a�^XU��Y� (O�0�Xb����n˂禆F}g��MU޶���J}�����!�V+��"=`:G�0׹�iQ0@$�?^��c�t�N�:p�5Z�K�8}w�!�5�L'p��N+w�6ن�_H.V�\����|�x2��wZ�1HXJ)=����#N^��x�.
!.�binb�5�����|\�[o� YaĒsZ2���Q�M�+=;�l�6�H&zj����	�O[ߡu��&lׅ7R��T2F�i�ww#�� �T����aD��9��r`����������aR��3���~snJ�N��'Cb��2�L2Z�z:��dÊ \c��qm�%_m����(	���8'��a��?�����y�ċ���/�PI_75����j�+��?u�	"��b8��J�5>�:K̯gÈ@Qs��*	�(�p�#h�5r�\���R~�k{��8SǮ���y�����#�''�'�i����#�>Q���T��Any�T˞�J�{���蝾}��غ����Y��G�Ld��=&B�^���0d�X����M��աh`���a��\M�9�)�i�L�['��Y����P,�e�!��\({����Ov���Qoo�Y鳈�Ƿ8���k�$�ԌF�M���NҸ2�΢?m�̦t�ʫ&�k�*�p�2Ml2�6�[�����٘5�I�m�;1ȿ��'j]�MϘQ��N�i �b�Ǎ�G4G�S�-S�4�X���w�������2>/"�`�5�-��+�� ���vY�t�¹�}3$��'��k�H���B��/)�ӓ0>f�\~��,��VDB-��yߕi�4$ [��A ����B�к���A�h��N��!�%��7�ϡI�ԬݎW�l��QE2�2�����9��F�\��6գ��&�0�g�)��@~2W��A��_��2�1WC^)�UԱ���5R�|�\z	(�aϊ�@���j�y���>�y�2���x��C��*�����8p���.:�$�5�A�(��O %ClB/�U�c�J����ת�*�~��O�p5��zf��>�L=b�ަ��n��_:a)�6�S��m9����Mcv�%�'��s��!�"E^����Yw��v���p�J�F�*�s8��%�e6�$]��Q��a��b����a���b3�g�����yg�R���p�Sű�e���{��~�Q�ha͌1n����t�*!|^�J����|������j�A��>;�<x`�:ߧ�ahiK�T1�^#¼f+��ޖ#�� �<)�j+S)��@V�<�Q��;8�L��E9��i3��e^	7꛸KZ1���E2�cn�P&����6?_G���\1
��p��o�6�l�\ 8������O�~��W�%]�(�=�9g�10 ��.S<5�7a|_��8QM㥙�e���ZQ�:�ݑ�j�i��*�nͧ"�W�)_I�b�,�50�c����m-�{�喫��d.�~��g�E����b�D�Xˌ��N�Nk���50�(� 7����`,��eXU\Կxd��B
G?������"z�3Ҧ�Y���Yb��3"�+���Ϗg8�l�t�{��}�0H>��>rrj�^��M�>�S*�q驸W����= �}*`�G}%%f���2ۖ�$�[������\eŖ���t�6�� ��������vlS_�)�`��<F9�H�K�&��!L��r��<�S~�qY,��tf�T�7W�|�tmF�=�vba���Q�(�jNݶ��V�k̨F��箄�jg��z��^9*�S����f(���w?����<�A��R�@V��
��쫪`!�z��̊N�FF��� [�0/Gk�O»�[Pك�{�'t�T�Ό� Տ��Ђ ��Th�C@L���1�u6G�e������$_����,��4��[盟�N*F�T�\7��S�Nz�t<���4O�H=��VsO��:��,M�����c曂s.lAO]3�T�Jm��S0�?{7);-9&��N��y��'��~�����9�/#hPT��r�L����g&���2`Z|��/�4�N�r)��뤗�)x?0:9�R/G�� d��%j�T�]��ES����~Jy��� j),Am��=��]o���5���{��my�p��苨\�qk��I��ޗ�|C��Sٜ���Jd���Gr_c^�{�D��ܐTF�ⳝ��@���6���Yq��Z�J��@�0!G,_�C ���-��\�SX�s�U�v;H����{�e^�y$�H,;�i��z�~� ����9���� )r
|���R�˂����KLA5ҋ��GoXJ�c�m�s�aY�����r�Lz�ɪ�@!�{*��pL�J�`��ݢD)�.�D�T���
i�o$l��2�����O�c�8��7�s�$�n3���j�v�܁,Y|�B�(�/�tr7�8�����0�e�8<^� �SB��,�&'�s)�[�X��8�sWj��:��W�?M6�������f<�r��L���\�u3z�!c�K�iE{�x�H�7b��aJ���pЄh70m�ES[�#m���Ȼ�Qk�O��ۃ<z�7X*>�N������̒OVk��pJi�c���'?`�@(��W�5jo�,����"�W&~�LrmR���ozǷ�+�M�]�@�WJ����ّfT�i���t܇���$	�l�x�t�6���b�����X
\�oЭ8!�D{$�x����d`L��ގs^9;�������֑�v��ה����6��?���}�E;.�f+�H��V:H��!oG���q�[�g ���W��6�R��i��M/�E�_!���,�j�Yj��3��ూ�e_M������7Bg�) �ܘ'�| ?&O�8w~ՠC}��N��d�f>3r����[X�^��,���iQ���Ƙĺ���E��}�h~k�0x����Vyȁ��9��z�3o���(b[�dD�O�M�a�t�[,yO�Y����}�����N� ����+>������;m�c[��2G�@�G����e�	HZw�l�&��hM�T{%w_��.�۴r|�#>p�=\��q��\�����^mh�Ow�&��X{�5�	�;G����)6��pH��9'��-EX��E[]���O�7�T��d���R7��5�?��S;�����5mb�"�$�@ƈ�;#<��m�m�aQ���k��*G'qf'G��%�]& �Z~tFfz��$����"��F�6K�	�0�}�%3X�h�H6v�B��BŰ�d���QЋWJ�:�2��9��������M�pѾ#����h���㓏� �0~h����"�ڏ����xz�r�A�c�"��4�k�C�x=0]��Yb��� �����C7\
����8A}-*Ѕ�V@���<G�K�VQG�1��s�xt�v�] j�=I� ��	��Mv\<��Տ�g��r�(�@�
=d!����c��V>1�-S4��[�#(N�VH��o���;feY���5���a����n�f�`G������u:����j����$���Sw�G�ѫ��$/~�E{k�ו��m؝'M<���9�y�����v�"�xqK�7��Jީ�M�6�Ȝ����(����"J��Md�H�4�3ִpp����2	\�8�N��BC`�9{s�﷛�{�1q\L����bB�{�aVj�ˁ�s(�a��&wZ�z��oB�a��SG��*g���E؉蕥e��(��l���U���k����i��FdZe��/M8�[\��!�0/+��U+>Q���$o�*گ���C9�͖�ZY|������f ���d�Sz���%��R	`�W&ľ���B]�L܈�]i.Z�T�D�N}mkK2��"�GB9K=��n��t`ܰ��ŭJ��k~K6n�j{-O������r��u�ROqc �p�����>�	Vt����Q�ׯr*{Jzkz�b�^�*0T���i��ή�cqd�"�H�+�d��&
Z1��6Gx�?�5��g�R#
�#� BM��Ղ�U%��,�E�L1ǹ��ϒ�L��������&��y3��3oۂ(��L��^�)���>k��d�)�������D���tL���%��O��s��l�-~�'�4XM�M�;z�N��l��1�5��(��4&�d�Qy��`#��ᮇ��GQ�t�E���;5H�˄��X��SV�Շw0#�C�i�/<J�T�x[`c(U�Rh8�bn�3]τ꺯Q�h��t	w�|����s|Bv8 ��f!�@�;�����2�n�����OJ�g���mP7�E��{*� J愾F 
��E�~8U�����W1⑾�7u*J�[���}�`!�3+��Q=S��uHB����b���C��7�Q�ܩ8��UoZR&ƌDQ�scu�
yS�bT����[@���،��IK��=���'�����������i��� X���c��f"�,���\]ah�VB�8@ �^�]| !M��Фh���"�\sB��[ Su��C��$��n53����AH/�?�9\~�?�sK�s�J[[,W���*I
�`����Ϡ]f�A�_viPN�K� ��3!A�]�;�QDqf�BKUlr �e)�˹�����\��\RD���C�s*���7�f{��1�Ǘ��=����ǩ[�LX�E�ʜ�n?������;9�m먵�/V��w#o��t��DV兜Y0�sn�Zz�k=L���:�|�D�H��&���=�Dp}���Rt�7��"Š��oJdj�`	v��T�es�q(lE9���X$&�k��>!���=v_"ƣ�|��m�QI����%F ~ѝ9���D�X�t��F�)FW��1����L����У}=�v����W�/k�ٛ�f5o*�����cW�L4���Q�^���R<�я��[���0=-;�WD�u��$��w��	��(�'W��{��](p�zq@@JT�'rȭHIaȷ�!ɜ��G���+ �o�eX����]Ie�O�V��ߦ:!c�^���Æ@���2�j#n�P�]��;��"Ƀ���C�V�}m##rWǾ�Q��nT�S>mi��9p:V~U����㖗y�&�˭~���ئ���`���B-�5cK�|���N�(1�GM2����D�a����mh�����
Ǵ�W����w ���I�zy>!gpH���M��ϾU<�`��!�>�vtN7J���*ݦI�X�Ȯ��۫���m�����C�*�0���0Ue�M�)Mh"��n��N&�2�.��i�{l�n�Jo5vm�hJ���PJ� ƅ�PNO��~2�V��FM��*�˙8�:�N~�#%�	4�������w��.eW��Z4�4��5��F������|��
��ЎL&�I�0�
�@Z��dl�F���rvQ��ϡk͆	R/��sBj ��h"��͗s����I/�G�'k�LI�H�E�y�?v�\+&�R��rMʐ�3�΢먹��2�j_�=h� p^�f�I�[԰�j�
�K�wPz+ �mZ�+'^/{%!w�́q��k��D(dZ�B>#�H�(@bn��z��=sr��*n*�����)���H���4�5	�i#���<����H<��I�Q��`�J�&xˮ1��B�O�dBI..6hC���33����6K���7Փ�MU�����-��\6���]��Qh*�`��s�o0�AWq��(���2���{ԕ���oA�;XJ̏p�����֗G~/Ӎ�����d���G�s #�;�}�(U��R��WT���&���f�:�$���2|ZmNri+#u�w[�)_6��O��Ww�����BgeYgDbA|s8�Ks����t��D�!T��k�C����NtR@�����L>�/T���x�y��������ו���+�R�?|
w� �\xe�� ��!�Z$5?��CL�pJ3�����b\��֡��,₶�P2]f6ix��N�Rw6X�/���J/B�n#�����닡��"Z&.$Ў;O�Ӡg�o�`@���c��f#O���5C
)��}�Va��;��,LV����3,��Q���a�!��rM{�����S	I�,tng�����*��w�5����c{�N��6_���K�����|o������\��77��G�CO]��%,�F?�@����7ǌk�?|�(���]3��r�,Y-�MAZ8voTl�?$���t�q�0���{x+�o���J�H�����4qr��DN� ��
x!N;�b�3r�K��>;�G]D
I�������{F��O7x.��^x]'kfG��+�Ĝ��(R����4��Y\���iD�)h�c ��]�������2�&�yV��s�
�O}j?��� i��OMV��sNc϶�:��	E�f���u�w*���Z��T���c���-��_�VjA���cRd���܎x���FXY������'oO�����% �ׯ�F��d�?^()b�"I�FMPT�!"&�_�Q�E=��7%�J,����b&Y_�	2\��Q���u�NoL܁>S�Y����QQ�8|X�(�l��=�3����X��_��Ԗ�]+[B��MO����^�[(���Lz�p!�g�M����B�~yxC�LF40����m5�G��B ����F�\�Kh�4`5��JZj�+��W1T^:K��b����,��|�L�$�6뵪��W��i�W�KG�v1R��	�?���M��Jh`����mЋ3a�D�6��q�")$����Jj�����<({�w��Z6�}�M��_�g�1�.qo�
Q�O1��˪�}���w�@⑥��&���
��ς����+����{P�h�FD�����_#[�R���p��j�1;��,%��.'5��׊��u�awε�|Cxg���$�����Y���)r��N҅<D��<y��2���@ӳ]	��V�����fD�L�TA�N��}���p��#m_���0ei�~��m�1@B�+�_�00�KZ��U�w�I:O�+~E����]u�X�A�HYֽ��A�xݏ:�)y���9H�\��P�[�{9ޅA�VHLD352dF�͊�>������a����S��/s b��L�	G�Y�L*��ݝ���h�Sh�C?4Һ4h1&?+O��hL:y m�[�+����w��2%��;Rgg�|�X�-9U��Og�9 Ȓ�Ğ�=�V�D&8dK��X��1ɄC��Z,���>���G��/�f����؁�I���dhu`��A]��d����K�,�Uv�s�E#���
�Ef`E�alm�l3ws�9� ��]r�>���(5K܌�pX{��t�g�q������c�T�`�^���-��o���a9�Db�����r]�.)e���{�>u�-YR���zc[��h�qj"��Z�*��`
?�X�m�������[�>�Y�yPkYq�7�C�`r:C�m��e�}��k��?�vE_h� �EA/<�LY $�,*~z]7��'C4�j����.��4���Q���L�F��AgUdft�����(�J������+90A�Q+���\pe<�#�������r�F���zw�O�E
�D��ngZ���S�S����M�ݜ@��iB��g�\�X"�t�y�cd�; ��ǷĖç��XUtI/�k�類����	6d:dG#�����1�a�w��I����3K�����A��&N�`�Q(���B�:K�Y�;lX����x�;Ǭ9���dL���FVN�[>�f��y6ª��Uoe���ū���Ӻ���������u尾�>��M�˳G�w�/��ۂ
�%3)7|@킡��z�������I�����H�oU���QVo�!Xka�n,-��]�?w����x��ӊO_����]�L����c������o�i�+(p<z	Sn������ꩥ�Ⱦ���;�eK�b�0s�ǿ�aT;��k�Vg
��R�O	E��r(z�2�.�hq�3":���d�ĵ����{��n��)��Q����.�.G2���Ϊ���I�������ö��x��}k�P��k�AŇ�X�Q^']��!Z�s��#N	�8�^���r�^��B�pj�U�&W%����$&�k&8��e
;�0�i���b�C�Ҫ�ߝk�18*����:��b�?P�:7ў�O����󙜰q��}k'�/�'X�6h�ݼ@�mסEn[U�������)J�i�s���sR+���Nږ�����/�3����n_�xw��C2�ޣ������b�u�����3�$C,ґ�8��2��Vm�1�G�D#Sg���.l.��$��(]��%�o�����Ь+IS����`��h�����C���,��u�ӝ�$�a�uS��yQsU��>譸6�C��3ַ� �Apx��";03���t$��
K���?��f����y�PnA)N�w���J��c$}
l�I_��dP������-E���w?+G�*m�C%˸��n�۳hx�.&�����Dy�r��G��;ş�h0��Xx2V]<m4z?�����w�&��2��׭�8qե��:-S��{�c�h<��w�[�y��Q�ORڹ�M�T�BZc6OV�$\��à���0$ _E�Uٖ3��@c�J�х��y��T�	N�:(��)�U�������/����; &.�έ���} �wԊ{��B���
���-ԕ�F����u�����DW�-�4�Q��=�d���'�G��|�u{$.��>�Z�*@͙�]jB�Zޫ��B�7��.��>� �[���0�t��g���ů��_�ֱ��M^�U>��)ޓ��8��hX�g�I�C�I�.�ph�ݙ��j�8:ꋙ��l�DA�����6�&K)�t�G2;!@�6�b))����Q*�z�N�6�֢׫�0�1tZ.�*�BS�qd4xN���,��w��/#fH{8?��y
9�U}e������~��8��m��
��ٌ�{{_o{��(^e�7b�E�@��o��Yۚ��dզ#(�Tm�����82����!D��t�=����ͺ��{`����0:ع*����v

���C����/��_'���"��7;�����J#jP�\�hzbJ8�T�
mp'�,�	1"�F;_��K
w��x^U/�`b(4�$���y��`�Lڏ!%�uH�}V�#�Z�^�i��&��^�Ujs�s�9QĶ���xui���-b���W��2]�E��Z�#��>���m?	�]�׊�ט~�xe��T*�(��zJ��Hs��%4�y�y�1.��l�(Os��覎a��.ݖ�+�P��MB@�vch>%S����gd��}|�J�v�bp!oP�Lȝ�\�T,��n�z�Z!�p���{���!��=8X�{��3$7�h��c��K�u��߽�I'�4�pC�_��uE����:kg�ž��G��n�f����|i'�UD�����h�,�MP:lO�*g�n�|����n#��B{,(�7Ն��GO�T�8��}����KcME��W��H�,g��"���e_�������J�r�4cC�R�紅�hG����tm(�Eשּׂ�~:���g��L�~�W�ƥޟ��R��!�f?��?��B�qwT1��8��dޮc�g��MKz[}&�-�Abw��uDȡ�R��k��1Pe.���#G��P&��P��my<�pbx�l�܄\��Dh�|�?�*[U��S�-�T�ɣ����8K���t=C��§��U+�7%v-O�[������%�^��A�ȧ'>�cOd������_!�R0 ޑ�p�Mq�A �c苂}&�L<����[h�9$l��~�)Zz{�-R�v�<��A�W��v21Y@��b;F��A�U=|�I�8 N�6Ӟ )�������CA�B�˲�0�N�=�\^���0��O��}h*֡�Eݪ�	���p_��d)f���#�Q5:��0=tHI���k�V�w����Z�&�n�;D��z����������p1��,�������3���E�^�3W5C�S40ғ�	M�e�aC�'æ��� ���!c/yL��.�sznj�Oc��?\��ܐ��K]3PUo+�:��R�?� ��fWD�
�`i�?�Z-�Ow�-У�^���B^�H]�&��x@�kjͯ���k��&���AN۟�[�w=�OvЕb���ǂ�~k�N���=�^�PZ�t�r0�'�� �Ұ�x�o�B_���3����kA��@�7~%�\	XF I��t�;@�ފ�!]���D
�tpH�D�3mT-����I�Z��3����Y��1��ʹ�-����r�(�d�R�V-�9�8��EE��H���m��?a�@oC������]�l��qeW���R|a�o��^��z����Gq:�W[����� ��ȨC���C�����ï�r�-�_(�ة��A!�e�� ��Y�u�NH�汭����+Y��#�l�OoW��-���:}�7����ݥ]�
�"-�(~{~�=�������1oZ�u�J���W$Ʈ�T=�o�v�I.�Y��� i��)��UG�UCh�]���\S�M� �F����݄�C����Iq�&<mS������¥�ll;s�+	�O�!�GOx���K ��!{����!;��_�n��������1L�g.d�XV��9�̻ϛ� /�;�	4�+��Iu3> '5�eJvbl�ͼ]���u�5�`_���lQr�7K��$��S-�k�d��8�ӛ�V ���@S��LO�h�2�C�;�`�<������Q?^�8����]�T���ߐ׃�A<�QcC�܌�83`Ԓ��ZC,�`�Q��sȕt�^@63[�4�_�T2'��L�����S�iӭ�X��������վ��Xtt�1�
~ ���L:fk�F?��_�����w�
���=�.]D��ln졯��כ��J�V��V.�l�i�;k���b6X� _9)��!����$�w,���$]��
�*��h��8n���	�z�ڹ5���ʱp[�eC*��Uţ�(Ԟ\�cxOtU�8;�l�P)��b-w{ӴB^?d*��6���
�4W��!0��0=3���Ϟ,�Pi�Fҡ
f(�"ֽ�����l[u���c�Џ��#� m3|��M,�_�,=�x�1"�x�Z{>Ѥʊ)|X����O�����X���K׶r��OB&����TB�__Pit���u���x}5`Q�/��Flp�Yט��O����+���a�Xqv"V�ߖ�<�FL����\Epߎ8T@R����Z���W�����Њ+��p'_>��+A��u�y�.�N�X�5����%d_
��beV~�X� ���q�ş'0u�w��2� �Y����5>7{�lcT�wn���v�	e�Pi��{tD��`;�k�6�R[�\,��/|
!����i+�޵�8;�a�T�o���)ܡ�NQ%����nC7�Nc��BpZ��\O$h��l{����-�K�;�_�b���&t�p��:"��������ȡ�wYW%����E�k���;�a!�?����;s�E����Ӧ�5@/�$/�k�!��Dy�H�	q09!�zsCG�g�̛=���Z4�o^�O��w�x(���p�z���5ȇ��,�<�QG�p��OD2,Q���|BD��Q�F�?�LcE��<a�ց��p$�}ƪ)ȗ�#%!S�7����N�,4h�g�R�����=�y�5_���X�M�c���=���F1z��4�EE��FQ����Ǧ�Ծ�A@�Ot��Hʜ�t��Y�u!�8.�z��G��ȃ���L�[�ZQz�o�LV��?M�Em���\8�<7�J�р�!^��L	��m/L���~��Մ+k�}2l���~�}��㩌�IR`νU�FX�i��\�lC�@xL9G�Ĺ��Ȫqʄ�T��7�!���񦂡��!�x���;�*��xh�=��L�`�]}��{*��>��m�큖� fJ��?8�Y��=��KV9\�z��ʵ���)���t3nD-��~�D�=D���jD��oO������~nK���G4��iD?	4�J��gH���C�8G˥5���aov�2��M�QL�seWes��U�d��/�F��7=�����?�V���ɥ�hD�33���{m @���Gd��r��� =���T�$B�?� G>A�湼���7$8!޿">��y��}1v�'��W?�b�V�F'�V��咙�[��/}���{_D�WU��A�ɐ�6�����+��;I�����"^�4[�끥'p���3���l�:~{����Z�����^]�����c�vȔ_O�U���[�n�Yò�I\J̮1H��#��
�W��V�ˋQ���dQ�����a��u���J��r�����p��B�{/i��7����<c�-����`�0U���?����h-{�����OU��x���3������] ���4ܡ9(?����o��,�$~`㿟7�'΅��s���~���NU˩4���>uSތ����y�g��w��^�/��d�����	�1��1����zQ����z����Ǳ�ߜ�~
��.�إ�l��A�4��]��aǋaG/���t���U���,�yCf}�ˀ)��-��ƛ��#��ө∁��bjd���D� -5�/Uy�r�亾r��ȴ�����-V^T�u��y�*�H�YE��u���7`1�x�\3�b�;FШ˹\�j|.�T?*/�tA<y�)��{]-���Q2�D|��č��R��p�9��;�^��T6��oZb6Ȏ�͏>At_U��	AsSC����EQ�F���Y���N�:�LM�!�-��֊z���R��͍ �.��
D����05�a� �M�W5�	�a�?��D;h�b�a��m~�r���v�Žc�i�u��(��EV�ة�D�7�S��=:/�i;���l7���#a�n<�~�A�z�@Xg�v�ņR��1��yq�V%�Q,b�{.�tjT��>up��e�;�tfk��.x�
�%���h��a��h�����+��e!,�d#������y8�nϫ|�wf�4ԛ��{0ܡ\3�	#i�v��؞lx�v��.�1�$?��K�̞qB ����L��N��nF>�s�����O+F]��X�v��l�2�P_X��8�-��89����jp�{ȇ�2�簘�`���,���9����!k�2�f���K���~�Z�����u���c?<�F*R�ඒ��?��KU��D��d#�4/2���iy���V��2w���U ���WX�m�ƦVӽ�pF���+���)�g�T��#���k�TOU4ҭ��<���z��^���(c5�#*�P�r���|��t���
8Z�ݎ ~�R�6�v���ղ8? ���Euc�',��J�4�C�K��s5(�A236ך8�JUA���fD��6�C�e��3BgiK���}Om$o���������f*�z�|��&1�j����L	�Lδ��.%b���J��2/+=d��s
�h����i��� ��.�G�	�YG�3?Ͱ��Nz7�J�����g����ꂧ��\�F�fNju�V���a��e�ƹ�&�4�z�-c�3��j"����H������_> α��P#/�]���ki��ao0	 ��oVs�.h��"<���y���.�/S}�3�ۏY�L;߃��+�p��jQ4�B1��W�E}���"R?9�N����A	ݘʩ٩�������4qUmő������٪V��0�sIQ�CO��G_KM/F�@�Ǽ8�{�<�}�5f'�x)ƕ��!���?���d�JjC��8�'L��ۜ�2+S��|G)��Ƒ������.'�7J�SU:�Y��	=c4#��~���]�sD�K�#�,��6�s���"�����Б�$����7�2ZMK��u��a��W{\��w���k�?sB��[G�˛�w��M\r9���ɚ˧��w�M����J8o'[(��Kh�HF���_����L����z_eά-m
�%}�g�cbA*t�Ua�-9E�<�m���?�y��Z�l��ݼ�no�������
�;tQͅ�`�Iۺ��=�|�d�A- sM);�X�R�%�~�{��O��՟�L�� ���m�d���g܏o��N�,� ��e����ݝ���o��h�D�Ox#5�T*/PYn�����-��lg׮�	���0N��*_Hq�<!H��-F��7,C�ȟ�v����b�,�<�.��}w�N9��?�p-��g+U�n���W�=?�HR�K!���`<����iT߰�ŕ_c�{�\��c�8/H��=��X�� �Y]��g-d�Q�c�A�g��%}��U�il����P?��a�� �9����u�4u}A�k9 p�QMV`̆��k`b��hs���4�0�-[�m�>V�
ȡ��0�!��+��d)��!8�rr�>Q�<(�kZ!��|^��.��1^�4���ʂF1V�|/-2?�z��}���tV����S׶���zE� o�mp�������`�m���O�v���Ve�\UX�tn����!�8�_3��-m����^������b6�j�[]���P�c�Pz|�ȩ�U�૟�?��\��s5�ǚ��YQ��:�Ka�ҿ$�Xtfƹ2���Dbc(c�W㭫�Vzc5˦��/�)�;/�!�Q�dr��I�y��C�P���DxX�~q5n>=�,�(��Hs�������g=d+2+��\��^kf�)u.¸}����xe$�4�w�h�i���jv_]�ZC�Q<Cc\%ܶq@	�aW��%Z'��9�3s�D�0E��c�Am</b�����D�Ids�#�g��dġ�����EF�adIf�T�:��4-�}�|�j�w!6AG#-��Č�9��odN�p��f�d���q��9���'6��m ��ĂT�
9���Wv�6X�7�2A�|�iy�z�z8N#�v�О�íTR�>;ۥ�AED��~�q_��Em�k�$��$�,��x�y5|�[���<�i`�`�k��Þ���q8��p���u�姎�sCLKt�e�Q�J��Qħ����fa�;l�Lj'����ҷ5����`�MȄ��A����)����A����~��+eŪ�j�KE�qy{�d7���9�=M��R�t�N�0�(�2�)�j��`)��a0L�C���x�p]��{��z���4����:2\��wA�*��
��A�>���	��=w+V%���Zqol�}�9Uޡ���go����t�J���{{�-iD<k%�o4fϙ�A���F~�-k$���&ο��ם�3�N�_�c�Ap�H��^ȏ�W�}J�d��Au�մ��.�UNHT;�j�ă�0A8N�Yy4m$�;�>�y9�&qAm^	����1!��I����X^ۑ'5�!A�(% f�`�����:��]p����H��.S �#A�
2�A2&��Asԑi��A%G��ӫ2��|��XR9(J��b���A����P��A3/a��P�r$8"��G���a`=�@��ɢib&���7l6�Q蜁+r.	m�9��_D_�vx��*��֓���M�)4m)�pί����j�����	j�s)p��5�K8b'��Ʋ-��}ٞ�:`�+�K׶��w��E^S�%� �����a���v��
�[��Q���D�ѿRLP��N�m�j��$QF���1P4M^ )��e��Y��ZVb�=*v��%�bRs�|��<0j�.�,B�~� ��KJ�����Ȫ$v@�����p�!F@|]����N�A6N�b���f��%k��+o۫w���)�^DA7���QE��#m򿑚�;�n�R��O`��1$0��o(KW!��(:��Л�^r�]N\ƶ�]���#Rzk��
Z��E
G��X�-�ᣧ��E��)$����i��1�Qt�Yv���a����SY�	�t��"������@G�|1����[ME��Y�Z�0_/��$�fە�z������,Z�������2�%��$�P��|���d+t�)�^`���h������0w��K�L6�\�O��r���&ױ8�xc�#+��ܜ�}e@�[��{=�a=�����{iDX*ޮ� �,W�t)7E�0X�Ӝ����h�m�U��E�R._8F3�Juf���Ct&HZ�2.��:2�A��4��E��$=t��:�Ϳ��]��S�h���@�fY�^y��'�p3�r�A��"H<��^��6��b��̢۴��h����59E?�,j�O����?�I��h7�W=W/-�~��䂇>F_�3=�5�m¿�MJ-n#u\�f�x���ɦ����P��q����!�;�G����O���9���w�!sR�E}��׉���u$���#i/�l����%�� �'��>��?��X��h���2��t0��2�w�S��ɱ��1��ڱ�~�	����5;d0�;Z���[o�@F�`���5�ra�ɣ�G%<�J>����~��c+�2�U���|_<����
e2(aP^��6{9M�����E��4eQ�Vlih�d&�;u�����7�����Ud�N0o���-"{Q,�R�
����ȳ��|Tǿ�
c\�Cw�����H#�4�N[x[��Y>��]�`�;��d�,9I�jc�h�����A8�K8��	�tb"o�D�V�c�����s�<��? y��i/f�R���M�?-��Uy�chuwi���R�*�*�1�s 3�B��f�k�bl���<�'T׮�T{N�*P6�j&˝	��Uue��5�r^Ѫ�|?Nb��X��J���l�z,;�隝{��È�ǌ[`1?T��j�0�Ys�,�<Z(*܊� jIҷ�\��l>��[��C�e�j'�����3����K=N�m��R����
y<�O�_I��iް���fI �|B0�0n��튇�n�G�0���Q�Q�^�8=n �����H	�'EI%?�C��Oo7�#%[6��)�2qHl����nʶ9���1��:�N���Ho��ul��)":q}�\���dxV\�����s�_�a�M��ڐGI�C7����*����G͊^�5�V1���v�2��%�zNzlК��F~��4�2�#~�D�E�R��j>]^�Z�Z��rA��(nd�q>�Q�I���������(u��zJ��m9r�'���{�B"���e�_�?�3[�אP�?��M�jLb��"|I���7�F�j�]O�"�s�כr�t��y$�����T`��;I�`!�7�\���#��w�6ӟ�J��
#9Yu���UN���Qk�)Xc�s��GN-��}M/�$5������w8�e�vf��G��RvP6Z������jqXI�F����Tx^MAek���;�Pm!4���Zv���V����8w0�u���`}�$m�5��I�Ї\58S.>T�I�?���&+Ƭ��J�#~-�ֺ�5�8.s���[E���+�~s�4Sz�� ��Q������I�D��{\��P	n7�u'��?���)��� G�ۀ���?ZU�uZ�'��N��O���q��U���A�V�%pǆ8�$�f��ú/3<t`�D��K���%3s�"���3�����|n�X[0Ļ�^T���+ ��F톴amIG񤎘m�e�qr� ���oRM��	n�BPx�f���.�]۟�Y�|��ּk�kL��v%&.�T~���0?�~1y��C�o����Mq8'rm"#nɷ��<$|�j)kou��Q6l.n�P���+�P�
�� F�WL��?��&Ūl�Gꌙ��,ޘ����n���cTJ&c�Ԉ-y��wD8z����Ĵl:*u�܋� Bں��*�%��O�����|<a~/p�iԠ������	s�CS�x!,0�=�O��F��V����@���a���i<�FZ8�	�q��Y�C�,�ހ.o��0�9?�r��ɉ�p�7ι�����'᫬��j��$jaH���O.�!����ʁ��qa��6��r!P}��l���YOu5OGE�kI�t���L5AtJC4�� �	N����:7dT�f˚��ZԂi���s H��ܣ1�d=U>DI��]GoЫ]������N�$|�ၛ���/g���$R��g��X>Y̆�,�ݩ��ZE[k�X� �Y����[�߇�Es"r�H$80�E�b�����[sg�_�^��ҕr�����
�uw�Zÿ�)਌�g ;�F��˥�#O�zc���y�dW]����N�U�R^��5MC�1��p7�N�c�`j,M��.URB��/��g:�����U�S��:K=Ȍ��@wM�1�~!S��d�E�j�ikw| m�b$a�Y[��;/g_�R)��d�lH���!Rʿa�:.ws��vq�d�`��Db8_�w2��)�6V��$�G��K(t�v�4���� �&��䮻��p�_\,��Xg��޺���*
���J��i��>�=�v�u��!+�K&����nt �շ��x�1�T���LgB�epW¸���'|^5�Ճ��!�t�I>���h���g8G��:�@�!!-��Y9;Fq`a�Q�oW�IC�zڂW�V��*!��� ��I����G^��UawUL�g�x5�A7�)i�䤹_�Fy*	��s������Nd9��%͇�`ӪOG���.j���1�}�.;%#:�3h+;N��Rw���]&��g;8-#�B�j�LR�>n ��E�U��4�'���fLR�7��V�k��@�E�M��10ib�	U�e�t��f� M���� r>=�rh���B��q��0���V�2◺iR_8ruV�%�&(J&�6l�N����-�n����նgH��~r�N�d�
�Oj�Qr��rȈ�H�h_E����1M�,hiLcE/o�E �f�
'��e
�5�g��m��[3T?3��ucsSO���4��k��G��-\4^��ѸYL�ti�YN��JQhΩ��k�?[(�MV�>��u7M�����b�"�
��R��.s��gT�hp2�N�
ef�
��m{��J�D�Cy�����2�w}�?G�����O)�߆�>��!Ԣ�a'� ��P���4+�mA+�쌳)�{��i	O���HW�'꘰�J��[���|-^r7���;��]��~auZ[8!"QmM=>�c�+�
�f�l���������+���D�;�֜���!f�U�μe�Y�����*��U���N��6���R��:���;������>j���/=���Y˳:�>�˱e{���F0+�L/P�� �61�3���s��6<��%�� y�����>]��{ؤ��ӏFZ9Ʋ��L&	�T!����ѸM�K����j�x�&��������W��T�!�.}��K��ŝ`66v����k3^��::*��Z>�"]}�ܳ��$�C�vz5A/���6Uա����
��$J򜉟]<d�pm9+�Lu2z�!Z�ڃ�3�]���5[v��G�P������*�B
~:.���C�$y��u�1[�J/<�5�RHF�&.yM��	�cL�~���dv��:���*x,bV�Wd�10�!�V�g���-��;:�^?�㇌>AV4C���~7rx-o6K�~ ��ɖħ�����<BL�*e�U���p��P�̏����8\�~�
)�M�x5�E�V4���<��_9��	 ޹{��IW��hNF��^�a�J�����e.R	L��x�r���%-ӉP�{2Um�7�`/��&E^ %�5�xrp�i���G�
�
� Y=��7G��OO�՟r0��y;q�O#,2��m�l_���ke�Yyph��N�� ���+&��+ ����I�ayd* qI��(�+uu]6Yα:Fb2O��:�~Eܑ>QA.kT��sSZ����(G}�M5����l��)A�Ӡ�6#�E��D�-������	d�+��ʱ��R_��H#����Ȯl
9��+J�G�0�M:��9����j`H���5��E�Z�-M�>|`b�}��
�╜JCa�����у��X���F~W�5ෙ⫻�1���
�g���>�3 ���`� ���Y�L:�V�� �|�]�02�5��&#h��ݳ,|v90��!qh��ؤ3�K/��3)ԕ�c���ͻ�	IH���9r�=�!|zTk2�3�K��萜��qa���/1��c�e�ȱC	��dv!��Hp)�{��"��H,�5?M�Τ�-���W���R�袴Ӡ��J�YH�Ij��q	i07a� >>b<HK/!���.�.���Gx������o�ľ�CC3<����`�F�}�d}�{��Wf�L;cP��sW�ǸW�YK�,��l~5��U��N/)va��w=ֳ�2 �D�������;�\YU��ͬZߌ��W->R��B(���G+��r���[�w�j�p������/�l'|˥Qf��5�:?�k+RF��	��� �V<���V޹g7���̝��(���������Rx�'�/�ΔA�l���X���hJ1���I�{^�{��ҹ����,�ު��(~O��H@\s7��<?5M�|��%B���鲯�i�),��*o\�8F�J��� ��`��+�v��ì���ُ�:j�:@�o�/_d	���,�B��ӊ�G�ZՄ���~�Fi��&ר!'/�]UIΕ#��U�=�v�Ez�C)/���� �:]f)4�"���6d��5�Pp�4P�l"�7D]���-�Y#��K�����G��={����}���#55dI)�������2/�J����;�ɬ��	g���(4	�5-��
O�K�W8x�"��ʌw(9M�OE!?K4�s�4�����͂�v�ES8�����?+f$[; ��)�ܮ�~�$S���_��0�� <�0`��`�3���[/�@�7\t���Y�1���N ˤ���3Cp4Y	�L�TsK%�8�}~�9V3�+U��|(��5�^#X_ ~$��W
L~yql�R8+PR��R�PfV�1��n�/ő+���A�`��(��^�J"�OJ�g$��_6�1n5�mi�[��;ս�b�e��X�����W��}�����t�"?oKK�V���tR.�M"���{U�~��^�=݋�ۭ�)�L����L�T��:�ӔW�y�~ Mv��L,��djR[��Nv�u��Ǯ'"�������Nn��{R���z��4�?��Ԝ��C�
�>>b/�=8�"6�a�t=�d?��}��O�[�H��3=+ n�G9��?G����g �f>�d=Z�������T���L�8�͒@;���#Mۑ����B֡�5�׫�C<���Q`����U{EA�X,S��r����y�&\��?]��1JO,D<I�8���N\R�O�:�Z�]l�f���n������M�3�	�pf3j��'"a�g�(r}�w���	�wtV�u!6yrc栫_�-�9���|8̻$�M��4�$_n�n�6��'(�t�/�H����O���3�L�ә_W�[Q�mƟ���9�'���eǿ
�������Jn(i�r,I��>���B��Z<O�Z�rv(�?�?�5阉R�+�rS!�+�h����\3s,+\���ǝfߒ/������~W���3�!�u�33�I��ҽ�d��>��)S�?RA/��@�	e�8vV:Jj���f�Zkg�#��.���R��M�^Oټ:(�	J�Y6_�-鰾E�P�^�@�GHCۦ;�P����?;��n�yї���	�{ A��:֭�3�Cb1鏍l��(�t������*@�6�?'�h�*Ї����K�~��sϱI"SY#}˛�st�r-
�i�o�`g���3��\p�9UY�%��(��(�.VL/�Qkk��T�%`J����X�a�:��i�����#��D�u)��g"�?���
��YP��{[b�~��#��+*�9�f=;��K�ȧ���a���-�Q��W�3��z�ۣ�w��p��Kx3�<�����˵��⨦��:9.i���d�i�Z��ye_���EɃ��@�3���[b�<�,��ˊ
�E*��/,;�l�E����Иb2�������y��}+I�,��S%�dCl7�.-�I��q�f(�sq�t���%�ӌ�\��@q|��VΑ-GE�YWoѫۤ�rmqr��];H{���qf�2��/.���un?�o�޻4lu�d\��Rm�n��|M�.G�]��S$���{]���n�*�@`a�����BNO��^�;[mK ��[i���'�lѾU3@`���%�BgSf+i`S��"��!D�BY�^Y�\v�ڨ���w����V���t"i]ЀwB����n ,iDe��PY�5.�;�9[0E:`� +!Rֻ�q�
�xnGN$�f����=�:���Ի�Z�"�ΠX��o�b����7H,���UWޥz���z��Թ36�lo�:�;Pՠ�:����fa�E��ą�m���mq��1�!ȿ1Fu�T�d�1�o���'=����	hd������
X�^�[�bZ:D3֦w���'�a�d"������T(���m[{��};+K<!�}�/-	J�#��%a��,���K9+І:����sW
�����i���cv�O�F�$��}e/����4g�9 �.?E�ɩ�õg�f�Ť@B=A�N;���G�Y��Y�֔�䩊tJ�c(�IP�O�=��V����������R����s�a_;g���g�Шϧ+�B�'�G����D'���s�r���W�k�r��N�\���y�͒����� :J�H[!��}����e��K�D��n��j�F�)�Q�s�����b�V�z������`ԍ��ԃ�Β^���1?��JY�NO��k����?�"	=�`����C�3˔�Ӷ�m���f̑����E��!��Z�#�7�� ���M�3�;������Y�{�zM]#T.Ö�Ej;x	��_`2��,6�c}��6��@P��&~��z��8�oK{	E�!�{ ��S��%f�(�)#��')����Ⅺ����&��MbY�h����>9��<kA����.��R�9�qy3����2	\�5@#���P�	�&% �	��;V'��l����)x)p�G/%�`a��ꋆ=8�B�&:N���Q���2(��D�'V��������J)[� b��;j#���*�@�1�9]��L`�-�����? <>�W)TcR9ߎhXE��\P���Pi�wx��w��+�1������z�&.t�ůl�ȡ!�6�yп���o���i1�����6��#�q7w����&�z(�?θ[f���/��p����t�H��,Q&M8�3"kޚG�<�o��
o��o-@e�>�H��&%n{|�<~�q�м���{�A�-&)c9i��POa�Y�,�C�#��t��+'r�x�n�F���N����z1~vX��.��j��D�3�O�w|�җ68�>��ve?�1濻�ǘ�����!��;->36�!�'�L�,�]�/�e���N�����{#ؼS�QPc}���S��$����� �Q ��k.�DS�ǆ���nǴ=�`X�6jRt��3�s�0����eNg���u�թ��"W+�m���0!�� vtFB?t:\Ų	����&��鏪(��7i�L�a�$��p�JU��/jk[�~x��5<��O0��ZA� _�`E�'�#ϻ#6��,5����g�B��_���my�O`K]FɟH�+��:o^��{�0A��v�2��?�ȕ��aU��Z�y7�����А�8�s�Y��P�&��Lg+�R������,-ܗ�l��J3��vY�\q�iQl�۰���|���Z{k����Z��Ӿ��]&��!���E���ϑk̄���"�V����=�Y��PF\m�֢��9�q^92w��S��8ݛ���`"Y|PvZE���4O�"��*� �A���(\�{ф��&���]����>%#��M����e����	@)��=���Q�訑�8��$��W������3N�u#�`Y�BN ����L3��aU����p�Qp\A<�9ף�3�{��_�@=5^%$��:�ⴷ�1l|�ިyv�xK�:��I�f�'�sNQ
)�|9���T�Wu��޺X!�Y/RU�갋�i���S��Ԭ� e�C tte ���j+o1��s�D<@0[��H�6��"�Y*���/#�����w�ZC��N��PƻQL7��ov>�|R���(�sg�a�G	��$��p_�.d�@̺"m/�6����F"`�7�c����R��^ب������*��kPh4�-�؊�3�:�(>W�4&���X��5f������FIG�r���� �-��`�&��w�[���EtgEAF/���LMmB`�=�p����S�&JD;^�6g���#��5��G>�r�#��$m@����t,�Ӆ��L��KDɡ�A��a�g�&Ո�R�]�N8+�^1C0֕�w�xE�b�.<j[+��lխ�(�?v�K�o39���Ve�º��\R�l��2��Y��x_��I��b�$O��U�f��������p2K~]y������1����A,s��4��tG���C�Fw�c}ڕ�?I�am����Fat	���u������
+`�aՁf�&������/L��nxӇ�?���}\N�o�d������z�S��ߡp��G�E&�}� �h����1$�s� ٽ8�������.�f,:���ƫ5��R�r����f��!1��z7�(l;��u����D~ u��W(�Ha
�|ԩ�Q�j�fϮن4j��8Q��9�Gz�7�'�}�7KR��~T��(�b�f ��S,�ŋm^9�l�Z���|�:D*��&N��+pn,axZET<�W�g���8m&T�&hp�)��~�9��U��4�]�;N����+�ۓAd�ý�"u���G�A[j�M���d��5�y��:���j�^�E�8��V�H\��\[6PED�>�I�m�\��/�-���2�џ�.����b���y᣸�ܚ1���p���LwF��r NM�先1uX���&�����H�ϋ�S�kͲSP1k����O�"XZ"v��H�Y�5�)TK���"d�`��� �$lu�@7��q��>�m¨�M��;	�gX_4�0E���C=�Q$K���ɽ*�ӨM���g��*�J�+S$, l�de�笼�L�f?�^���J�lV�� V����W�+�0&4C8�U��{~N�E��dΆh���sEO ���m?�j./Z������Rs:u�"�-��X(W�Y���ې�_R�ш�k�h.n��7T�2�w+4O��خ=�T�"4SX��~�OGl�����?CV��1��Z��V�.����[��aZȓ�|�^���R4�&�G��B��q���HR�d� ���kp��2T�d��S��+�̘Inf4��G��a\�Q�("
K��+�C�{oy>��-b�VA���E�j���npG��$�����$��>�%|*�NleS��u�Q�<����c�]�C�����C���zZ�h��n���6=)�`�cU2x9�ϠO\2�9H�!o�P��{-�h7�~�)j�3
�R	<�j����nc�3�N)����e��۰Z������;O�6�mL5
`{�?�xm_��\�n��P\qQ(�Rf�����*�"C��Ҍ;�cvػ@�Lr�Β�`ӗ�Nyٛ�#�5�(Ʋ~f��\ c�Wq=�N"Jݲ�jCil4I��|Ŝ�*���\C�o��ϋ��PyQ�z�sh�}\l��'�U�j�����(��{�Z�wqr�	�)g��~@o�(��0�pmɝt�}�h:ƣ�}�5s^�������߄&��/�0JԋE~J�������D�{T��g��g	;��� �q�{���
9@�c��y���f�q��MI}e�4(����.�i{�R��"�Kn�rN�����԰�h@�ΨZ�N�$��L	����V3��@�E�5�X�W����r��a$�9Kh2̳]5�k�F'S9���f��i���5��nŭ*+�\N�++H<�6��d�3�HR ��р8EF4ӫ������L���e.(�AfK�# ����#���b�0�&hy�z0JNl��Y��W�}�&��z�e�1Wfqdծ	0}#� �,�+~L^0��Ȁ"���a���+��r�ȳ���;i��+���M����I4&V#��*�I�N�m�|��Jy6�b��W��Mђ8?u;��,����U�$��Ѭ@��*����)��d����&�HVJ�F�p�c��5�$�(��܎�X'=F������f��C�]|3��Ie}Cg�?-��>�O��i�߆��.�`�*�	�[�0��=�����AtUlx��K�w�:��-��p��"'�<;���U�х�~lkR�KYcK}#�c8F2�pO�K�]PYiJ��.�x����C��(����%
��͹�Kb���D��b	:x~_n�1�QD3����46EԼ��)���\��r�e�t�Ԃ ����)��l�2+�evrF0��=��k���j(�f1�Q�8WԖ����#E�E܃��
1��
��y��{э��\���u��: ���F�h��/(w0:�v��$��q��1~Mo�b�jk-+E!��%x>𳛛�̲�6�v�,�΂eD�|4}�Ow�7y$�������p1�;��z9'�Y���c��#@��t���jV��w��l���=m�1P�dF��N����
��Ǌ�TAZ%����bm8m�l��j�Zb�L:x3����xd�wy�b[.7�����ґ��;��	�h�oD,���'��DȰ����ne1	P��ir0Y�/l���AM�;X��3hG�����>z�WiU�r,���,rn:N��A=Q���-��	��!{�;�j�^y�h�>�^V�:Z���QȐ(@���s�8}LO��1������+���Nm���6����BW6����~(��V��f �����#@1���Dɬ�Y����pe�Tj�Vf�(%��M�R!�݈r�ʆ��nH�!�~/Ȝ@��TYU���4�W ��,+e��t�]&�sx�Y�ŧ+����y��S���Oſ�~�7��
q�#6ꝋ��8���x9����3�d�Ӽk���ҧ1ل� ��epќ.�=�3$�FhMlA�ư�(�G
�.�k��k��HHX��T}�3᢮మF۾\L �&ľ9wǳKJTޤ$��&��t�|�F6��z2l�����4�r�<i�
����㗐0'��|-8�IL����W� �3�����S�K:-��D-����)�p�x���ҧp�\���U-���z���]@D��Fr:v	����> dS��)�\O�#�\u�D�+|�kK�Ӻ�:\Ĳt �)��Zv�����vqpYz�u*7 � ^7.�-�CU�--k�Upj��3�H1As�_�+�+��ʒ-K�'6�E�`=sZ1��&��!!g�'Dn�5���0���]�8A�u�ڭ�ؚoM�q�IB�W�F���*|�̇5��z��- ґ�ѷUQ����n�a8
3��D�1��T?bM�����]�+��0�^<sٷ�ʀ�;�A�+�� �o�g*QiVQ@�����Jx�L3|W��U��2��)�&fDL��[�^�����1c�h8'hw�M��D'����z锷"p�o��q�:.���LOƴ�^�I�,�h���(�mtr�e�޻��W���$�բ��e�\3�J�;�#��\�:�����"J��7"W(��e�q$y�FyO����G�H��~ �x,ʗB_z+T�&ā
�P�%��}��TN���Y��H�;�yXC_���Ş�S��F'���;��-�ƈgoQZFV��d��Ӷ\e6+U8�@
Ͻ�X �����9+�$��¿o!d��B�w�!J�����g������3"�!o�@�bA��O���*&����A���ӏ�k	����ɸ���8��AA���R�CNN�6&l�O����?���d~����sq���Gu#�zt�ξA��2��v{-�C�Fz�y�3��6#(h�TEAk���5�jT�p�1�i�R
� �+�>��K�紐@��f��m�4��*_��Ќ}xᐮ:�\�A<^��rByU� �p�<d�*�c�5F�byx��֬+�n�VM'e�*���s3�:�#�*�]��6�f�L4)�?$������vo֭�U}�x��{�u��0c�/��&���J�,��P�U��:�<>�v2b)9���7I!�?�g6H��e�q	$m�œ2飙�%1K�s��Z���	�ǂ5���/�/�5W��
�]�䅂���RɅF#��YM�Ԓ��3��r�Q�9����78Pq� �>A���W�X�J�goÂ:#RO�w�n����E�*V娐�6��WVcse�<�X�L*k	����9�>*���u��7�Hl��P�-A��'ׯFalkp���ld�[���J6��N��n��C�B���^����7V?���_���f�}4� ������sㄗA��I�D9�tu6w_C�G\++*A�_6,�w`1{��=s0��?W���{���r��hU�LX����4�V\�AT��nA/C�!�0( �(װ����%	�	�
��)hA�L�ƾ�3w���*�ښ	y���@��o�Kխ�K�ѣ~$h��M1��-�x��P����
05�Hz~G�����5~ʤ�Q�QkGĢ���=��tx`� �`��ֽE��"3D�V|*TS��H_hD'�ڹg�'_�x�!�В��MY��գ�:��ه�|pǻ�B��_!�b�����gBx�WVE'�|_�, |�F�%��bb��"4� �(tP<zNI��'b]����,~�#��P����3�/�u��)4��ϳ�*�:6�M`�<���as�|�	��0�q��>o1o����2��N�D�F�!&���!�P�$�K���؜ӗ����ؔu�!чuxv�700�Up��ȤaZgt>�?�o�ܿ�ޠ�#��Q{���S�r���R������!,玙��R�r힔C�C���{�ۡ���������hoP����
�剓��8¯�%�)��%Qٛ#�R�C���o��>�||W� 9���� ����/̏w�%H�Ճ$��;��щ?�2<,��]�V*�_�#.�,[�����Es�:��2���m�����$\;��x81̫|��d�0����p���wf���t����&�@��U��*��$�n�*�
��Щ��iǓƴ�M}~$�!v�խ���Y���~O�8�\�����
���^�+�/{���\�S�A(\���F�����kƙ;�G�+Pg�!�����$gPo7�҂����k���c�A9^S+���n���3���a3�7�3]�����;��[��Me����\Z^=�lұ�ߞg��U���E��e�E��U���SP��(\o�$�BXl�!g��TA����, �<g��s����z�Q���ݍ��Asp�^*J���
��Km.�עA>��=��<��!���1S\a��ڥ��X��=zE%��k��v��e+�e[�h�{]'�����R�PE�* �Pw��]�}�_���I]V�p#V����r����zi/��cx�1����f�v!%>	Q)�4Ĩ4 2hM�#'�������\g�*��7�%��>h_�篌K-��ru��N_Րn_�n�Q���&#�ц 3M��V�,���"rUY㽥�������J���dg�w0qM!+W�o��"�R��^��j�i���/���i�?�=��kM��&�(�`�7��L�"�;�!���H��r��/s�i�;��>�2����<�b�n��i8ؠ�Wb36�z�
��`�~�]�ߝn��Q����'<�g_�xp��[i��G�*�<Q����o;��t]�fP�<І��POQԜ��T|.lC'�������l��t��W�^�T��GMeM�q��Ɯ����P%�\���ǀ���v�Z,!_���o	·�z]V�T"�Ey���� 7�>Z6��6�4c���C�u�F��y����O��D��hn��xH�cV�7�� �|�<�J��bk5�Z�x�,�7���<����=�6�>/��B�h��i0�{L2/3&�*��;}��&����_�2-:n4B{Rh��������m@ڱ�ün�N�3��Ak ޘ�U{|�w����0r�I��f�x����bP
�t���A�ٰ��N�m�zh�gl%���������'.�6��ʂ5��2*9��[j�g��2�y�ѷ^^U���F�䬑n��O`�V��ȯ���)I��d��[���4�|�+:�êLd�q���.{��Q<�P��u]�V;��>ծ�U���kZ�Ojt��NG�_y��LB��њ��Q�v�&@Re@���#l*�p�R�;������w�TΤrcz�/���0�g���!J1z��U��B����d�~>�=!���5�����Oٗ;����%���.��*�/! ������5Z�}=��ޓ�ҫ3��kNM���r;<�Mӽ�ypY�� lW^�#�'U�R�p���
��<��B��~4�L�H�.|�K�?�f7R��#tePRcs�֧�m��m�BP �h��t�8��5�;�I����{�5@�������5���0�C��"Cʭ�{�����A��O���fmO���-Ǒ�i�s� k�쓓Ne�Ř@:�x�ޟ?��6� �[J�l` ��y����� CC�.���8P	��K��o�=����<z����=�$������p�D��l��AȤ��6�d�&�l6�;B��s�g	CO��a�Lm�\�W&��SY�~��5�1s�&?yvz���}̿4jG3}��r=H�5�+p�*)�	�c.�g+9+�c��������R�uQ�*WelM=K��门9�G��(Q��
!����m)9�����d�	�64�[�n�9֟�E�V�׏B_��f���L<�ڟa�!�j6�NS@�ۖ��Eˑ��&y�����a��-l^�vx��=I���t�	�o�f�w�c��1���؛�c��+��j���x���Y{ ��G%��w�:��f �Y��UH�
3@�;b�)'g#ׅ&��G���U�Ţ��CQ�/�7�y�/�A�{'���
��U�O�	�8ܲSKf�Q���ǻa�5�����Y�� �l�m2��u4)&.n�m�?'��z<��	�ާm��M����T\�I��@I=�CX(u�b���2���(�ZK��l=������
�z8�OF^�_y$<�.�&���V|e�D&����)��ʞX�ԜÎ�n1�#�!��1\nV�%���n!�� CE��ߜ���-\K.���?]���u�
f�S(���22���Z���/	�tI� �rj��2���I�:����(��E���㪢���{��h����bT��j��g'�/f�sf٪YV��q��X	'&� '�c^��Ԡ����j/UO�>���p��K ��}7�ʶ�<��PJ�����n�C�-�n��w �d��u�0����N��C!p2���]��B�YO����e2Y1��v+���t$ň_�&)�p�dG��jL� ٝG�N��ʉ>5�;ͦ���jg�R�_�������� �9��cLO'6���_0Gm�5��Q��w*�[a�Di��>���"}A����@��04�Ol�/�ə����V� K^�\5�>��K�k\涐1�P欏i��ŀ�%�7�I'����=�Ӻ󒵄�Sa�V��@�~(a�Z^��>���6I
�s	�̺���v�	'"�=��_�3)l4���	r48���3}`��	T�E߅Q����Mh���������?�A��X��C��� �zE��D(��޳��x��Ϭ���X18���������l-�U�¨�i��ʷ}�,:�^�3�����b(�V�m��T39�?Du�Lh�(�b����:�`�R��ol�yBT�k�!u,��U3 �:MSԝ�F"G�Uӷ���KlA�Ȋ��m�K=��ѻW�mQ��i���Vi�m�m��t�ֈD��g�4�3Y{�?ܸFW��>֢�k;��OI#�毺(, ��
~���C���"��F��
1{q�9��!R�����	 	��&k��8��[��x[?��ѭ��]���n�Bт��g{�Wpd��/�����s��~$�^S�j���.�	��9|�y�G�N�֚��0���qU��E�*��CX(����V~~Y����R�f͗v��?!����^��N���8*I%�gt��-é6m|���T���ko����|ʵ
�jG����L�1ۼ�x���+�\��8y�rw©><{�����~e|���p�%��[qZ�����9E��w�9��VL���R�ҋi0&2؊�w �]�}ً3��D��N����%d �����D�i(�[D�Ê}w}�^CÚsu���)�,������-\��>*29�$�6H~���}�eS���ǧ@�`��2(���y�Gb"T��{����,��
j����>� ؙ�]Z�wf_��E�mF����������/ؚ?�|U���/0�h�֤@���9�yba]pF�R�(��
�g��T�R<���3�]p'I �Z%�S�=]`��h3�m��`�����[�_6��D!�o���Q/��/~$�j�"�h�o�ه��,�'2d?!�Y���1C��y��`}x�>~s�Aͱ	��E^�vP�-L�Ӵ��K	v���u'����/O��N��b
��^T8�z ���� jS��V}
��.qInTߣe�At-f�]t�vl>�$+�hnu��Q�+}��P�f��
ptպğ]�hvZ
���[��V�K�,�H��A��
�����*7��m��$��Hl�\z����{F"Tsj�5qYJ��!u��#�+�\v;Kg��ƕj��E�2^+��0A��.la�2��۪K���-{`n�72�}l#��~g]4��X�U���xO�	N���4��[p�c�R� ө4C�@�/'����8�EI��p��T��j��7=��
k�=/�Hl��r%�h#m�:1�n o\�j��?�2(i@ogޚ3�x���d�3?|$M,X3�Ŗ-�ʴUk��R���K_"�����n������ma�.�Tǻ��6W����R�1d�>��R���Ȁ��8����;)98�r <Y˷�����G�9�_�����E*���[�VO�*c#�3�?���f@�Տ��UG�W{Xۭ,���>�@�~��X�<�0'�?'�o�1�Ht��h��YMl'h�����q�ľb;875�13ٴ�P^
1S�B�vЛ��4�$� ^sUj�w��i�Pv 틶����U���[������aۦ�d�q7֤��x�^|�����'_#�ۚ�Љ�8�d��A�LۂrUM�����Q���|B���<Ƒ��8�n-�t+	s����3�#�v����`��{�/��Q��e����>N��o���g�t^a����*oj�uz=^"0V|Ԇ9J�?���'�k�,��y����kD��X[6Np�"#�|}h���rG��M��+ 8i\-݂\��
��5���;�I����W��^�������9�'\�b�\�N�s�*� �@^{����d���?�"�ipi��\���(�,��Ph��	�r� 8����:���ۂL�M�baH}��9���Z(	�֜ve�����f�H*��2^�l�po4}8FھN�������ڟ�+���DU�g��d%?���||��3@�̷#2��Xh8������;N�yu�ᇁ���ΥH�{(
�%��W �S���n!-�6�Y�*t��E9� �\�x�[}! 2�M����/�q� �~7lՌ��Q�����3D|�l�]��y�bxzD�&��:3�G�u�&���y6���^>��懁��Q�m0�N4�wpAG����FkW�L�ՙ�R2Wf,�b5�*�f��yL�/HLS^�����	%�9F1)QQ��4X�1�NO 9�ಣK�ke� �mA|?=h>��S	�CJ�+� ���8[	,0Oa|����F�2�|{a
�{�K��*�0U�&����ݻ���)��iT:��<���%[�b�%�������2����6�|�ۂ	�����n��)��)L,�k�Ʋ���Q#N�S���^&rLc
7�E�^4q���h���Qq{�Ҷ�Yw����Gt���8u�f�g�2��dZ�/ﳀ��B��Mv-N+��T��ܦ#^��SQ尵�AldF����'f�a���� �i#��C�A��6�M�-4�Y���S��{����V��&�+��x=O�+\�X�usz�^M�h^�5%�/p�H�\PO<�PwJN�)"���� �Kǒ�:�9x@�1�N���\�ض���#3CK;������p�~e���'s�B(��q|��O���#�����2��d��"Ƥ�>���	)_6�/�lܴ�EF�a?a���ݝP�p�kT:d�G���<9��DY�=��װĤ������{Xw��-�|�����_�z�Џ�~P.l �PO[�g�'Ew5���I��ߋN�G���SA�"�|¢�8��zx%W�N�zݵ��_�:�jnà���M	�U��� ����ʴ$�˕!�`>���ܶ��O8�f��z�rf���MH+��w1������uc��<�/�G�3i���гDΞ9Ԫm;�gR����-d��f˿c߷�1̲���(�I�r.�w���D"������{�RA-�r�� ����-TF����#�-"�Y�k����liF��Se�\qL'�W�h�_X�*��W��--vW�/$	c+$��=���� "=޿�F1X�eJ@�=8��$�T�4���֬*�zD��B@�J~��IW��R��R-m��O
.�1��V��͸��D��"�_5�1Φ��,��ȳ2��
�VQ�w�(3��� r�,X�V}<g���yBoI�D"�N�9�^�����V�n:a�";�L���Bz)�#B�=b��*t�$�5���Q�����U�,���V�"�q�g�Þޔ؊ȺبڮK�0lk��۵�.���>�t�w��RSI�'�4EХy�7شH��W�F�7���-=��p� �@+���8����dX[���_'t�IJ�������X%�jJ�o6��(���v+?cR.���H&��u�{�0����r��G@Y��9��!��n#�LN�$��&Kh�"虓7jl[�F�G'6�kA���z��p--hUU�}~+����N����Xd�E\�����|/�K��mگ"�ZB�*�O�-C��q�)�rv
�u��uߐb�3T? �1
S��ͻ+�6�B�Vΰ( �g!Gf]
���c>>�|6�	J�lv��$Yv!���%�!�?d��L:�6[�?���a���,��M�D��+�LWP)U�hVF(=�ǎod�P)-��W�l�yɳ9�s2��*�p����y~z�X�M")m~ĕ��y��'Z׊$���|��32����Q��3Ns�MY��W:��&�O2����#1o�/ox��2d�oW܆�W��/Һ�	�4S���r�3���L�L~as�R&�kv�.��3�9��J%i�JN>!Hy�i!y�̺T0i������,&lܢ� ��Yẹ���{��"Cƚ��$u�&����V��E�xb�F9�_Q�0���"8Z����6��<|�~��e<��_�/�z-BK!��裛�*Gm*��A|=�-!���z��ޕ���v;x�4T�_cCM�h�%|t�i�42��<Xl,W��9�a!a`����T�ɣ�}^f:¢�\k��Ӥ�~�@s&��ؤ.y�;�Nf8��ʯEE^/�y�����ç� 
�
Oى�_���͐Bx���e~R��8������gl���f��T��W��/�<�١������N��>qM�d�B+��#�\�7�gξ�,��d�[<�f�$=+�ѫ����"B�mYj�ר����9"�=i]h�/��$��q���.v��>b��~�],��\�Nx�kT��f�[8�gٵ�?@� u��o�� �D��"��b-pw������c5���i���;��P/Fȃ#$���7K�U|B���H���N9���ş~�^�=	n�!ŋ0h�@ޗ�7��1;9�ʐ ��3�S(M�
%��b�\�߱��.��gU�Vg�e���9šʙ)�����7�� Ĉ�;NV�!�C� %�}���kV�ǓjO��؃Ƴ��ğ�p{A����Q�8U9.�s��+IW���;�~�����|��	���"�@��sC.�d��p���c�.Pg]���V�ƴT����"���ϑ�T�j�xu��Qbۅ�A@Ŵ�\XOK��`�d*V��T7�����U�FH�v��m3��܊�m���A�C|��TSJ��ћ��D�]j�qd4AxA�ډ-���#%K%%�4,�����hW@5ѹ��3�DWǅ�r�7%��0|	`L��N����o.K��p�k]BL��]d�B71��q�l\͑R~�E�����OB+�|�;G�� ��G~���C"�0f>��1�Ɏ���j��ª��u	6��g�99�*w�N����%:%�`B��~�ʞ|�{А7��J�n�0b�[s�JUSf�Ļ��=?4�Ǜ��awK��("�!���B��/�mv���f6�������
��5��ڷgpt�+�������x]W�J�_Q>
�!�C�	/����6���GB{�N��t�c��+�Q��x��Qs��� c�q��LU�{xX�}�|A)\E���<Nӻ�8���lYE%��ځ~��t=��i���V��3�,g�][�S���y!��g�a[ǉi�X��j)����TŇ�i�ԯ�ҳ�Q;�����  י:���~�橁������f�t0�� �l%?B-�b�sfN+�`͜�ȋ������oS�[�Kw"h8�9���i��&�Ί��O�x���/&~�	����&b՜�F�'�v[M��&da��Z�,���"�:>����q���+���7�|�FǴ��Y��>D-�l&��ߩ�)���U!�.�TG���PV+�T<�0����'x�\��=����}���R�p�8���f�E��k42��W�x�$n�&�ݙ[���rы+����n�5*Vٮ1BB&�V��/��[R,�3s�#ۺ kxv/O/���Z������J='�����6G��K��L҄��~y3�M��Oj���a���?�όz�{tk]YS'��-;�\�[E(ؽ#%�;Tq��B�I�%d�ei!O��+�23��k
O�wW�W�YH5�Z7rN�K�[��ǩ����F��(�+��';�o��I�_(��|����ײ��s���R���� :$�Ǻr�����/ƙv\-��6��t4����z�` BE��+;���fC��N$�7�X����z��<h|x���*$s> 3���aʔљ��4&��8��!�`�����=f	4�44�'f�o���%���2;2�����~��Rge�2� x�ϟ�]��T�N7���~!9E�:��X;G:�I���G r��PN� Mˡ�b&�(�d��7DM>
ؾ%���c�Z��Tu���>q�
p�����q��Rҷ��*qq���������W�a��b�q�A��Dѕ�!��r������w ������+*��@��̦X���ol�ь��Ws&��v�/�� &Y�<[�N�8�)*��=�ɴ��"�I�./5���f��y �~��-5hD��γ�}Ё�=_�#�1t ��:r`+!V�dO<mW<E[%U��y�I/P"Q�G<�62 �vM����G�ن�m�R��Y��`=�x����� g~��ӌN,m�/���9G�UPh6]2��|���yy{��Oi���x��0e��QH;��9��!4!1�����7�o�t�d��An\�q\�g��RR��jl���Q�z2�C7���fN�?^��i �j&	&�W�1ʐz�����7�����!]<L������ׄ}��O6n �u���(���l�j(��I���yn��R@�b�.P5{���i�A@9�+-���L��*$V���$�Ӽ 䃦�<����(C�ɅKG�O�ݑ�����w��H.���R#!^N���o:4�1���Z������:���I�	��#�:�4�O��ϻ:�~<���iy���
Ng�w�Uq�j�q��g�4_����k��`[Жsl[�g|	����m�}[�v�Rsѽo��k��s��@�9��Q�P����xM��r"P�����#P_y���/_�hxu<b�R��
���U'�Q#Ak|0���4��Ex7x
��͓O�AmLf��mC��s��d �QK���V(	2�#���2h2��U��+�XUn~eRT��W�di��zÊ�l=�X�:!w��+}$!>�{q�qEO�;���/�s�I?��
����9�����
�⸠uq�C�t4��}�$	�M�3�q󋙙v)���E��kwz��q"�wrCoĄ�mz�C~V��1$8�eʹ���z�o��Ӌ�(�WP|!V
?5�z�w]yŒ��*&̊�jy�rA�6� �Ϳ�='(��VwN�!&������`o� ���ڃ�#�� 1(�����c8�aXI���d2����9��7�X&��T��Џ�v�s�!X#5�>����E�	�ܿ��I�x���a�/�d�(u�l��@��J���Co7�T�[�K+,�az�[V[P7<fP
uc�j��C�S�.58�g5�;�����2���h8S�V�Ý��-^�����UD'�m�g���7����cX���T{`}�`��5�@Kq���jb9ɟ����[C�u�����s��Wa^�>��/�/c�0������崮N�
"�d Ꮢ2���6�N�l��V��("Ek�� Và�y�	���q$2�+!���q=���S|�.ʭ7�10���t坿�*�+RǙ�S̙�����4��W����J�(B*�MX���]�����ϗi읮x��F�"k��']		� �:�+�ДA�U��!v k���Ÿ��֏t�!�1"�歕��������bs0�c��*a��z��l��д�4w{%(x
�窇@�i���F��R�}�c�>	� ��o��#�O�H�ҧB�(.��z$>cjT�e�b�a�$Ox'���*���Q��\>wn���͐���]�� M�@\%�G�!&���x�"*;l7��g���wQ�`��[��F���rø7L���%����\¨a4׾Z�Y���+A����;k5C�7\�xb��H����vX�W˟G�r���)E�����bd�m�
�&t7-׉�Ā	���"���\vn��*�y�����+����g��/��f�pTy�a3H��:�X�Gqm���4�� ��ўÀw��������f��{�Γ�G�2�Lw�xË�������N���^>�F�҄=ZER�z�.q����̂Rْ��G	g ��L���^�����"<�!��CR�����������w9���U�o�����#�j�ۨr5O;
{U�z��G�����R�J(��?{#�ج��G�/jN��;�`���ܗt��d���[��$\�Ѧ���[ �'}�nwR���b�Y�~p��7-~�C�	?�<:�u���+�������a���<흅z��L@�WO���<x\ �uxS�:_~�Z�S,�+E�Z�� HQ���L5�J�S���e..�;���Bv)������<y,V�sP�BEʲ��<@�i�Cͣssyt��@8�e �P$tx|���꧶�c7P
� ���"I�'ܑs�RG�j����R�	Y:W��06�tl��֎[�y�[΀9�$� ��_�1�[M�ofo&< O�d.��c��O�97N�� �rl� w��/j�kC�]p�."D6��'���Ah���|��(���|k���h��U�2S.���9*��a�{��֗��F���v1%ðŵ@=	U�z����)�%B����B�����)��Z���L�%V�hE�{s�{)������FV�C	~�Q��T�gy
��n��*5tG�.pFH��KLv��7����N[�Q� �{��Hcb�{�$��w�c�W��);�N8a�-���I-E��;� q7t�i�����mn�|�!���4����1P�;��9�����W4]��OO�	� \wW�&�.E@�Ta�t�!�ދ��>�K.R�!�uq���M2(�`t#���W�r4���B���e�x��{����n�M��t��%��)���2��'��H�εd2P�ʁL��(�mO��ϯ;�h�P�$�眔(ea�����`�' 8ֲ������#G/��Ŀm�Ų�@#���/�3�yv g�!����xid⊣�܆=g9�{�*�y*�8��1����g��;�\W-U�|Ң�Dp�M�]╰��d�.c���I!�(��G�,�0�n ��P�/���@IE ���dz4����H�Ρu��o	����r��W?���1�}Ե%\n)�<ø�	�eF�' ��r?��.p6�K��i	�.�O\a�0o���17Z�%���
Ŝ�8��9`&�{�(=
�
�B��(�W�UG�e���S]F��o˃�3yk�ѧ�a�J0�::Q��vL����fL�����	n�ƍG�cS׺��rQ������ ^R
�K���.Y��s��D�e��#�O�!���T�ZA2-?�A�]�-��/�F�Sr����$��.��� D�{����F񹘱��k���\�m.�G��mH*~��7%Y��ꬫ���ecp��9�7�)Q��v2MH�j��`q�%^��N���(a�ѫ�~֋�W:Y&�L��Fj����A�%h
��qWXg�+�x\��{������ȭ�z����N�/!7���O��ӄ�$ɨ�)�
�=��@Տ��f������ʶ)A�d\��2�һԠ�$zz�}���?��*0$�yA�#��7�.��M3�o�,�:��.��:W)}��p7�?dVWI�n̍��sC�\r�����4> [�z$�VAَ�4��nG���ut��\��:ۛ��㯔�9���д9>em���]�!NX)��:�5dvH��������@�i��u=}�7�O��R�S�%	������.-Kq`�o��g�:<��Ii
a#�y�7㹕��IB������7G}��d�N���B�Ea�7����s������Z8"s�\���a�c;D��S�([�I���'UL����Ξ�j}^J��г�"+Z@	G �bE���/Ew���j�l�]U����A���zh�Z�CȞf��2Ϯ�qZeBM�!�Nf�<06���l>ŏT��6���_�fl�PL*�}���ZCF_�لDo�o�·BV�ki<�?�b��on�o�O�{�N�a+pĽY�0�o<��5op8;�W��bF�I:�����2�-Jm�?3�S�WA�qlWfE_����m ���Y��zt���T}W;a9Mk�~XG�Hlm����ϫ�$W�g�D���U�+gp}��1T��\�y�~�s>��C�z�F�y��M�N���y����n��U��1�q���-��*�ѭ��;��A	P�׏�`�}�P4R�ɇQ����S.i�H슌[2�p���f���1�/=����b�L?E��|!�u�;q<��$����.ϽE^ʿWS$����yJ�,���s�g�+���p3�{�45�]X��9�=76NY_�ys �����*�_�PU���E��Ek�5>�v�qcY]z�����'��(�����A��B��wgT@~UYM�1^5�O�	Y��ٰ0԰\�k�R�31-=�|�8=�#�w�wjF�SY���U7{�����P�J��E�_�A���д�Y�"u��*\+ J[�YB���Kd&ۥ�X^o;L�a�A�����i㛦0��¯�3[R\��ç���"C����B}s����/�OɈ-�:<���W�BG���˖��X%��猃�$>�	"�a�4h�K8�^2}��9:�nA}#N�/���*��� &9���w�) pI>��� ���:\̞���ĺ��&W4��3��+�˭�a��"
�M��<��%�����-�iW���%n�q��W��WƲΈ��'[ľ�V��SCI�qqgn�J�z�p�JL	��Cz���P��j\%0�ݢ��%wz���5i���w8Jr�g��Բ.�S4����aE�u A�F�{��J*�]���T���}���i�'���t2�j�+�1��ah �brYp���)�����r2�SI���im��7�Q�8���NoYRRn'�'�r}B�Y����Oe����Rj�M�o� ��x��@A��4Z�籐����1��f�-�ZF-�i&�x�C=�W�n���4�N��٥%�y�p��`��|(����`}o�0���D�k���V �g6��%�.p �i��}{L�x�n|�\A`a1h��8q힣����#��6u�9<:d���$A��j����O$/U�H駬�%�����1V5M��V�?߯4����;lDwkGn������aH�H-ڧ9���ߏ�@�+��A#'h���d.�I@mń#h%o���H��C4�܃��(rQ�i��(,mFߋ)��sf�N��[x� o�����]B����o�vSǑ_�����>�&���\,�d[�ђ��A���s=�U���z�5K�a�'7d
m�}@|l\���@����}��� kʋ�L�	��^����49�뒿�L��T�����`�LZ]bs��{�^��#�6(;�a�,$eW|�tB�2[��먉�1yؼ�gHwmH�ld2Aڏ�>��8��ٞ��'�$��b#�<zo����a���>o��܁2�����Ɛ0R�&�
]s�|���jt��9��c�R��k-c�܋�%�D�3�#a�<$e3��!�R�Ï2�Z��tlc���F�-��/�&?�lʇP���{���^�'Je�zqidxH-h)�r ֟��-�D^mW�Y�p���G�Tm#R#�_7(DOPt��>�{t[����ف���ՌK�n=y�2�$�K
%	r�������&!`�WH>�d��%�ű�E.�����bsM5Nd:i!��D2��;ŗ�N� 7x����hߊ��0�0��U�}�z9��܉ļ�ZX�eܯ�c,�H*T��J�C��K~����ag��j0�Sbey�`W( v�d�U(�&��V���Y[�)�䯔M�P�cW0���9|U>� ��#~/��d]��o}�x���y�l��dd��Y��o7�_%����c��Ѓ���V�baEVa+H�gKa!GA/_������o��TU"|���UԴ�J[PK#�(c�u_r� p�ݢ�ˉ�:%��;gT��U�d?��h��f�}=�ֲ� ڸ���X�i˭� sﭱKO�b�͆�W��g�;����`k���;�e����a]Y�jU�FU��p\�03��[����9}���>�ڪ��ႎk�2G�]:�pux�'��W�WU�G�3h�6���rv�&1؃UxM;s"E�`�5�eu*\K���cv���!��(��[��A�$�Z����T���v�Ǟ�x�pʻ9�.�g
���h�,�=&P�|�Yx�E=g���� ��	�L�� o/��!�#��rr΄1�N)�QO1�*CPJ��7:��:0�w��T���C����쯡����Ɵ.�A��je���@&ӕ�������s�>���!��9 x
�/�S�;
������R�4���ݼf������D���j�Q��{��=��������ʬs��1K9;:�q-���z�M���d����ީw�P�⡊ŵGd��f��e`'�P�s��3�#�TQ��6=��֬��JB���grh�WJJ�@q�gbA�Q�8)������z*`^�RG�R���iLd�+ʙ�?uQ�#׹�c�?{��CrcI�� ^��OO�ТP �B�,!�ʙ���w�ߌ/e$��7Y^O�6��_�׽ml��	F��Q����͛��F�����f	�-���MG+��tCx���Č�����xdu,w{�x�:I.f�h��Ԡ�^S|R��y�w�H��B[���f	zU��s���7	��t��V�UA4P*�����	,�_��3�(Q�!���.�w����N�Ǎ{���@�W6!�3ԇu�y(�;�;���\�����}��E;y��0��/[J��׸D��9�]��Q����Ϊ�:��S���lg��F�#�)#q/����-�d<�n;�n�M@�j��z:!峃뉔�f]�N�U1T��ԙ{�?�H?[��|��n��*�����l�����b" ~Y�VV��F��H�=J�˟�|h���k��Y�� 4MZ�p-tJr�#�mp--���6�n�K�)K�_r-�[� aS��ee$U�h��pBJ�R�a�xE�B��uk�1hᓆ6v�.�G$˓x���y���`�X�Ǭ���Y#W�?}f���a%P��xw6�-���	�gK=]��빊��D�Å��I[r�[�>�����Ƨ�ܷ��`�ti�s/�l��b��n�瞆�:����F3�������D���JD3�^�/�֡�hN|{��v{��`�tj�%�\�|�g��r�_�F��>#�k�h�3�wT'~�9���P�C�9:��Z%k����n%����������Z����vBB��s�`�T�3pW���Wy��_4a�߆�0b��ɍ������P��fD��d%9��P
A�S��)B�-l3(ڝ0���IĤm�qi�ݟ��ܼ1�lzSS#�<F�6����++���$�Ք��ا���_�[�$�A��]i�=~��~�H�������Ŕl�^��e�C��3C����q���A6P���A�Ё�
hkM��(�G�)��_�e��)w*E\ģɟ4|����\�=�1�I��"�:�h&�ʪ�{DI2�Ce��-��G�6
@�ێ�oE�;���`y9[;;��s1S��S����	ډý��k��p
r؍�8UA%����T�/�FU5]�jN٤�f�Sb���x�~0Lʮ�1��Q��޳�a�3E3�$M�J`��x�|^�u'#�J��:*�$��^ZX�&��&��z��k�8O� ��5��p {���IC*c�)Ⱦ�zv�9��<i�\��>_ai������c>i�)[xpʹ���8�w��',g��D�F�C��¾�R" &��K~ku:��E��=�@���	e��蓍�W��hrE�2�:31�8t�p��v(O��J�3�4��+��j(��W�?9r!��M۶w+,GG$1j�Qq N!�<�nr=R�H:�l�dwim>8��Mۅ"�v�dA���Ժ��@�7[� K�D��^���P�3��h�/Q�_6���xIA9���m�F��݄\��
Y��!&+ө�W��2�lA����U-�a��;><T�����A�/�ˎ�f)�<K�s��hM�{��/H��x����#���ܑ_Uݝ�N9��qA �Fn���ܫ�����ݐ2H0�����v�z���%�pj]���Z�^l���F��ܡ[Ю��Z��8X����~|F̎a</t��'k�:ɝ4&DKN�S`-z$��eWڥ�~���v��BJ���O�H���9��h�}�*Nd�P�a,����,�K�Ds�	�a"����a��a¤5��-���'"�H�<13���
�qH����z�B{����ZO\����:�^J��m4���z72>�q�lx�B����;L0��Ԛ^�(t���T�#�y�?ݳU���EB�C^Q@'���頻�È&�m�}�0mYS/� �����XA�M�s�l
_��� (/�]�N~�v8���ŀ��\�<�C:�V"h&��C3�N\�צc���VB���B��^����x�3Ѣh��k
>	i�gJE�JP��=1(�y�A�uB��x>��W�Q���f��ޙ�
��QaLԼI}o�ql$K<dkm���A�i"�iN�_/$�=��{�i_:��UE_vvHn��vA�ɿd���z�2@�r����fpG>4������Gmݟ��#�꺙?u8�-��g�0��'�&�=�i���%�_U}���I��u!t<X�(�	�k�� �_t"��G �w|��"f�?
��ԋz��A�?���!vl�y�"�z��u4n����^	�C�ˀA�{����}!����Bi��B:[Ϝ��p�9�5���^�Xvfp)o��y��Z~��л�C'-�Dr08��T��%�����8M�s�a� �K�����tL������n=Zn#�cJns)[0�Ga���| q��@�J �k�^m9�+���Qu^�sh���
��tׂ[):�����$lͪOB*z��CjJ��a���v4@]ކ�[EVc3�M8�G�39)~؈ǈ�/�#$�A�<Z�]�n4�� q��3��������&����zS�n5M��Ԕ0Y�6��˺���
��2&�&da���ݻ7�u�>��L,#{�1 ���\����4��I{Ib�y�N\��z�Xڧ$9}���(��a��XJ�Ft-yrBV������m)M���U���I���+��<�{�T�lp��>��ƺ��xmz0��4�}�������8�$Z������[]F����r�*�&s/���V��l�E�L�W�h;�o|���C�u����lħ�1�4�mX'�A�?6+	ع�
\/!�}�F/Ԉ��E���}��0�����T�DI�y
F?�4��ȴlڤy��!I4�R)dNҶǶ��>��{*�^8��k��@ǖY͖T5=>PN�,�r�|�$c�-����e�y�R9�	�N���5�
~���F�F�`Dysc���WJ4
�R"�%^b��Dʱ��/��8�	Ld��1�`��Gq�L*auY�Ix��B�	�i�坍��i����f:��b�k�J�0<R�F�Y�SO����IsNj�/��n�`��MWӚW� ����V���\���	��&�5��	�|�relq��dvq��5@;̫(�B��@�E�>��Nۢ~�_Jy��v�"�e��H���}��o):mQ �;2�_�HT,��!���]		`�t�t�sE�Y�x�DGv6:�^���v�{�{X*�SO�w:�3�JHxy�J]����P���>�W͗G5�H�<#9�m|�
BL��x������*m)�t�H���$�P���#�]Y����ܯ"�|y���f.��[&�C<%7��B�a�g�'UC)���'s�$�t�8�����y�V{
���C&[9V��������]r*��V<�1����AjV��(r���+��I���� ��*��L��P�a��\��yp?��ʯn��`���_3��?����"H� ��ɭ5w����Պ&BbZ��'�xٍ�3�S_E�������l,"��SXPxM����R���1Y�Q�)pkf�\�U-�C�7�+����C$��<��tX�z����H�Ǒ��򂳿��uUC�Go\�}��i�pl�.�z��y�Yek[\#�rqx��T~�ӽ��4a�m�C�����'��k!_03�%�۸��}A�Ub �]�9���I8j�%^�4�L��c�̊�7���R�a�H�@�-�i���U��l�Rs�W��=E��>�l4�"L�S�V�Q��op���Xpn��ф��J�qB�d���A�\�P����:�:�5�7�0}��R�C��q�}O�����v%Ȅ5^�f�,�~�=ɧ��&|����	�mȣ:�$��X�j�2ͩfb�����G�<�،���d��$�G�~����$����Pǎ7��A����Y�#_��������M���Xv�v���kVj�T�U��s��.�	6��U@&���q��;� �4A������>^*�Ҽ��b��aW���0�1݂�,;�g�H�5y@U�g-d`���;��{�ʡ#N�|*'�-n��<����ׄINB��Fhi�0�;�ڡ�5<��]O���/:�2j�y�ɥ��~��W?m�o^�n�j�����$k�'�g����v<�ݮ�?Dɵ�o8��t�M��mz�}lbą�ڪ�1��k�ы ww:\���p�7Ad��y̘l��C@0y��hS��K�ʴ-ş���h*#t�ޓs&>OU�:���5�����Rߧ�;�>�v,ԖWƤ���<�Z[��M�?"��=8Ɣ�Ew2�uʦx��D�s�7�G0�Rh��J���r!]0.�'�iQ��t�%@3�,�3ucc�y�z�P`#��`Cd�А���h]�KNy�b)
�.��� 0i��PnT��-^�A�V#N�7|�����#_�<���;�ޓ0�lQ�%��w1�)`��sɃ��3P�cY,{L4�@>�J�� �� �/���-ԅ9�w����Y�Wqnڤ�v������ߴ�i�b%Xs�L*X�`�؃޴���l��IŤ�wVKm�N7�7;�8���aB�V,	Sc�G����l��1�>8��t�_�D$�ĭ��\��(!٣�����_�~�G<�e�e����Q�/-g3r���}��)�~�״-xG>�4T>T4�S(�BeZ�������yN6QK�1�&6�;��@��HkJ�l��׬*R�\Si%Q�ż���Q`��u���A���eO?&����?�����9��b((��f�#)�D9B��V�9%�����P�:�z�_���k�Ҧ*��"���Ly��ܬ|$�J �;m�畁M��eˤ7�K8��.-&�� L$ɋ7������5R>^�o4���@5�C�jx����F-t\v��d�,�����h���}��05ѼĿ��O;��ߣd�
��ѯ�+P�&�4H��'Z.4�ͱ=?p�-\���TqFHؐc9�V�-	�� [���d�����bw)f���� ]f�K$���̃2�[��^�S�D��۲���6��t3�BA����	}K	�|}L.%/�Ҥǣ�y� ��I1M�J��Tc[�S/�$���2�Տe�ө���]i>�L׹&v2Z���I�/3/N�	�V��"�g+vSʽm~� M-��t�Ni�/��;�[]��ǚ[�͝'�A�p����e�jl�?�	����M<�7������ma(��s (h�7ךq 4��P%�?��L[~�E��5���1�A,��dSW��[���7�=�@ s����|T�|�i�M��b�H����Je_e/X{�[�>?�I ���)կ���*iU�Q�Gߘ�?g7,-��K�;�Kv�c59�;���{h�2􂺠���V+CL�N�g�R𐊼66�����#���i(Qu�"��C�;4v�	8�Vf��@�����D�Vqq�1g򊓓��\�Ƒ/S�E��2S�i���v�qޜw��P��p�w#����˓�f�����ZT���8S�ot�(�d��U�6�_��F������K�=�Z��Z��x*��6=Ў	�.�:f�v�7i��vGVP���~�\�@�&�2��U3a_��{��V�L��vCq� 
�} ���5�P!���D��237��hD�
�X���2! &'��[�J�ﴙ���S2�$��pnhaD�&'X-_�������Q�^R�0Ex��@�zݩf=o/3����,5��&�5�CBB
pr�	@dʰ�&ä�cU��$�S��f���d{_���8(d�ۄ�݈�\r`x�U�����!0`�$��@ �~]rQi�Yy]�lԿ�O�8�Tӹ�BAS	x�ڍ�Pdg�r�,�
n�ڶ��ò�[�y%�ZYհ�����QiE[<�0\G%%�Fl7v I5!e��1���m�r
ɮJ�9�0��vF�u���sX�����{vN��Z{pɈ���x�}���ب,���,q�~;�-殰�����͎�d~!�f�q ��:���I�ͨE�c�����j��u�!N�3�v���L�?E�p|*a"Y]�8rvz����
S#� �aƻ�Qڂ�3��ۣi��.���z�n*��\��d���"��D�/q�%����Or��)c�<���7�g']�oH��v%ev8�J2
��L�Fb?kf��揙���U�Mo��{�|�nй(|�!ڭ�Q�]�6��~#�/��|��P�6
��Ô�Sx��h�D�QT��#�@	�~�!�z�/�b��rx;���d����e�RŠ�)�V2��2���d�c}-!Pl"oUZ|	c��5�AKK��*��P�KY�.�e0���]��D5���	�;�kc�6dڸ�]	�PyJPvl)M)�j�ǕR=����#qx����;/�Oc~5]��$�\�� i�n���1i�6\T����IY8�Z�g6��a������uG�p��g�{����判���+�Am#���ue��A]�yw.�ȅ��5߹����RV�H^�YS��3q��Kt$I�0 ٟЗL�
E��M��g(�t�vS�𸣒���
i��"�����44.�'��fB2���i</�m�",�FEY.���kY$�����j[��0�~C��Jg�#:��7��Q�����O&��5.�L�×C�~ɟq-E8�{<`ѝ�/�{D]��Fv�ݯ������(��'��<��K���Y���x#Dsʍ�5���3"�:��|�� oJ�s	~D�NA����뻎19�yN
aQ�
��4XrC�ǋ=���!� ����*�v��h�Ɵ� �}>�\L���a�ݾ��(Lۉ��iz�)�n�Nr�0���N/�h�G����g�~%��� �!<�%Y6��z3��6"q�$� �Q#��߳���Z3�d���i& ɐ��-֎��s�Hxe�ŉRQ�O)�c�K+�/�S�P\�SP�5 �ǅ�e:p����� m]&�]�8��s����yp,@�k���k�C��V:Ũ(B#E���t��[!�L�8�uF���
��	��*���,p�}>��qr`}�{h�ֿ0�=uάL�����I&�I�E�� ��U%�f�������B�#��a�~aoIm�?�c�a��^G2C@A�<D�_���ql��*�n��������\����`��L���7�_��^�����6���m������R���C�U�ȡ�� >�4���ꍠ7��.<�2�5�,����6;�>�*��;���L`�0�d��<�[82���F�����c�θ�H��.	��8Ϧv+��6M ��Zm�_?�#����2�C�NƓsN��$_rdh�͛]%���e;�ѐ
����]��SY-	�"R�. ?�w��L�is[n�E�Z� ������rF�ɟu�"����ɦ�D�y�V�$�\���s�����c��2���{y;���|Ԡ;Wd�?���tJa�m��]�Z�
p�x�߇�B3H���+�`�~LM��,��?���R�):bEu4�|N.�ů�[���,�EV�����;j�7��e����;u�����P����C���4�?� ��f�$�'��_$����&W�t<�F��|l�H��l}Gh�_؇%�b�h�;(m�� �H��n���\���$Y������3(u���E�Yr���ͳ'&�)h6�Q7-�7���p������1d�.��f�L�����:�0��g�`4�3y�Խ����p��q��^|�5q��9ih��jcɡxv���]����^"%y�)�|�L�X{�|�4�G���l�{���b����K��J��H��e�p5@^>����گ�w��k�������Tw�̫�Z.�	�aLjf_��)�*[��O�-��,ݼ�JɅ���Z��}��`��a�
�s��#�4m�>Q��:��B�,�e_�XK��Q'�&�ŧ��2ىs�݅���9�{0���)��.��i�bk$�u��`�����͛�610r����!h2A�~z���
XuB �x:��	C��Ш�%�i<>c��Q�{� ���x���WL���iH<�e��X��CK1�\�!#la���u�NBeV�R�,N�R��\��柁l,�W�r�6�����ׂ��^���]�p��H|���H"d�/��R�NQ��ṽvڧ=�"��F�Îl���l9ұ��s�Zӧ�:+�D�\e��fE��w@�����Y�I�H���
mۏ���\��Y*]@:�{���B:]IBV��-}@���-A#�5����5M?u�_a�H�tF<#����$��������ӯ/ƴ擥�jW}�	f}�#�͸�������C1��V1.�-�t�<ٓ(�3�4@π���l�E{�j�}w��M�o������Ҏ%�RT��MκL�� �%\�N��7+Yb�K}z�^��^f�Ĩ�"����g���� Z��Y�B�k�E5g�T��\ �ǬM.8TU����s�o���F�®����^H�ԅ�%�<����r �ș�`�A-\V�ED<�G���0ުO�;	���rD
�o�Vty�����������h�/���r�7n�#ԞF=��eU��=������\7�W��H�hg��`��Χ��x�U����{�8��1?L����d�<t�{j�h��~g����P��)l}K-�i�m(�B��vb�
޸	�=4�� ���N��طF�����S}_PV�S�%��E�9v<�����{n�����Q����L�������m�w��|��(N>���	=��W?��F��Q¶1��٧�b���o��⏈)�rݾ*n1����JJ%���?v5x�A���ٓ�f�������-�����x��gI+�3���jN�ud/��Y�ʝ�GK������V`1M+��?�:��$�Տ�n˼Qh^~��7��h8�K��'q�x�_�u�U�$� QS��V�yV�y���o'���Ξ��DW/Э���nkǩײpLL�"ES���'FH���u�u�I�M_��ϛҭU���j�8�UU�.�렷�)~�b	C%�>d
V��*A�s~��|!vt��K���H�:�[��w�y{�����ksL��=ǤwQ����ѧ���ޛ�헥��đ�� ��/�r�t��܃\�?�����fP�ϰI/1��@	 �MtMy���d�Kt��gS�"H�Rqf"ɃP&�� �p�M���O�W��Qq�j�sԝ��[@3䟠������nX_�+�.�*�PRp:�^��������>B%0�J��er��E� �̐FG�kIe����fQ9y�T���|h[
*e�:��4D7h�W�!n!�P����O��A��p��5��yI��:���c ]�\@���O��]p�C��T�]m)����ҧ�D>�4:|)u����ˈ�tΰ\C���>����$�C�H���׾7g-�G�_O�y}಩����1h N�lDPi��?��'$;7�xD�lpM�b~:6X$R!��p��"C�In�P����{��d�dwUs���f~��{
�K7�̀��̺m��jqc��͔wcEj����l����n��d� �GyX'����_SFOWƕ������������'5�w�@iZ,���`���vь@j���Z#�R<|7�=���c�{�2��%R�d=-B֤�M/w�%��i3�h���g�0P�zEuV$�Hb���}��q�"P�&-@�o�M��%_u�M�"����/��{����MX����u��;�3N�i�w-lrVq���vn��eG�^ؼ`Y����}/�y9��ޛ���켷&�B�#;n�z@���b���z���|~����}-L��Knc�|���PR��Tl�`��T����d"C^�&4�$5�:�`�SJ��~&���E�s֙�'�k:~��Qm?T���`Qi����];�V.��̪uc����Bmͧľ&KSD����8�W�^(��"���lc�N�x)sϨ{1�����p̟r�[�ޮ+��5-����e��]_�F�E�.*���1K\g�`Ȝ�k�����(3$L�gCq}A���]
=	z��L�KS�DP��Lb�NJ0�����(����Q$��+ �A{���&[�DV�(t�T:1"�m�5�Z���}�{��\ �Uf��T�ZJ1�"�Kz]j�ХYn���Sڃ�Z::;��g[����x \���s�;Z6P���bL2�v�/��������KY�cX8��yyoK�3��
0��|ZU�?1f��� t�	V��@� �qAq\�7�,���M]�	��
������#�S��P�6t�"٘���� 6�鈯���ʀ$v�3��1
_}b�����	;J�\nү�6'�A�����a+�V��[���حiB�=��@�9���RdCee����n��6�hz��x���jC-��*��C�L�>D��S�Gh�0N?���j�!�ˏ�����`���Ԣ�:���:�X s�)�y��X���es"���ʸ�����h�Ͼ��8_f��'��9(���Q���춝�tե�yW����ЋI�/�jH���$�J� ���^z���Z|��y|K~ɝ�e����\�|�-�M��9gǌ`O���|��pxxCdؿ�μ&L�,vc�X�J$A� ��]�v1}�[�������Cj$�LB4�Z��t{L��^�"`���[�;�㒖�N�)�͕��bJfE��|��io��cJ�Q��-K�����6v�� �n$�|X�?C\�TF�~�kb2n�ph�La���(��t��2�6x�Jɸ��V���]S�X_]�t9�3���S(�:�M8�Өi������Y�Dۉ��U����E�u��f��ǀ��[CMŁ=-��u�ha�'xw]+,Z��q/��Z*���u�[�e�ŷ�0��K�я�W3TN����ã�	��R]5�+�6�N6a:X��=�m ~��?� �n�Gk��P^^ht��IaBr�%^͖G�]�������������⌟�N���:i�#"���?�D���E#�2���y��ЌO!�Z_t���?���8*6�Xe�KM�6G��(A����O����p7���j�c�e(�@��C�Auk�@`�4Fפ#=��Y۹�/����:}I=w�\Zz�"�+&��z_g��R��5H��^O	�7U mR��$6t2��/7%����~MhV���S��^�����[He)ҧ�;ڟ}'��YMq?sa��Hf]�us��q�/�����m�\j�`D�`���q/� ��6�-U��/(��T�.��+���s���
�a���I�`�g�и�I�!�>��r�h`�I�>�<���|�E�{p�� ��h�pF��o��)7�>�1��6�G<��f6�%<�G�O�ޓf���2\�/W}5�z�j��=i�Xnsj�9��M,�aŭ]C{!�C�r�H�T֐̈
܀wE��"N�*�Cu4���[t������W����&�b����F~��y�G"�{��oOm����?�lc4�vc�z��~���p�W���r;!I)&�O��6pN�p�M7�x/�,p_P/��kY7D��l[�W�Xڅ�r���S]&�CΫ v����(�
�G��s*a� �p+o�y$X�Ex�@���0kYޯ2Ս~z�.G�}�r*��̢����!K�sU�-v��J[��&�*N!{5��k$�t�i4Z�6'������^uFW�J��q^�b�>���U���Gp�Yw��34}���kF�ɦ	$H����C�P*��|�y2�`�i7�-�e���'t4�m11;�YK����ID���m���3�[>G?�K��3Di�8�`���L�mU�r�[�kUQ�(��^�>7����ݔ��'�+��SJKh�]-H�Y�ZҔ�n��;@����\�ӭ�ڑ�X.of��W+;A���yr����uyUWcًу�Գ�a��V�nC*��c����J����e�	�*����63��$VNo�N�(��=��~�o*ޜ�$$��߰g�ڠ��OYG�k�Ж#��b�e�읙�	�Q-��s-ų��@)�Z�2��GjI�̌�$�P:�y�>��ѯ�G\�Ţ�VH�[1S���*7�����L��cğ+0eL����98�Y}���2��۾����LYsRLL1��h@"�5��Yh�v�YFo��ԞoB���Й�K��ǜ�e^-#��?�lK��Jo$�g!��F�ӑ�L��n�h�2����_�+�s4����	'��`|��7�����
��	y<}U[�w��⮾"����Ŵ�^�{(��5�q�bߥ����w���d�J�̊j���]�Ӏ�m~��X�ݤE� �GI�f�A-��I}_������ރ(⭹�e��?�O�$�c����d�TW<�S�z|�"�E�y��\�0zJ3�W	�����[{���1S �W�5��*z��q��Z��H0��N��в(
'`E�������¾�q��K3���*�!E��Y4�7�ݢZ���,g���P?.�	/�7K�[kSq���]��-���4�����W,a�z��j�/aU3����Դ���ܗ���WB��ҝbM�R7��fSH��o�>v?�R�D�xo����0����7��LYgXB6h�N�RL!�`ǆ�&� ������� f�7���]�����/���؀�~�P ������������d��6Y%�!�����L��ao B=F`w`�\W�Bd������^Z:������F��2�V՜z/m]x�FOއ�u�ÊXS;�Ro�E�z,�w�������Ý����R�N��kiz!����n�"Q�rDR�zs���!	�(�����_=M>���X�YŠ��h���ȶ����Uz���ac��9_���_Bѧ��.»��^E�ٷa/�׭��[?�n?�m���	��fL%��E���ޕ�έX�Iל	Y���j����w��(�v�M�b�}6EaҘ�u����̲��!��S�]e�0�\v��b_{�� ����^�M�-����	���b��J��Х��~8�P����E��o�a���r�>1s�^�_��*�T�ˢK"iR�
�e'���@�����֔ �Q�=�_���2bЊ��J[B� ��Օ�p���������a�e
Pny`z��
�j�n�5e��]	��6��^pM��ѷ��'o�{H��y�|��XS��'<�%���n����}�gt�k[�����s|#��s$�UN��k��31�KBb����|�w���g�ߟkET��ћ��M-'@Z�:�jr̹V-��b+G�(�~���Z�s2А�S~���/w���`����QI��j���"TS5�g�w�)�i��	�nƴ� :�a趪���k���g�؞Z���e;�:�&#��Γ_�RޢJ1VueE����}���$��J�A��C�o+>Ɣ����uЕ4!� vV��W�~�f�o�Ѷ4���"rt��2~�=����]�S3%�5��re6P�����Y鹞B79�j|A~xW��UA�V�4��?cm;8�����`K4%�7v��U.є��sj�|�닩ab,o	��,��d�,���`'�S�m�/q��깆��,����@7���{�v��P�Ι�L�e��>�����lj9���f͕K�}x���;\]_�&��3/_��oK�'W���Swu*7�Ǩpw"�:T�e!E����~rϔ���Ȇ�v�~'�/l�Щ�Â��,�o~���In�i?�(��b R�:��q���6j��	-B�@b�-{������;����;�8;�N��S�iV�LFc韴�� �2�SBς�zC;���h�����ՓEu�)����}p�ƨ���J�	��om�@�>lX�U��'@c=�C��Zp�z�G��Y,���)Q9#Ӆ�Z�km	S�!7�Wnߌx+���1�S��$���m����%f�5Z�Xȣ�D|
c��]�M���M�b70�
2�rp��//[��#�Eq�r��t-��7m��F��zc�a�p
�⢟m���%ɀ����X������$�K��=A-�N�7�����8 7d���!�Kv&1)}��F�-�%7��B���ZՇ@�m �_w..�H�K��dF�B��Dp��3.��9���+�R��" ��3���Ɩ�6�$'	�3e--{�� �N���o�����yf^����a�9����|[���4Ds���t
�S�I��o�z z��VWc`����}�E,�Z�#��6h�������,K�V�E�Uu<��n?_�Y%�{�.'�|jw�w]<V3�wo^��0�>5�X{�#T��&a��xݝ��'蒯,��͂��$�*��`�����م��Cd�{�G5l���~�ۅ`m�v?N/V�v[�%7N̅L�j���ý�QvYR�|���re�9jV���'�K���I&Y�_���c4 ��+�Ӡ�G����f��9pF�ܱ�"pv���W2#�� kϟ���*߷0�Y�x���C܏ĵy���z0��� ���k'�n��������������Y�s�D��V�ƙ��S�g���$�m�?2�?��D��T�.ć�S}��$*�0��
���C��4��r����G9˭�^����B:�����^d�}�O&��/�q7@��'(T���o�46+�l���\���gZ�$d&}���bud�����u�o��x<j��@{����Ud��+`���\5����m~��f"��`fv5��6�f�:�R����Nv��!7��~�F^�:}ے1;(G_à�9���$k������Φ��̓�p� Z�ac�^���8�y����^��GN�n��S0�C�$뺯-�U�g����N{��ۚ���	
b�\�B�~kO�(��~�o{X�L��ps�z`N"kۆ��T��"�^�t~�k�f�
���(���k��C�����=*��x*��LKr�[�q�?����p�����f�4e��X !u#������=ԭ+6|�`�/�[=��Q�;���$��H��L�I?�'�$�RknJ���J�}�׶X���� &ˢ���Y�l���T\�E�w�?�W��Mu8bj�a���i����0d�8��r��e!�<��q��t���?^�����jN���xht�-��9�Y�"[����zB�=�2�w*Ai�F74����A���2g�_@h��݌�,�^=&���R�R�q��|�&��"�+���4uI�߽�v1����bm��R���H�1?>��g�?��$°.h���\���m7����=���: h�<<:k��	�`���Y��o���#^g2�1��/`��2��W��(s�15��p.Ƥb��Ur�v���m~�pX���g(���=�`���!�9�2�Z��z��}؁X�Gb�x�K�"_�U�b�\�94JN�Ojd���r���@ xJ'��}�� @(
GZ�*p��ug��=�W%�/�#�y��C����$�2c�������C��t,�r��ů�>�[7B�k����B�ࢡ �`Ck��/�r��2<�V�oZd�+.'�a�2qg�F��fМ�� �)�2�Y	}���w����4K���\ϭ3��sHU�b:��������Hj��pťc��|5���	���)0�|�o�[�,�e�p�onj���2y���یC M�(h[F'�+������-� � �p�2;�{�����`���)��g����mZ����2�,��<�Q��p�X�1��юL�z8�k�����"1f�-��A�,R[���d�n]F&\�U���r�b�	���L�P��8�֓�,%��x�س�G`�(� Ru����{4�оgÝ�|?N`���a��ɜ��L�ͱZ|w�� �Y��»��NE��y$A�iދ�to�P=P>�y��W��1�����V��ױ�g���Ts��D�e�`����D��v���V�����&K�cJ/;v	���E31����3�*���c�˹��V�X}�8[ ���05�c���� ��1����E�e��P��&��=C9=/�ǯAz���=�X5��_�C
����v���2��N1�h��6c�Z��-f�Xr�����/��l@vÑ]��d'�0�Iכ�p|��Yhm��v?-=圫�sh��^$xES��E������gjn���XP��p#�^3v��Y�sk�V���e{(�+>',��"�רP�VX���;�^��8¦����� ׳qVQۜ��U�XUZ���x�������k�9�4��W	��=��w�r�U��I��-`�*��Јǅ���1�v�7����z9$�H1fFZO@KcQ
����9�"ɘH[^�Bb�~�A�DЅsຖ�Ξ@�|�	�|�mq����]f#;AZ�ot-�(�u+���Ǡ�3�Io�Y`#�>t�&p\ނڳ�+�'�On~'`�����Z������h�O�Ԭ�����?ԍ����:�bN���T�*�(Y�,�׆E=���>�7 q�f�-G��4��~�T��)� �q���B(�j��].�TW l��2��h��th�v����0�>��1�\ڃY�b4H2<�ZZ���y==���WA��8L�-u�Z�k"������{r�>zX�Q��og=�^-��ؑ���/ۼ�C�r��r��:[��`u���8�~��i$���~	���mzOKCd�Y"���V`�VV�c�A��-6�x������B����F�n=���	���H��
�>���� ����D]%�=9#U{����R���&K#T��w!��.z ��N�H�{&ˆ��3�t�m�';����]��)#���m�
]�����zJ�NfQ�xC7��o��%քƲm�2
��Nb A�?o�3��^ma�n��є�G+hsOU�E�d�4M���6r����A�DSw�NQ�{P|<���
m�ʵ�������+�-k-�
�����S�:�1��s���o�O��yO)���-�z��� ��o�g�-����l`��V�3Ո�N�P��L��ѩ`� �*�p��בn�������L������\�ӱ�^����H�p_q��ƷC�8,~��E-ӵ&9�fn�k�N'������w��4$���cU@��6,��w���/�hݱ`��q&��1�_�Ҧ�a�\L:�D�f��\����A��:��ֺ� h^ר:`_�B��B�X��}������p�]�X�U�{T��^�w6*�e��q�]%��h�]�����/v��Z���W2^w"mn�P��^ez`W�5�&7G�W�۞�-"�(nw��$�!����ʟN��:��$��bS'LS(
	��#��8R)棥�H�����LةMe�Q{���l��c�	�"y!��J��	�M��.�$��{�!)�����I\�<���3��:f{B>��1=3N�V&L��#Q��Ѭ�P޲w���{ܡY{	g#�y|4�������d��2�08Z�b�#/n����gH/��"���K�E�OM�k�Z����pߦ�X9�SF�E�#�d^�M
��D��b�bh������kd!o�Z��?��X�Jl����U����뮰�A4%�؄�lƪ4Dp@�Z��q�ӎ���bu�PVzI0��2nC�oʨ~p�q����0?�{9�_�)��&��&F�<m�����m^*,���Zk��6��DV��n�K���Ll=�Avp�悈}Ob�k�)��wf}9x6&��vt�w��9�pd�e��.�Z�f[�t�V�7v�V������Ы.�Z'�gf�&��L�']��!���e��4����f>�<.-?�-Ծҧn�fdF�%K�C>��O��!�v%?�DKlؙ��{�����l�i�q��?�����W�
�^"c����R}Y�S���@=>ֽ��)��qΩ�6]?����c�4��c��)q����e�ѿy����];3Sp�ߥ��F��Ք����&���?�	��u�.Y,����d(�ۮ�_3�4sI�䅅�U�ͯ��J�kG���vy+sh+B�M��Y���2�do.B��뽐�T+f�o���嫍�tL�	�x2�<"_���ku������1�*�2��k�����b�
�D��0�[�O�e�5QS����G�_W�������[)l�}� `1��v��vr|����riX-����?�F̋�|��v`46�u�Ӏ�)g�_�ҳ��B2<�G�H�0�����\8u7�"7E������CW���j��������0�B���X������p����� ��
�|nD���d�Gۅ
�w�?��P��у���&eS�J�����d�j�BV"i
S魁�Y,��e��Mb���\�sԖ+�2{y`��iz��XN�`��e��+��M���(p.��A�BE�HQZ� �"zВhJk�!�,���M�Y���m�>U��*�4z��������J�/�q췒��W�l�h}�7����K��q��>��-�Rf7�Ž��,s{�&�1����,���E>� �J���R>�em��g��[��鱺��ߦ��9@St�$�؟Ӄ�lƀS�E�i��K�t��L�_�{5�J�HC�����Tr���ڧ��4wFoM[�}V}���	�N��6Lm�AbO��x�X�.ǮyT� ��L�=����ϪD��kp��[����u��������L#��q������ץ������E��k_:WJJ�G��}U�����o�(� }S�%��*}�R�l�ZȉӼA.�ߑ#ʄ�E�K2���0�x���X�^˘X;mf�n{)�Q��*.�s��6�50����NG���Q��ڮ ��FH��{�P��z;�8��J��@{�鸆���U� �)>��7	��������>"a��X��0��&����qUㅋ���\֮�=�1ĘP)Y�d��<�b	F�b���&�+X?�nͨ+K�G� u�����/���-0�/3���ثξޟc�¹jh��S�7�B���@.����f�kU�������2f�'|�078)��1?�Rm��!�\���r���db`��vD��L�K��j�5`�Pe�N������$)����)"�ܭ"��i�Ș��Q�C�rfk`�d@gJ�pϠ ��1���$A�
kۜGc���`W��?g��F��+V�ߛ��G"��|��0�3�F,�"�:�~�C����'�C�+R�Ш9yc�?�[�M�s�#��ʳ�T!�����T�G����ji[c�_:�E#z`o���*R̊�6Z1��h�F5�ֆ� of`8��2�Z�ը��du��_/kј�6�mZp�%��"�E��44����uSǸ]����Yih��6ΆCܡ�5E��ե"_R౾6���"(�1���E�M��?���̦��]��S0��T~g '@�����"Ҧ�5��1
ٻ�J˗��l�޻�#3��.���f<�{쪖~���r��k7d�V��g�(e(�%&��R8�C7"��,IٶB�H��P��,:��p� M{{+ ���2��Y>ե��X�c��t�J����Y0rvS�]#k���Z>���񗺩��{�F�D�D$K#;� ��bM��̓��mhq������7��Y'�!���8kZ`�pF�Ĥ��ù�w�
Y�d��U��B��(��%�'�kˑuh�ma����@�i4�Pzt�>+qR9ӫ�t�x��c��!�<��c���#ڮ��V��o�Ԡ�Ի�0i������k�A�"�/����3@	Z�|5	^"х��b���9Y��9}�>({'��@��k�Yۦ�lh�Ԫ-���ح��3���4��^q�%3=���-Z"a�c��v퍾�8
df5�(q2)�(�	c]�$�(!�oKA�"���/d���|����
����Dy�SB�|��p���'#Z5��w�(�Ru3�B/���s}��.d>x���/wVn���[@`;qB[cƮ�qJ�������@ �Pm�Di�k�7�l�uyjaf���Z�}:8��$�0'�]��&[DrF�(ڔ��D\&G��ԃ�È��\n�X���lra {Wߦ�nE�s�^�G3_�%�
lB~%������9j�hۣ�w��٣��ϲVW���F3�\y�rF)���=CG�k�[��E���L@��Tg|��֛��;1��\�ǯ������Ys����鞀%a���i�o�~r|�S _@�y-�d��eyt����iO��ǉ�	n�m{.�Ș�_����A�e� �~F"�P2������A�Z6~�hL4oG(�4$3���Ӑ���|��4�1&��*�Y��I�"�HS�kLl�����7-�Z������ůkP��
����E��.�o_�At�W�&�������i�w����_9 6V�����)�/y���o�fk�{��c�}&D|͔�!�"����%�n����1��wJR�Vf�#�$4���_���M�`�,d�&��p0��s�B����t�Y)>(�	͙B��o+Լv彎��Y�ʊZ���Ü�]�%�_5sa�o�k���1���`p���QJ׏��+8����`d�K�r���,�K�� �xm�=Gf���������?ޖ,S�@�2l�����D#�lޓ�9�$+��1YS�"��`� =����Z��u[��@�0��2�����g�×2���NC��T �.S��D��|�j�[Oz@庈�'s��|p'�@W��+e�p	`��b�|�bLp�$�!]�1��|
���Q��w9ӪWZ��찂X�u������t>��X���� վ;�2�X�&mI!��s�Mg�N���W�;����/6�4�H+UE�d���������o6��w�����X$b��8|�~`X��h��X���'+w��,w�\���?|��
^��Kf0y��WI
���g�9�kX�������-7�-��(Z+���7�ȧx�|�~����tZ`��,�O�Ť��tK��l%�i�i�s(��By���-�f&IOW�[=��L�E	 �Uo�EZ^w����gʫ��Z
��3A.R,��W���:;>��.kxy�[*y��[�p����S��ӥ���@�5�ΆT�B��Z�}^S���w��2�����8]��f3ܑb�H*Q�j�Ɋ8�-�'`/��9��$p����(��ՑTi0���:|K�����d�X�M�����5X��'-c��Ԗy)p
�f|8'W�	�&][����XD��/���_����I �?=���m\�@����`ȩ�P	%�P<�^\�7l�丄�ʄ�,㏼���t2	/ͷ�q�P�I7�����B-��Ý=���G&�'M1�͜03���F�KΎ.A�u<�����O������s�}�N}{�l���3n[Gt�¡X-
�ˁ�r�kKQ�	���i�%�Rb�?�]�B�#���P�-=�������?�e@�5�SE��'��ǬW`��;�!ضt�b]��w�F�X'C/���u�g���v7�
���)ǆ�n�6��A��׃� ���I�T�'t�D���<�mùϯ0�¸��ui����8���q���0Ɛ���N����\���~I�xF��ps��+^�0}�	�z�8L��l5����TD��ʌ�#O�.��/+�a������LxF.30@Cn~���O���]��ɢ���!��ʿa�m�/�fM}�������?^���2=�g��t;�P�%���5��3�ؙ�M� ���|�m�z?0G��؉�'A�ҫSX�?gul����Sd�~��r��>���f����
z���i� ��5��}t�9okx�fO9��\d5'�eĈ+���.���o�����T��7y7�6t̝��lTu���"�G���L&_F$��oN��s�c�IU���K�{����Ȫ2��lS�3�I%c�W�֔��&�?v��S���|)�q����5X΅_�x>k�O4"�� ��_'��ߊ:{��K�m1������p�-|f��$���c�+��6��e���_�CC�'�^r�"��Mn���"�t#�����Xe��i�:�첀7C(a٘֌cW�I�_�a!��nm��$(�@��&��k�GSr^������Q�S�ߩ�W���b��Y�,�2�:�����T���c2N�)���
y`�(��*O�]+n9�6V	��x��er�(\�P^�)↛Y�|����>oҙ٧N���'	����q�������4�it5��[�*�ϑ����-��^g�i{ϓd��8�锫V@R�N�I�2*���h  uq��^��M�pRI�5�ZC�ob_��o���߉��&e�0�E����M�8<�(��x+�G�/9��7���i_ךu�$G�i�E�vȢ��[.��q����~�e�C�0�Ҷ��Q0pՅ}�<����n�v�k2T��s��pt.�`���X!�N�
��+�
u����m�P\��WIS���T����"hdj�	a��.����l��5�����7��Az�<坹�� z������c,�ҥ��\�Swr��^�-7#���H�$BZ*�?A�]�ئ��v��9�%���݋o��:����ЉZ�as�&M��W��o�&O�0rم��3�O)դ̠�؅%�(�D��5]A�r�%�!���:=��Z�3Z�����"/��
&�qm�L9
�g�' v$�`�0�6�9�<g��52��e_ے����P�D�v�񳶞�J��Lu4��v#�Z�Jf�S 6}�W���CNjSp�"�?A_��N�l&��p�.���P���Z�dZ�G��$�1t	1(|���I�v�t��fE�ܷ�]>�w�az�y�0%�V*9�	F�}��dർuY.�F��c�<$�h����z+�Y�ns����vv�A(u\�e&d�i
�KN�˚�ѯ��뜋�M�k,�0Z�{��hS�p�,1��k?�.�%i6�%w��A�ZA���ӲLy�TjlUIZ<Kd��wرb���izk�m+g��vL���^���<^�Iu�:����.q$�*�@����TϦ�dH�^�}��L�e5$����X�0��_��5�-J�J�Dz/% ���K���4��F!������i"�[|<�HY�U�Im�A4`��]46R�h��ɴ�ׅ��%�����OS;���S��"���}�YNش��{��"�^)j�O�~�����4/┪i��nD�[}��̦DO�/<6׉U@�@��_9W'�UP\فEB�#�Ld�<<�7�Q�QY���~R8�G�đ�O��SŔw*�M�7����%��#��G���Ua,�	N�����xtFgG-�Ar�?ݱ���p��LӚ�d��&��9;4��Bb�����!�@�8E��pr%+R讽Z��O\"g�l�soE�	o�H���h2�/��ٙ�n�۫�����L�ۘ����pv�2�'S��n^�Ԥۮ"��Wo�U��
5��Ba�$��0����k���s�&���(����������Mc�ϯ$[3oe�4Cԕ��G����z�s�z҄k��	%�
j.j���B1�1-��8F�	~�b1���l ZT*kb~��%`�f�r�G	&����4�RA��w�k��]�ς���ؑo��Iր�RIUw�(�i斸�$�ø[��u/U���(�!�Io�/&@�7���ސ��_�B>*ҊAm�~�q쫈����-���`G1���(ϱUi��͢��i����Y������6d7�l�ȩ�)��qU�z ��C..O�z�C�v�O:�üS����R}ӽ�츈��%uT�����lhw��6l(���M��c�M~������w���<bSGc���ez�͖�@{�Ǖ
<�h`xB6����������B"�ܝ��M8��n~o����g,���R���v@��ö_��I9u�%�'�,����H�3av��ӻ��>�ݳ��dzj�����=�)9 d�Jϫ��G�%��6���r������F��)8��9*����♐�fN�����3kG_K�cε�1��N� n��S���$�ѓz��#�/,�vMf|W��d��A�%ܡ#|2����:Y�k�>i�5?����V-w��>Gڋ���c#?��w��!��w&b39_�<���:�&�<#H�P2���|���)��S/�c�<"Bޭ��8�p�іB��m��rwt�>/8�;(��L��O'y�A�[j��5�y�=�^ð��.l��Q��I.�����:6	ac��6;��]���2��(t�;)�^�S�˿��%�8["��/�R8>��j:hc6*��#�N��WV��l���R' ��<��%�L̖��kGÒs������(д�B�#�T�8�9�Y�M����/��M�)�����F���ӱ �	��o7�,���y3ER�"�'��N�#���S��]���
<'^`�&�`�Q+C)Fgx��M$x3b��B
(3m�\���J�	�Eϟ�`��[�y4�������a�c��J�^4���G-�b\�`����Z�<����5�Ww.OƑ:�6^�f�ϫO%y�Ч�=U읩��\z$�>ٰ��tW�4� �
S�
=�'�I�<�}��r� ��7�	�g:MT6�����}R�3�ņZ���7��L-�dL=i��=�v�����B�Q��̏)���;��^��CH#�ʶS`+�FoYܔ�0�Z=w))��RC�j�I�?iaZ�N҄�o�
2�d:��cNw�5�>D�؃���R�I���8��!�C�>ݞM��QrH�&/�۶G},h9�����+_�R6���A?p��G���Y��k�1��K� �r4�t��ⱦ���,��ul��
$�Q
��C�+%�_�EE@�p�u�C���A?'^{(�a����X\����f1�F��<�. ������B���ג3�Zb�G^M?�������)Gt���Zr F���ɏ��.�>�����0,Y��GD��f��Cf��C���O��� l��I���"[���Z+���"h'`�+�'��כ�������ع�e =�*5�n���P>�*8v���B�:7�w�,w+�',�[&M�C���ꏁ��`d��!���V2��/������?�E2�.���������ٟ��Ҳ�B��Z���|\�͍�Jd�NP�9?� x�Ȫ̋�l�Bp���Lc�]�����/d67���Ή�ɂ� ���,�ɟS���!�3�I�y���0�9,� ��wf�7��o$������i��A�6?k��S�I	B--6?Nd��A<�T��X�,�ȪGk�� ���� >��="�����p�"���[2����7�-���/��zGa�o����D�08��s?��v�=L9�hx��[��-�J��h����8ȟ����A&�	�E�ҁ��n���.'��X>��/�^��L�V(l&��n�u����D�)�D�_B�|҄0ְ��wv$��:��ġ>�
�ґ�mԦ3|?�3��jT������/5*Y���F�������SPL��U��ߏ�%%������:_�np���b7k���=�zOޑ�����]���#^|���!�J�N_��i��ށb�;�.q��}4���_�P/I_D��_v��|�&N��+Q�t�u���<��I9�R}v�ፖu�P�}�o p����%HV�:,e�x@J��[x�@�ܣ�vJ����F�3��B�!B:���1�YA#����p��]��{3�4/
����9�2���V����}l<]����qTj��������66[��g�I����i���>C���Bw"S]Ţ��[҄V;�K�DF�*����h�iZ �2h��kL���ˆ(�Ø�K���ٔp���5�� V�݂�|ךs"�8��.Mw�T8�
�Y,�p@n���eޮ���]'Ŋr9�a9��V��Y�v�K`�\�G�
�D�U
����j�b�ǃ�Q�_j�����uc�$s�dZ�Ƚ�y��`���~ı	@ʇ`l��F�7e���N� �&�wv�
����2�@B���U!;�A�.8���A�FIA�<�u�����X�y��< x�/�@�[��+6��JTX�],;\%�O��iA�T^z,���!p�[�%�`!yȗ<,o����K�Iò�C��&�R�:��v��RYMԕhT�#a3)+M@�cT�>l�B]���Gsj=��v�t#��$��&;���,�ȇ�����r�	��4b^[S�R]��ED�*�.#��x8ھ$��%n@�Ll���(��ē�W��|>��f;mX�[�d�	��P/}�=nr�jnD�h�t��D�O1�ݟ����Y�T��SъQ��?�_�N�-�,4�����ۭՋ�����PK{^��[d ��Tc���0y��:K!ʈ �hrC����'�m��v��q������Xa���X�\�E��wU���j.,�)�%��5d��d��!iFzq!Jn:"��h�"�A��v�¼�*���b��c���1��+�z���j� ��|�YS�uM�] "��ψ��e�,���ws��Q4߷��K+��(��9'2X�`�D
+�[⣻)u]`%m��
��fø^�E��r��J��IR����X9iKZ�bd�&׉'�0�\:��pb�D�0�R4����&`˼ۂ���Yחo�Af����
�,+�-.�'J�^16Z���Sy���yU.dd�!�VF��{���MZ�{f�~��c*�3k�&��Wl��N�'�͏���1�P,�n��r�ŪH!�t1��`�=��^vUJe&�EG�3��C4���7{������r��)���r�WX�e]��:I3=J������vk �L{�Yh���u�%.{���]W�b�}��س�[�7�Р��\������m�h��@4~�|%!=��F�j
arlbjH��G�v�qұ����[�#-؈���o��?�%���;�S.-SjY�j�e�K����$^���]��6!h��A $�d��ؒ���o>�d�驯�{�������{�▋�e��,�\mŹ1`�j�iF<΍�Q�����og;4,���5����yyN��u���]�5��S�R;������D�/E䩢�|�f�g���&R02�U�a]'l��H� �`��yu��ȼ���n����Pֿ�3��o%��\Hw�ِ�z^C�F�vhd��So���q.��j��C�����M�n�px�7�e\uT����o�6�,�t������M����h';�� �.�0	���?����n��n�;�ua�e��&��8x"�����UB?�Q�:.e7b���=��z#�@&m[Վ��qSSO��bv�_*�76{-�9)EW�u�����U�C5J��JR��C����	���Yʶ�X�K0��.��rGk�N�=�B�j�)�>��&�^����:�	@��Ʊ�B7К\�@9Fa̓�*t��"�Gf��%b�8���aj]ل�tH�˅����|.��Ѓ!
ӛ&���"�A� ������<�r��|<�y���j�fR����擬i�R�K����o/��|@����WzBi-Q4��}>l���͒|28�,�G+4����T.�-m�!H�S��W��r��0z�;tW���ϩ��~�e�JkiǮZڵ���3�*�T�A���K�[ݰ�����zkgn�զz�E
G��?�2)��|�1�rП���1����N�M�"۟�t��2|�_��LY]��N$��xC�
:Z��k���_VZqkP"s��O��כ�DC���n�wl�1��� 8��z�0�'՞�t�B�蕳�~��J�<I�uz��	�����g��`J����`\���ϻAٻ�F�FUU}�4�C�,�8�U-��g�l�l�P���S6=�HR�{^$���փH�:�H��nķ��tɶ��JdP~֨a�����@�Ljx�ϓ���/8���t��v%�PVL�I|�<�����pɤ[�.%=����E�u��^d�s�4�H-+�2�ܧ�߁�^��A��QHFU�f��ݪ!�%׆^�a�s:�teV��EGن{��;����=�KԂ��aN���=#��u� �e���4�"�zZ-���l���F���x�4�GGm!�γ�C�.;�y˲a�'z>k_�V�'�:SĻO�/�t�-}�����c�f;�#��E'2�vl#����|uh읋;�83�;�(����H����#W��E�4���]��6��ʧ�%p�x��!9-�-}.��%�ai:�c��}�K��3�/kC�P�[x�N���6Q�m�\�w	��Hl��InϴEga$4��X@�\��s���Q-� ���=�{�ػ<`��C�xW)
�/�7�F yI�8w�'+������o�Vנ�d��0?�C�V������*�T_Ȣ���S�E�������5��{I���N⌘��J��<c ���-f��=)p��=�Ж���^:�̴W������h�YL�����ǖ�Mh�K�*2�l��EןC�I�� <ez���?$��JS��o�=��s40������InR\�֛�<��	qmq��]G�fu!"7��}zO.����_v���qX���4���t3����Ԧ���3f�?���+���qɬw�-0�<Y���xwvm�hU��� �u��y�I�úa��x�3���:�����hkJ�4�ywX������e�tn�!s�T�<��ccm�N
��Ee0�OJ,t�ƺI2bBL� 0}q"����?�4T���D	��y�,��C��J�N-\˔4=�v[ڤ8�Q7�)Y��7�j>��-p�3��H�:w����p�ε���R[0�ɾ�kd\G�o=�C��U�*�E�W� U��[J�	LU�[�F�mk���4s�O�������*'*�#�'nO�����g��F�nQ�(?����m�OfLЮ�I��X����5\w]o�䙬X8��!q������Ol��«g�o�=D��ql�I��<Q����X�8^G�y
7ְk��G<be(�@�-�q�H����O]ܻ��Kք��drIƖԢ�����@�uA'�[l�/�R�D3@RU�N�6��NA����8?����݄�7��<W�$�Б�X�Z�v��D�(��Y\�" g�'�`La�Q��4]�v8�r�rG�*�(�^F��
k4�������)��n��`i�;�C�u�[���2�tƕ�Ҥ.Ji����O�^vXL!�淝�>�l(ԥ`�D}�`����{X�3�wVHz�.�^F͸��UrI��̮ۧ��ݭ!\�D��©vɘJT�TQ��7Og �̹DK��v� �5[�L1�T�;B���Z�S�ƂVt�}�Vb ��YkHH��k�'�o���R�H�<�9]���I��t��:�FU��ȴZ�CSJ@.�8epo��[{↴B�ƒ`(J*|�[Vw���������42r":H��/wZ��*.�w�'��C@�~oq%����
����T����gx�C'B��X�ƿc�H���|ܧ�򗰼�Y��d�_*Åb��5b��e��	�
2(K�}� �(+��ޯ��X�6x���p�OQ���1�� ߡqĜ��G��G�~.Y��}�(�@�j���?���_X[A�엢	f�P�����U���z3�.�ϊ@�*2��-�$�b�s֛4S�bg�#���	h__��c�i��sg*8�^�����S��X�y���L6Gd�e�$������N�o�`��#X])����:��#��i�`���X�dЙ����G"��"�JBK���;�����݂�pO�߫3�oa,��ƒAzE�AF���	=:"l%�Ϻc#z���V]�Hz���(D�G~6�qSS��r��kC: 6�*�ե�7n�h�n�m��̽�
9�z6�A�fo�	C� ������9�<q�X2�Z�F�o��z.���ƦF�o�s��u�����B�a�W�ei�6�N��܃�����C-���*��$r:k�F�~�N'EH�M�.��bT�u�ƒ3B��D��Y)��4�Ӥ����r�Ssi��g-o�6���7�9Ͻɢ�����,��G�K)�-z�0FP8���1�%�=�mŒ"e<�^��%ؘ1���?c�7\C1gsn�oj�0��&o�����^[Enc��ʭ����dq!9�x�N ���T�$!�:�T�g$0��:�&��⦕9�۪ԫ�;�..1.�#�I��1O^$�Ȇ�W.z-���|��5rMJ�W�@9��2�KZ�~ǽ��Ϩ�98���i���� ���k��>�,��(�z����eռ��Ǟ�:y�G7��$yF�t^!Z��uE�����I`_ip�g���k�GX��i�Ŗ0�J�ƪ��#w�K"�����1<�uA;�������|
�^v:�.2!B��'6�k����?%׊�<� ��|"U�z�z$�?���RO1~�F."�~-*Op�A�J�%�txzd��_먅�4��yz���B}u<��dE�e�H'TOe��
+B���C\:���.4�8&�J	�2���(+�>��ɠik�^�85��^�1�_I��'���Z�AZ���t@�,�u�y(����T*@�x���h�BUJ�;�D�8�Y�5�{���D�)3���h�T��4w,���1��R��Y}'LU�l��8��s'ؔ��^�f���"(������2v��8�U��`S���E�ʍR�:���G-�"MIЌ{���HD��g�
|�������`�	��l��q�LP���An�Y"�-��&E��٤��r����v�1�Ȕ����%,n��`�T��~؀�ھ	cN�����+_��V��!�ô��}Tt"0��_�C�<{Dk����ӿ�~f�6l�
+���E��QX�q��mT��H�V&,��-{;����/�!�vQ���5z'�5��;�'���[��|�A�sw�-c��_?ѱ��+'+�f���Pr�3�L}�+�)�ٱ͆�TE<NFg�
�Z�mG�/�4]��P�	(	�E=��c �!� U�Z431`һ-�C0�H��gΞ[̍��O
:��f�a�ƪS�q�7��A��Z��VP}l���O <D�:̇V�?_�j�� �v"�Ųx�:�N��V�p�-a ����:ag�4�N��=#�����`6n��/k��Pz��Avcke\"��:��
L��Vq����uOo�N+��U�U�>��r��.���1��G�(�H>8���^�Ʋ5�TJ=�j��4�D���eJ�5v橄��E/Ysq�����,(z����ij�_�h�<��wyz4�]�AA'�^�Hg�6#ǐ��e]�(��Spw���.|���Lc�
�
�ߜr>i$�3����[6�R��Yk�P�&^�}Q[R�d�u/�ћ(������>F}N��uT��0�Sh7�E0��,F�8!ǿ�b!
#�9;�J�� �ֶaU��w�:�l�n��I=m��9>��X/����}h�ɟ{V�-�yN]��;�۶����}�7��s����L� ��t�j���y�qT�,v@�xl.��4�)h\
lA�ܻ��:aΩ!���(p%[�$��W����d��*����n������	���w��,�(G%=4Ao����h�<��Q�G�u�sn���@���O���W�C긴�)[��'a�I�2�q��`#�mO��-�]�t2Y�/؄E[�=m�W�w=�����f�#���g�Cr��l�Gɦ�ַ�A|��/�)2`�"�)5Y��?c!�����n�	�� Nd9�G2�*�%	g-F�i�Ф�Ų(U~󛞓Wٝ�J�ș1
���K%K^����fNg�,���-�8,��5<]l��$֪��Fyq�~��tmI����H;���ۺ`v��&/�� xj���<�9�5�^�-����9�Wò�'χ~�����'**�/'1��-�x	m.���~�J�Ȭ�Ai%1a�b��%n���:'o��@�jH+$�[�<���\*��G�>���,�T�f(�řm��u�+��+`��FNh�s�aoiz�:��"Mq�VI]�� �Vm�����fG�,o�J��	/��O/T>=I5��&���ǲ��e^n��� �#��b�B���t]5c"e3��ǁU�;� W��-�?�����F\{�Y?6W0�zh�������Gv%	�Kl��Ʈ��d�c~�18d���6w����~I�H�$sm��/�|��S��--����p�[���ǵ�^������j�Z��h��`��N��}"�3�R�Sǐ
m~Ʌ&��v��^U��(�WMY�+~��^�v/.�"�(��2=�����}�U���Ý\]Yß��a�|<���!�I��6�*�{�ӻT��UN��}6�f�˴RL�k�MA(���~��9�>�8��ҖMVƙ{M*��'Z��h��T~|����v�~�4հ����� ���ZY�a%���iێM���оkk�t�J�(���Z���J�S*����w,�z@����q}�Ա�.e7�Rc�Ol�;�"�c���-\���Q�����On�OFO�>$�Җ�{�����P<M��$*Yu{_(_�櫫�>�UOa�ך"�z�r�/�.Ϭ�MqgF� �������;�>�X Yiȭm9Y��n�>��Y�;�$Uu#)f���85 z�����,[ȃ���������1�����,�|������]��ti���~X��t�����`��᳢�K��OGly����tV!�~T��ܵX��.7B�z�66�+R���οj%�؆w�ݡ�$�rg8��3�q�QA��=��w9������B�r�t����!��Rb:����S+Mֆ~ˌQ)등p:�i�	Ȫ����t���N�cP����&���ȷi}���Xs��u/.qE��+�.L=�i��Z�_��w�T?�mB� |�EO�LZ� y�B܎��C�k����Iî��½�h<ڰ���X�C��p\����eBF����©���P��=%gAs	��&I��>A�Y,�{uo�^q���h
�\�dᬖ�7�G
�9� i�l���5ܕ�G�B��ښ$�:բ0�C$��W�<\�N���~I����v�n�r��*r����ȰNW֜���:�)������8X�h���T�A�8[�|�lż,e9�y�ƊC�p��y�,ʄ�����`�RT�U�(��7�b3u���ro�Gc*%�A��Md���
�,;⡻�m��CYݰ���_�� `��x�k|T��?�v�������P���r�|H$w����D��3|�|��A��C�o|�诨�N��<	��~�
�9a��rfn�i�a�k��˼یOf��
�`�����D*/�����۩��k����RK��)D*��Op�֝�=p����:2�px<,�ᆈX�y�ٜ�^�����W2Z��X������?��m���_K��V�:��9'�������4���ϩ=�;��V��\y8� ����n���.ˉ���}k�,��݀�1�	�Ô�7�$҅su��ڃ[�v踞!,�Wԯo�b?�A�箯H����J�H�}i�#�u�Y�Z�d��z�J�Q�B�|��>[W�g
G�d�ښ2qn��\���(8A���A_�M����O̑r��� ���l�#B$:���",���Ր��;g�.[��
�njF;�#_���p��}5����hْ��@�'�oY��&�đ��#Ż���D��8[����S�-����& ��K�q�Jr���b��������˷��j3��ߎ��ܻgCM?�P#ܑ߬a:,�	��7T�@���q1
�|���Ҹ6+V��B@���B�ߕ�͸o�����<�i����Iܬ4��3�г���b�:{�ᢸ H����80xR;���{�δ3
+��ն&:Q�:�ZWǜX��<��4����!,�i��PH�� ��+����:n��s���:��=a��/Pq�(� =��2�3��Z~E���$�R��Y��Y���9�[��i��vk >Uə�凟�`�ԓ˒�o)G�!zMǹ�8��M�|�P��]I�1��\����P|u*����YՉ�1Wl.}/j��6��R*��mk ���#�n#�k�nާV�ۿ�/�� �֖Z�o��׏�������G<���Kgl��рt��+|���r���	�wU���>�f<7[���5x�Ԣ<,)J�jd�R��1��jHW���>c�e�N����%���I��k�x�!�ߩ�5ȍ�:�jk	z ����Ri�pY�aڞX�5Ǘ<��{�~i���
�Y0Ǉ�?��>caPk��m3�u��c4D��IN���P���T.B�з�V����-|">�,e�7o��N[��J��O�������;�i�sk$:o-5W��Ƽ����hg���Y����Q��dU]ꆏ�U�l��FE4����n�*v����4T��evM.����@̕OB�_�P�#�b��?�	�.󇇝#���At[��@
n�d#~(p��B�	'e˃�]�&+'.�7sc�x�Jq �-ٕbw0��L"��U�� �ߐ�	��T��օBI��#RnO�~e��zo�r�2���)���2�'[��Xc�t~l@��a���箖)��^�[��$�x	��z_|�V��"jk`KΉ[O��_fx���3�ĤӬԒ��S���3y�	�v3<���aaA܌c���(��m�q#GgwVt�$��,�e�ͤt0�З�
�O�nu��/�2T5<OQ�s�~�Y�y�e� )�Nl%�N���|��bu�{/�edA(���2*ųl��e�#q��2��5�z�F�An��.�)����=�V�*�cTj3���8����o>	��?�Fj	�j���Y-�f���W�"p2��4&�f��O��ĤR�]ؚ��0(5�gF+Z�;�}�p��ۃp�u����V{|�k�'t�D�&=��Y�?��@�R��Zǥ�xJ�����|�́C�Oh�r�_���^q"P�M��ZFT���s��=F�����X��U:Yϳa̌l�O��;�er�ӄ�%r4�̉HO��j:�W^����_��_(��׏���������C:J1?ݓ�F
��p�x��I�ê%Ǡ�#�ZR2����V���u�D�F�9�$�'bm��M1�ñ�`-]��R�P}��)	.�v���9�����3�ms҄I��v��2�FF5[\��lh�u��x�蝦�t��ߖ��z�pRfE.�O�ƪ0��>���+.	�/����8U�?�.��<�E��!�DF�bN��XL��ޔb�t�#w�鍈�p�%���2
�%��Y��V�B���C���)f$����k��m��KP<�����H���)	p�� a^{b�B�p15y)��ݸ� o�@�;"�X_�����A��J�NT�̈́1Gm�e��,;u>��=/���d�el���ֹz|�����b�s�.�xF ��?L�m�*������$��S�r�8mPi}��\o�_ޫ�;
��2k-[U�`3ٞ�O�������<��e"�ܥE�:˫n�e�}��K��1d����8�	���1�M�_4�^E����Y��s+zTh��ǎ��l���AY�Fd2��9N�o�b��ٗX��?U�XK�LI�@œ?E���e};V;ڑ�6���x̧�4ص�޾��	+���]Jx��6�eΎ }�c~�4��r�T��9���cF��#�*��&L�Ag;�K�؇�H��D���aw�YC�'�����a�71�iW���X
�����_�B�3�4UOiձT�n�-����FZ�D�q%��g!y�Ɔ4���9�WY���GA��=Y�ֻ֚k�6ٜS�/R���/L����u�h�!st���.��%$)'���N�䍯���~�a�Φy�<��<&;��E�'E�c���6��Ą����F�U2u� ��f�]w�i�D̘2�e멠ZT�@�Y���(i���ݺ֜��흓�ۮ�xm�I���U�E"W�ì���{ɥ-�68�KdCN�e�0r��}��G�ښ�A��ߣ؀�B��[b���
D_>�BՐ����_��9p�r0q!&�"�Q#��,��M��=~2Z/\���|?�e��:���!IU�^�0G8�F]o-*|�E�g�ƿ�Th*�e�VU�ugb���jmQ�\f)�n��$�P�ʱ/I4.28�(x"D`���p�~M���-�̡5)�j~�����4I�1�Ǌr�B�"����
aӪ�9*P����u����:ʠV�f�]�B r��$��F��H<R�\��;���\03��} *�D*&Ò��Re�q�u^�@n���li|t��E��"X�����G������St �=���_�"�T�8e�a���Ï���[c��ᝋOTT|o^�"��\�Z����Z�;"?���a|:�>��Q��L<e�����-�=�*_p�x~D��QD��/�9��h2�x��rQ7���/�W�;4"Vuo��jaW��[j��2�F�+�&a+-�](���a��_#ԡ�`��JM�pz`��-��V$�X� d(*��&����4s�B����:ltz�qߔ��l4�2���p�o�^\p"p��+��Ҿ���B�;��� �Lx�z�ԫ�3�a��"��i{gNJ��S������:��vO�)��K*�S��{N��n>�6u�w�m�̥�Rt �����x�ͥ������`< ��DŠ�����pn�_U�>y����6/1/��'a�F���-��y�戨�,;oSx�Z�;YHE�vT-^��>J�̀�J��Pܫ6��z:8�K���Z3B*�P?]�P������G]+��GB�(�{�����e�k�}��bZ�C�bQ��k�e���F�RA0��HJ 3!`ܩ�V��S>��<B�q]\&yΓ\��3A=A�n8�"�(HV�h��M����xJ��b�Tst��׽��sL��q���.��y��V/4�
����m���Oʲ��4.����v�_L� *g�8��j+��X���o��.0��nc���ʦXx���A�]2�d�~�&��=�J�B���t�`=6ޔY�W��%q������p��;��k��U��=��Iԅ��Cu%RA��,�Z�ļ�+,ag����S��Э"W�f�Jm�Bd��{�ب�fRc�&�߃���ɰ���h�3�P�6
র�Ѿ��`�U�Kp~��15�0at�-�	�
=>D��uL����C$"��c4��Т�J����j��,��(������zi�w�kH�ۅ�\	7�G�+G��n�ػ���8�`��p���rsi��X�/Z��C� ^�}�}ʟ���>�WO��u^���]�~9�*�@�j�0{H�mq���vB��0.1nTn ��a��ґK�:�Y)��\�|Cۦ�dKRD\K�ى���[�DP(�{�4�kl����d��M�5�+�<"F)���A�3�>�Y_g��pE�`hY���Qݭ �d���V��b�}�4& ,*z|%e7�9�홨�f��ͱR�|��_<_g��K*�r�Y��#�_8W�$�� �]��#��<���F�&���nKHι��՗�� $X��O�N�=���������$��)X�)*Q�#�D��ό�ʡ�bR�$R�����ڇp���J��}���Y�c�+/ �X0*��TgXI��3��d0-2;������_�h�wz,��ݲe�L��g��#�>���N����3�/�8񬍬���z���4�)�bF��/vsd�C35�P�&�H@?p�	�"����l�G�Ao醚F����mVz�$\8<[�F16�ͥ���g�P��*���\)좮�M]$�G#�m��T���S@�b#��ϵ�S�}2��?~��.�o�K��K����l6lo��0a�Lc�2�BX�i���8?bV8�����g��e�l7�r� ��R��ʻ����̈�_"�GZ$~c/�?�}���WL������KM9)d�[�����ӄ�\�Vm׿�ЛXg����2�,�\��X�S�iV�2֬W�<1F����0(���􂈐n���ܵE3<��Q.��+�D�����8��b��J���i��:]���@� ��4�d�F�1��~1Ѫy�^�M���@]]R5g�Y0�2���ǚ ���"�vm������D���͔G�*MVL,ˇ�?����� �÷�-���������2{�Z�s@ Tr1!q53���5��o��;�C��Y��S]ɫкG��ŏ��=4r�7 ���L�{�O+�n�bY5�	�䅭��P�Gu��^��ķ��*mk~	�s?��$U�@B8-��H}����*z�WXY�E�-W�B}�ȋ�z@S���#.�Dq��'c<���ÿ�oPhH��Kb�������&)7y����!��洐����l&��z�l�@u��4�[�������'�8$͆g��Z�����㊰���Ay9O�:�Y"�Σ�ߋ�aB�0_�Vp�5ܺ���k��A�W0�2�һH�<�T0��1F��ld&U�X�3�hO� ��c& �J�c�Ȭn�� 8�B��/�f{_�}b97���H�#k��[�t����a��{}�l�V?Pg�б/���g�Գ{�|���U@�c�#h.a�+c ��Z��t1��8�(��7g����e(ؐ����a~H-��,��:���-b0����w�W<��
�Ȇ�����>�<��1���S�j���E�Te;��=�éI~��P���T>gK�"%�Ê��{J',s�Z�n���ke3(�*�Y�-�"5��MMd��
31��rv<�g�}���Q������~����'�;����G�c�1��=� ��'�eJZq�����'ڬ+U��4y�.AA���td�5�4���x�Y���c}��A��� �w��~�UDT�}��(�kV���I�$�2�s�>3�>_5��GR"��5��K^F�s��j}T��È:���?�w-|�1�<M�]��rb�I�����L�$ǎ¤�ꄙ�V��'�\x�1:�5�XB�p\;9a��`���RG8�)�a�缄���f�f��SB�$ߌ��7T���1��e�k��Y��!di9���Q��ois����\a'[�e��د�0R��<$�������#�h5k!��i���qmD2:�K���F���rR�#в�c� �{�XI]���Q���9ޟ5�G!x�G_����ؕU�ق�?*<G���0r �� �W�^yd�=w�8�R�Y��]��ܒ����c�Q՟�K����$����)�E�kߗ�u��a��mM�m�����p'�Y�o�z_E.� ��p�W��eoyO��K�5���bzexy,S-��n�y�
�O�������k�4�N�F������������|����t:C{���#�KqVbya��M�N"&(�� �����d�������e�\>d��o�
�y����Pk�ݵ���_�>���6s��\%�J��%	�`��|L���*Ó�1�`%�Dʸ?����M�|ְ�z��\�|\Ҹ󨊇�|b��`Wr��@�)�j�x���-�鸉gq>�Sy�g�=�� k���&��k�ׁ�U��q���'�U��ǚS�V��J'�ښ���B3��&L(�
��͎�z��@
���gP;\�t�0�H�z��?ʤ"�.��v1�Aډ9�Q��"������F���S��U�ytȄ�?�0��3e��)�#e ������ݤk{�8�C\	�˻tL@[��A6�L�*�Q�в,̈́��s >�g����C�m��x_��r��{�Ѽu~�xO��Sl�	��,P���*�q�D�#���y�;�D ��|~2p�n5��K-`]8A�-9+<Վ_�J_z3g{ب�&*�G�h���	M����z�����'M���,�f��Ƅb��]R�� k/<S�(͠ļ���H%F����2�k���Vc1�t���m���d�OtYT���Mu8$[�\e&�2�6���G�B���q���h��U�� [���fQ�z�E�0�f��C�mp��ёa��~�Z���TA݇�ݲ�0o3ǟv8���T�S��#zצ���F8"F�{�k�/Mf��S%/�u������X�+W�S]�ȦO��+nE����rr4�����M�]��l�آ�W[12��U�z�	mR��p�P�t����Oa��$��^ՐG0�,�#.�QACgd]z�D4H'����+)�S�ZV�ȡf�9ʾ��/�7I6!;{�
��{+s�'x���C.O��&t����Re�eBJ��v�|�R�AՉ�� ��ϻ�0e�}/�48��$�4�Hc�Cb��b��_3A��5<�@"i.�[L�?��~�����;W~�I��s�\��Î��D ��(��'JR�k�\�0���T�Uyj�K�:��'Y��	��@\q���(�$�	Q��z�J6��V=ם�ގ&7�x�QYE�(B�_���:L�k�)�n{H^X)#�'�B�eXʍ�\e��d�D���#���	�,�9gTP��b��!����pέD��f1��f��*�-)��eg,�!���bd��3�/�L��_C\�Sd�cGtg:�i�g��9���ߣ]W>A�:�#��A�X;�QYS�Tn�4>��͖-��3�-c*�Q$����� �B�nd���`i�ҫT���$~λ.v�i���0jI� 6�9O54��|�:�ҧ�6$T�"��Ö"��`���H���8��}�2�o���ν�_�~yC��w4�=���2`݀�aXKֺ�֘!���B��j��^��Ξ; s.l!�D�8��%k�VJY��^{�PGQP���bTUD.�`��y*{�v��zp����;��,(l�7X_(��(��fՐ!�\?��������.�4c���Մ�S�p+�]���[鄓��8/*E�{�jdUF�A�:4T7|�r�x�չ�v+f?WwGV���ㆮnE��.]�$��`� �w��������r�<0ӭ�7�/�@�0܈kS��(�Ґ����V���ef&�Pj�~�+��W��rIo�O��Z#��
?'&�Y��~V���q�q>���q��5�XMTS:<
P��x���3��.�@�����e#���-/�Br,�;�: P/  @��G@�Qg�9����m��m�X��`��H�S�K�F+v%2�OZ>�~��M���ǯ���vyDy���wR�+�Z����yO3	Vl�2jǹ��N�)�1��E#���^eCO�)��-2W3 K��|�*��ٹ-+�k0���M�⭘�֕��Kqϴ`6����յ�ø�,d �5����)-N�&�- ru��V�(�wxɹzQ"�ԯ�i�2���mO
��
O�������}=�l�.F2�����'�f�9u��u�7����Lu�:�i<�)��$\h0��'ȣ>��XQ���˾�����ޟhQm��Z+�w��V\�`}��4���elQK*��j��X�@�� �b�Б�7�5���$�7���e�:��K�%��snT���G��M?��2�C*nZ�:Դ�_]�v�q_�O���d���ic8ؗ��A�=-k��Ed��� M��(t#h(�`�����I����B�ꗩtc��w��SXLE��4��c7N��佊��J9�[�5n36�o�o�1;=���߭{O��0w�LI��ܨ�!�?&��c �5����U�mqV����ҿ����>�r�A��q3%xזFW`5Tk	��ѐR�]�&o�s=w�2���eW+��@�J���E��ٞ=P�39�u�D��Ԏ"g��R(��-ZT:�w�V�,JhN��'>�J)_yCS�?�RD\�L�:.�u��n��:D���܄�f�&
�G�<)fGL��eĳ�{)�7��u����Ȩ��o��Y�n�w�Gk�ă|_38~?��l4���E*��>��﷬㋣!�B��m|��O��J��V���T�6͔����.9_��`���VwZ,N7���'��ir��yo%�0�������Ͷ?7L��q���#�?��uZL6�"-�_���
��T��ܨMR���8a��x8_���拞����H1�јt�c���`�)�O۠�6�w���!���ī��A�T�E�)���<�|^Ʒ�Z�PX�'��7�nPcX�-(ی�M���γW1�[V����s]��i{�yF���q��|H��;���5�|�2�����d�n}WM��"2�8�����oR��b9�OժO�����б����r���Ll*,ұ؜����2R0՚��S ��Q�f3>�O�"4> �\o��	�;9����ҧ%4#��]��U4���[�)L�$��3(䷌'M
��TF>x Z�5)gTB� \Gi��G�ME����wQg�=i<��΃�־���������xZe�F��/т�m�J��L���hy���H�Ȓ%����l�s� �I��:�I��RQ��'� !w�N�s�v�vn�
�%�i����P{d��CM*ט4�M����r d�O�5�^���Blf�eK�x��_vڿx����&M����DöV�[�	��9i��P�']:�v)F�{U!��p����M��< �� ��Ȯձ]��*��(��N�bQʜ043�LL!�c��:b�)Aa�I��d���qн*G��Ue��v��!��#n�gRǝ{��"��A��pŚT��L��&9Y��+��R_�ƒ�<��?�V���ܼ��U��ozϪ���˦_����{P� nd�67.ʍ�Z �,���i��_',�L�?iE�>�1c�g��Ի�")�M�J�]\�AUf��Ֆ�ށ ��P�&�Z�_�[ �6��A+��>��Jm�墒�Go�Ad��<J��4%?�����Xh6�;E���6��t Y_���$34X�Ѯ��IhCϰSC�2;Q�ԥ^�T�1EFT? a2B��CL��O�g�h*r���B���m���iI��v���̊h�j?�v��X�0��3;�./���V�ƥ:򱌿�b̡)]vp ��ȝ�X{*�>v�@�N�kQ��T��01C���p��0�\�/c��僆�}�Dy�7̦	�Ғ	0<¸���-�J\_��1��:DR���	ju: 	��k6�Dn�b�8��r�V�T���I/e���P~c5��3��V�zȜ({Y�oC��y���Mn-m�O��w��BM�s��@'Ǩ����u���T�5�t�Kl⩾g��T���P| �ϸy�	�L/�-[V����Ӊ��)�ނ}r�O���5�fh�:w�XD�C^�ݿm����'Y�)r 9=�S1�OȐݧ���qY_<_0��j���˩�lރ���\�E��j�|%�di�����d�����|σ�,RO�̈�]���f^�z�Z(��-�.�	jD�Z2�PP�r.�5�F��}���8#�(Gh�ͫ"�x�O�J����^Ǩ� �-�#y,n{���KJ��[���G�ExjS<�PĴ*鿺p,�ٌ�+�����t�2�b(�,��u�����b"V�Ք�b ��L�U�c��cZ��r�Oˀu�6����zQ) ��2,STS�k-E`q2��
*�0C@�=U�/˱jC�֚ud���I�4��;��W�#����~�R�s�C'PM�:1��������K���0}ί���fg�M��8��t)ڕ)���?⭣��%c�D+��~���{��u:�u�jA���<����� �1��O�r��xX����s�&;R��˙��#6^kk��2��D�飯���"IO'fKU$���k�"�,5��ɺ�J�\_���"@��c�t�[��(��ŉ�qW�dw�>����+�z$m7�q��S2{m7'ɳ-��JD~�����@�D}K�te��ɷ: a8Mn@B��T���+�X!ct��4b/sL%��[z��'��%\���&�̼ѝA��?mW<���k	�~���42��������l�%Η���XE��5c���]y�6	��!�piV�V喍���杗���[i�л���zx��sP4��'����բ��|V�&U�dG�t�!���G~S�Aٟeϰ�WAI��FqfO���I#NzT�v�k��wnF�CNǯsB���?����A���La���涐ۓ�Q�YCPX�����	�ƴk�;�M�A�E��:�m�b�| ��}oiq��#Z�XCs��ϒ�Sh�H�\'���R�ݐj�d�̩B��?�e��~�*PS����w��8Ǹ\�L��T:����y~QƂ�R<�x{"��4��$<zw�zg����-����°�;�N�L��~Z��q[��sp����8�-����o/���f�����W9Qvu�$rB9�߁�;u�#�S-��O�Y��	�}�]��.Mi���w�u�=lg��cERvXWK��$W�k�"Q��pt���)8�����A�x�gr.���S�W8).x0K�8�|J|2�驩�Q��jp���,d��g�F�o����^ �L՘(�Q�N
�v��m�- o�I��ѯ��.J�C?�4��;���tb8�j �T��^YG���L�cڕj��57��__�;(�%�?�Y��U�Ӕ�$+>�C6z,�5��!��KZ �u�L��ONRMN��;��L
K�b5��X�t,�&j{�v��x���q���@�ОL��|Ùar�������C��mr�ݗ����Wy^ރV���1J<-�i��O��vv)�!+�\mu����h�!����(fO[g=d��U~� ���vc�sE���3Qg]�%ы-_��T]GΌ$y�#>��.�*֨=Z�Y#6����wU\_0��J��t�?GZ�6��^"�zN�K#�w�D��f���T�}�����/5�[_VYf��w�|�T�˪����6�Y5CLy�����pU��m�'�KF����u��%�!�3(�9Ns��		Ï"�����h�ڍ��Z\��� ��m�6J�n��������jW�Dwr3�oV�F��-8�8�s���Uw��)������O�!����w���2���R@��dd�v�T]�Hp�r�,���ʜ���4иrTV��S�K�^�^���4>��-(�R;�6�]`�8��J����~#�,y���<(C�ƌ�剰��8����VR���SW��U���i���#��]��/7u`��)[���M����e��ƫN �/80 ��Xi�|:�ڼ��v����=!�G�7;��6�� jJˢu�sľT4z�?\Ph�@�d@F�.��i2F��������>�2�$���/h���i��FMx2����aȾˢ����)j#魴����Iʂ���	BO2|�Y��ue��9E:�T��cV�Q�;��[�ͷ��y�8���?�U4ofb��m�J�n)�Ĭ2�})�M�#��^?m�W.
1(S۝p��_~B��G�
IW�>I����Ϝ�V*\+EX�F�q�֪qOi ����.�
����H��Zθ.��C���^/�_�7�Q�=�&S�L����e-�_h��f7��B��TbV/7�<~VtQ���QP��R-��įΌ���8�g���Q�<R�%R�+]�v�9��ϭ�nhx��Mx"���`�0T�n�a���5�(-������Z(ړ�������ܮ����yv��L|��e�Wt�;��.�jv��Oߪ��{��3��F?�.�����ove|�e)@��X���&���;LT�X�K� >1^X1;��_�Ϧ�)�6�D;��85MYuT�9ڈ0�쒄��wU�g���4x��E�nR��w���99b9)>�����m��|CO���O�{�	[
=��������_�&~��DO\��J��k^n�s�#���G5�_xT]`�l�LX}�֩�?�?uA?�F9�1D)��!A���kw�r����
���(�*9#�"�E�n~@�`�8��*� pw�H��%fZL!hָT�<@3|�����`�{����-*%(�'��z (U?aAA`�g�4x4y�С�ϪG7)gAX?y�j�S���-���>$��LA$�(.'}��YհU��/;�G����L�.ĕjĳ_o���D����}˟�0���N�jp�Խ]���۱�w~W�C[�ׁ����s�M�^���+�"��,MJͪ@��t�5�*�+��$�ϋ�1������"�SH�ɱL��z]do����X�;S�J4aHb?�T�B�~jIU0��'����n\Bb�gL�]D�]��hQ-J��җVs&�(��Lɋ�γ-��?�-���"�q����x���-#�o2e��^3���؆Ж�E>x�����~��`X�Tvڋ �1t��ϺRa@���,���Э�
	��Gl&��%ճ����D��ȿ=��c�ZTFi}=\>�{�A(�$��*P�K73�}�����r+��,��c�G��˒X&̒v�un�y������m(k���Q��鎟F�.�����g,{��,�\�z$���@*$�4�z�u�N��6%�I��0�j�Y1�(�.�U-��w�L�üAD�F��0t�'��B�#��&���Pō���n�έ�'aDb������

|�_�I ���D�!�;"-C�,�m�̟�{Q���(ʛi7���v���!��Գ���N���q�3�?��`�3�	e:�`��7`���&�B�^�kE�Z����d륒ˣY6������}��Fy�f��1����T5���Z�^��"`��`&G/#�4���K����(��+����L��-n-�x������Ra�1�ZB俈3u`!j�&B1oo��hD'����C���7��KH�H���+Ϊh��X�B'���j�U��5;P�ӕv���ل��W�0�U���q���kh��sZ�Q������
�R���e�"��˥2�.�4٣�����A~2S~Vs�|�sLQB��.0��GEg-?f�\M�?�{�W��<$���X�V���l� ?�(����
�wa�&q�-PR�h!��[ ���FΜ�P]_��'.X֙��){� &�B�
��3�dy@��5�����s}!q�&��A-�R\5���7�5�g��f�M��C{�f�_�K���o�х uD����q�Ԝ=�&�Q����y���:�ڮɳe����'9y�)+h�O��7����?p��Y�����ɓ���/`S�}�,Jg�Wg�,�zۚ��y'��ޖY˘��,�)I#��,;�ML �����R�q�$�������Hhx�?6��!����dx;�u�u��ӭ�_3��.���<��fыH?����|���V2uC+B�3�aIڧ>ׇF�m�L����q�kF�7&��B'7RE�������(��w0sX����w���Z@)Rn��g0s=����%�j�\�
`��!l5.(��wΦv��55���jLj*��n�`�/0R��b���I7F�{5���Ȁhܞ�2��~�$����ǘ���iS����e�����^�x~!d���@�*܌�]�*9���	��=D����2�3	��_�SN
f����>R(H����r�u	�|��+$+zu�'N������}�o\ǆY�u����sT�̣m��iఇ��̼%N� w���`�*��ch�f���i;��I0�N�It��?`~YvV���%\SV�՚"�f3$��^����rEr@��O�qP"��3��8-�����Y�e(U<���O�h
�Գ���̒@L��#G��[��x���H��]��j�c��ug/��ݰ�����)�����|���Ք��!>Qz��`��V�T0�;c� @�Y~q�q6�  y����8��t���(�8O�0zJ� J����e�5ĭQ�o��JI��������m^ ����3���,�����L0`c!�<\!8��Ւ�)k�.��s��!�-�\���98����!�r�k*����L7k�/�󱥤��۸�ϒx��9��?A@�&CtR>�V����F�n�5]�0�L;[c�AW�l�o]�`;
�^�iv��Y���lRݒ�a�ȕ�]�V�G�yg}L{�S�>��cNI��E	����W��	�i���m�i�b@��p͋���[�8��9�{v��@ǞLp ��9tR��b�˔?[���2�ⶌ
�h4 �e!"�$�|w��ȉ�K�{4��'�̧��$��7_Ky�����v����������T��~�B@B}X�/0����Ԫ��a�Ai�	��G�3H��4�1��h�"�iJی@P��ni?���_$`�0�jq�0j[�H���L%ly��64hj�4��?�r'8k������ZC��>�-�@��׬Z����g��-Ϲb�!˱�V͐�Z���1F%;%�GXi��c�V!������� �ɽ�Ӿ��>��7�S��<)qW�^�0 ����d�8�!�g߳��9��HO[�T�É�3�����6�^E���j��EN���Ƿ�Ӂ��F��.����l������NHU�CowqC	�-&�n$�z��\�b_e�{79� H�x�
����ދ/���B�
�e����l)�i\����-�<���iaޚ4��I�rh����@d��w6t�ݶ� �Uw�W����n"��d���|:��v�D�l;�8���˓��ɳ��U�7�P9H�[���+�߯>��H�1{=��}�����!��9z�}K�n��f����)z����s�;��-��-y��<:��:��l�Aj�+c��7O1)��\��yIar����\B��:T#�5�`\�W#N'mqN�k�.��x<<�u\_�a�>���6�H�	�$���ՉW�Ǯ���q��X�fY�Q�Ⱚ(()! 驤�o��F��Ւ��X��H:�!;A4��j��۴q?F5l%9��#�tҶIq�I��?eA���|��&�vl�v�ˑ�#��n>����<%Tz��W<��A|���im��=�����m#�C��(�z�S_�0"'�r �`���v�8x�����N�_���\�<� v�4 ��
��a���e���)eSGxE>��hR�n���	��F�k9���l�K�s��$�vʳ�H��|ivP�qzK�B䥒�F�3Fv��.��Z?M�I"���e�7�1�z�;l��#�7��_�g�h���5
X�Q'�,�-pQ@ ��}Z<��޳hӉX��j�qz-�:q6P�i�ӵe��T�sߵ��u�����F��w�c���������I��L��-�'�X�	�9�Q��)v��p_T����$���"�3T��}�gE<[�_Y����bkT�]_T�I�E�2���KJ3�ɒ����T��)����]��dG�	�N
^�սrP��7��5X|x���7�E_�����a�#ᠨ2dD��}�av���k���>'ފu�esr���8L�2�r�m��EY�0Z�J~�#����t\�>.�h
��:��..{��eΓ�n�S��Ko1?���r��߾��?!-�U(�7{�+��+d��`iP9<�$i����X�L�W�|1������u;�Iؗx�5teXwOc�\�#|�n�Dz��RY��Mg���7R;K�Kt�"y�j��v�P�C�=�;���l@FTkBg5���l���HASjQ��t�)���Q�9�O?1�iPV��iڝm-�8(b���d�H;g�t'�P-�7��	^���R�cv�C�s�&�?�������䋎�8�[og��C��v@���c����� �m�[*�Z`؋��$�H��t�����*x8��8�枏�0��%N��1���&r5ŧ<��҈ޅ'=E�p+�4���4S���|�@N�����T5���U�1?i�Ѿ.�_i�Q�[���!�����}�%y�	��r^�h䨿b�G��W&�	B]w�k����$g�(4J�p�j�
x�G��Q���m��c���>�X��
r�b7��3�����8�����%?z�JMI���׫�,�rmpv��U�O �;�+��}K����7
7�z�!C,w:�=��{u�t�6L�F��4v��f��l;K˶٫h:���#h9g9¾�_.�Ƞ�FKf-ŋC�� �;�n�����f��#Ė߆�J���"�/�����,�,e%"1^��W\�)��]����;E��ħ|�{V�l!�==m`�\��}=����͐#�r��<&i|� �Wm�X��o�gϽs}���k�yy@�߀O��t�/_'z����ӈ�~*��ۢ!<�5��ƷG��7������	�,͈?N�����f0��;:�RKe=A ]W�I�Ж׏Q�Y���qY��t�^������_z`���{�IH*�ގY�D�s�%��!���s�h����!��x \�Wl2��!�/Xܠyc@KwM�i0�߯�?�����Q�����]&�t
��`U�j4WX(��QҽA�џ�C�w��;�FAETl1O��U�1~�H_�cA���w� k���:���0���N!�Ze弨8d����/*4	M���x٤����)���)��]r��!�p�Э�$I�c����O1�Ӝ��#(��V��"� ��j�L���^\W?���'c����iz��e��G5yX��#���<�K`�t:�pP�bd��ݢ�@�t�����U�G�L-)j\�v)�2&#�f(�H��#��XD����C��Yy��Qp�Y`U^� ���m��<�q^lՕZ�<?���G8�=�vxމ��A�JyO�U�=�����p?Ϊx&�r��J%�}�����&��>��連��޻�鶞W�n�CU���=��I*;F��á0ұ��P+*���@�6�k#u������
E5{Dᥬ�I�� ��Y��Ll�#$�q������ZA��ݓ�r<��Fa8�J+1~�ѝ��#	,��st{��g��+mˎ�d��W��x�k1n�%�T�SOL���%)�	���s�t�VO)�;q�=�PP.y(ft�p��.�b���c6^��N_����`n���A��H_�che�`%Ɋ��X��������5v�G�(��oH��`�-��C<��Z�I��up澷R�[5��ca_n��|\ڼisɻ��}�=���C��	:.Ft����~�aώ���M4ڬ*�Q3���Ɨ�
Q�̪���Z�HJ�8���Jr#��'1�&|�.qC1����0&�,VωH��qۮ��SnP���`��7��w������U͎*����@�SY�d�Uؖ���
 �O�Ѯ��� !��n8X�<%�ʦ`o�����o5,ڡ�Ē�m���e-v��E�����jBN;c���C�n�7��Nҷ��OO��.�d}>��� ݆R�kb;?��,ގ/V��E���1�F��tsG��
=��bԏoޖ�<��dc����y@o�x*�;)�5���i?���ݢ�����m��#�-���Y��䴣s6Z:�G[�<�[�4�2�k�nq`���9���@"ǅY	{ٍ�?�<�O�O������4o��7.P�Q�&��s��k�b`P"��u���rz���rH��D*�`x�C�iO����򵇏�