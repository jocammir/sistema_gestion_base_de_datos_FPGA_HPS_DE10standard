��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T幫$��7��`��$��l��܌���������(y�U�+� �i��$�,ON+�������V[Tf�rj)�5��W����C)_k���>�PlG9
���EQ�Qh�v���@���p_�|��rkBK�yѵ��1%�V��dm��(:��-}�%��s�Dt�BK�x�^_as\�Ђ�E5�FW���I>4�q��GG���6�ۄ�	�9�����92���*C�6���T�0��X,��o����dsw�{�r���4�:�����ѣ���憉��L\��.1��O+�9k���vFg:m�hn+���q�S���,��W�#z�ӻ���!2l�ڧ*m���ZĄ|5n�~��[��azG�EF@6��2�:��ބ`Y�Q��mɂ0�rG96�z�ȧ�_�/���tъ.
y�>�
	������Zj�8��O=���-�y[���Z�cZ��S���q�J�ef�y��
�������
KG �j�cM������®��h�����u����!6O6�gR��Aϕ�L58.�Hv��^O������~u[����V����u?��[��{o�Q��L�/�e]���L��H�eCzZ��]YE�����E��A��#b&˷j 8Hd�ٽ��	M0A�p=�9;��m������. D�gd�.X������ΝHe��w�(2����2��S�S�/:%{U?"��m�|q�G�5�{���� ��BF����m�����.)�{>�]��ݴ���.qg�-�ѱ�S����$�a ɼ'��2��/^V�V��e��1#��"]�av�c]�zFdd�
��4W2��9��&J��I��%V�g�h5�F�b"4,���u<��'��_�����%��
v�Gx�t��,�A�S�!�Z��q�D1cj U�c��N�:�<��}�
��z{�ݞ���׎��;�E�3B�C��S\91_�5ڱ+;�Ii���vhA�v~��M���C*�f��ƺ��1����Ȕ,l�=��(��	��	]��E����eW����Y�1R~9>3�?a~NF�On��e���,�v����!5��]fF�젚�0�gn����k�<��}�sHDҩ���݋�|'%��<�O�)U�(�\�9)d �m���M��ۚ�d'�vû��F�ć~�@��ݎ�Ns�_�iܠa\�S��,>����}�!�f�5>=�I�SĚ3�f��6��N��Ԧr�4����@s��cfo�4��jn� 3;�����g�	l������|(������J���3����)Nyii����_��%s��$����#9Vª*&�ѩ�r���aS� ��A�&�Ͱ��)�s�� P+2��.c�qc���)���"����l��͞Ε�EE"�ƒ&R���p���TBB��r_��MB} ��l"�L�.q!9�J�&��Cx�|ơ���y�P_B�~L��G���(�;K���v �3���.�8�D�1S��I��ͻ�K��ךR�pnп�cv�淦��R�`��}���
�fܐ:�.
�?��*^���Л,�N�!
��<s��wە������B�ʜ�l��;�Џ�,�M�&^��o����6�\L,ϘB����Uax�JY��0|D�,���&�1���c�ѫ�O��b �i��H��X/&����首���?�'��I����i}Z��_ٜ�9CX�y:���/�x��y�#!_��c�Q�[�Tܡ��j�.9ZW)q^h9���g�x�%_��
_DJ�X���Jf'�V���g�`-��<!	�Z�.49�e8܋�3<��s6G����d?b+ݜ�hs5>�������#;q�����>�wQiĂMQ���l5�`��K�q�v�6(������t�����C�o^35���U��h�x	8_xi���$�L��jA��J�
d����7pFH�l��%�G�T�><I9^���ۧ�L�ϕ�ʀ���t�_��[1m�a,(��|�%q�[(��R��0I��g��k2��i����$�m�zg>#��B&���yS���s���/��Q�4]�S��ij�90�iA�<�O�Ô*��Ϡ�+jL��_������a�3y�@��pT�B�5(E[�������/'���t5MmmX�@J1�;q#L�q�*�{I��ҋb�g�S�,u�7�<�5)��3���Ş�h&�H�T>��� w���[���F?nh~~���V�@
��	�#�ٸ�`�rԄ���� 4whAlg�J�α������X�I��H�,�����ۤ2(S�w|J]�7�ٟ�?ո!�n�I��.r���1, ĀWƆM@���+��V��c�aZ�D�)�d�nz{��]I�5^�ay���8 
��Z�<�a4���RJ�ؗ.w,ɀ���5%x�:�8�|h�*�{��z5,�5l:G�:G��iv���<��	����~~,~T�ol��\�����&����o={i6���w�tV�爗����H�)�f���Q�jaIڟٷU��Y^W�d_��7�Y}%�1�ix��q$vl�F���w��qޥ�&QYZ¡����<OT��&����V,�o�MY��(~�Ki�4&��޲��Z^�],��Cm�a�c�	&k 87�����C{�f���Ց���e~Fh;�DK����-��:z��g�r"�˗F���5��.���<�X��CZf��ۜ.�<����%�t�߆L�����b/������`v"n�Y�iq��:�kA�v���ҕ�Ʉ��ѡ㪔�u��`�;=�HUte�\�-������XO���VE��aJC��&o#t�1��a[q���͛��S���?�Uq�n��,�y��j�??4\��Ni��O�hy����Mv�9F^I�8��H��� ~�w �j7te�8��f�I���n��P�Fƫ�� �� �5	��o�-'9e��m�c�+Y��&��DS$��.���8!%CU�U]z �Wv,	�J�H*��C)�fr'G��A��F[$���;ZgcU���1������㮈A����*�q�'
@XΪ�c�0��H�I��E�DׄRA��t+�[�r� ]X�x��S߉�U�v�$t�������0%���T�uS\\�4ar��'�#�{b#�傯~�����r :�M�}a����g�1p�(B=��%:|"�x���Ûn��W���J���@�g=1S�4��n��?�I��N-	M�zg8����9��l�vz׋�	�f^^c3��d��n�	;Ͷ�2VrN����A�@��r�sҳ�� ���-����Gq��yV��P��	�����.�j>ڛ�&�Ns��y��x�nX�y ���?�U}�RPY��ɣ^��7���2s�Jx�Ň���O�V�)yX�4���Jò�[�&��3�t\A[���+�I)�Lh�e�lIi�ٟz]��ŧ��!����4�쬮r-�Fʟ���umG�K�N�m�q���ڀ�w4n�*>j�;%j��B`F�����?uM�r�T�`J	9#�0�!r��	���� w�盋�|���e�?j�MX�X���cZ�@3�ӽ8�
�_�e8$By��{��؎���?K�\�{�B藀h;�$=�K�E�N�ml�x/�y����ѭ;bq�E&�2��ɹ����ۊ�0r���j_6��/�֟�ݍ Ԛ�)Y�)��HH�4i��pm!~\����9
?hM�T�Ǚ����A�ζ����R�J�H���sg�N�ͅ
�D7[4�W�)2Wm���-��p0〚RI�z��Sg;lv�7��q�`Z�n?є�5A��0�9�b�$0�'X�:+�Y+��W@IO���M��s�0@|#�/��Fw4䧌ݧ&�f���M��p+��d�모$s'+������4J۽���=��m�R����Ԑ�T�4l) ��zN%,O�ͫ�k�kEb�+���p���}g��?k�Ue�KrР\9I�%Nc����-l��\�V�����[�8���5�.��"��Q����<z��W�"/��X�ّ�f�9͂�#zsԿ���8�o��|mR��vX1��ȴ�p˹���w�G���1iM��S�zW��9�����#t�t�QI ��6���!T�B�$�EcfF�f�n����VS�Y�ʤ�Քv֢���Q�WQ�A�uA$'x�҉ܴ��,��FW�]s֦(l�E�� -�}K�]���E�2�K ��J�,}^��.�Xux�*)q�Eߑu����ky�/\q�C[uQ�pn/2(h���#��D��fm���0��<��L�*�w7M.��T\���e���w�Q����jTh���Yw]CҨ4�	Zx�%�ut�R�q;n� $���I��|�:}��E4B�k0g������p���I�.6B����6�{���#���˵�e���'��	�y"�La2S9��0��">�[-K�l��"i��o�(�0H�i���+6:�l@�P��.�@��uh|��v��Wx�ai8�eYmi�z�R�?�7`h�� ��G�V`�O�o��6�Ǟb-�Zn{�i� N�#���w�d�]ƣ�1��/ �1>�K�u
1�ao���l�d�'�ep�X.�\]	#�� ��,����Zc�:�>��{yJ���%�AE�ju�'e���CEV��[����$UfqN� '����Y��]u�mU��i�Zpְ��T��7�X���:�x�x�0]���4�Ue�
r�z��ɨ�="J��aeS���kSҟj9�(����~�ԁ��Z3y�4tI��ރ��_�Mp�f���c��0n���&�D�俫��?� ����˹����f��(�E��V"VS�)?&�He>��'��L�ai�^�1����k�^Tk&�D�X�|z3�Y�6�����P�O��u{��hK���L���bM^TQT7�ª� P����4.�����,��Z�����T��^�}0���7����}�'ө�$��i�34�w/��1�v���9�+d�igC��5���ޔl�~�}�q�<3�j�d�]A.�+c� �����/e����SXU�H�(;�m�42Nx�
߯+�t���Б�[CD_�n�+0�D��QҌX,V�Y�	pze�r.���(�8΃qXw~e`��h;�c��4nF�g]�v؂K��k�VS[�?0�øV�6~�A�H�r�;�A�O����RVk�a+�)t"����!z��F"�ؙ$nI!��k/c�%e]�qteC;�(� N-"�	s	���ZQ��EZ�v��*Z�Y��jD�0��=M�Q��v��TD?��d��͇_��L�oC�6�n��o2��<�}���\� )��S��I�h_<����u8�q�p��x�%����غ�2������"A��:��|f^C8�=]t�`�.eB���F��^b+/IaB�6gE��`Lt�ޔ�1�����<�9û�;h���[kA��+��ްܰѢ�H;��5�������^��=�����&���C�O3�Fa�7��_D'-�4)K�ŵY�u�'D4n(#E�?o*v��s�͑�Ne(���s�ѳ=��
��҃��̗4�84������`�m|�� z4�b=q^����O@�D��a,z�Dz����g���KJ=�+a���3ϴ�j�0 <�jŅ&Kj� ���	�E+$�����o�>.7��Na��@p5Ex�1lǷ	Xɶ'~c6[e{���^�HS�%�h�(���2<I�um���%��҂�X��EmR�D��	ґ�{��y�I�nS���-�57���PK&.O���:��%�������j�3Xm0�L�
(7��@BC���I��&[�,[�����Io�+�B�ؘ�nwR�x�\��/7��$�t8�F�	�r;}׵v�0�#9�I��_�Jb�t�6�is��l��ۯp��YKI�H|Usf^�I"Q��L9ؼȂ���G���ߑ�pO�zz�.�3�VS���)��O��ӡb����P1�괳��'�x2��7���]�������J�EK�(�.5Z���9ev�h��eB�ntI����{�O�i�d��l��q"啟��3 �oh��Ч��W_a�-2���f�� EN�焏���)���`�m)ל�M�>-��K��~� H�ۑr�b]WiwM���ad�e���tw���������=vlfD%%v;X���>�+Es�t�|�uZg<�DQƩ���m�"JEd�c�Zf'�HH�3M<r�)zO�"c&
;@3! m�@�弗.�
���4��	KBC9u�r�؊9?�C��̗.���*��.����p:�9)�F�k��H�����lf
2v�?��ه]��4������������>\R1�K�A�q�A�O��RVis�0�\w?	�Z͆�K�U���R|t!��ܒ�'̥���e_Ad��z�Uv��m�> Y�";b�.{,q���H�ۙ瘧�c>d9��kkZ�Ḓ�	���}�3�O����9%�Y�_Q����n�
�I������������R������BRq����K�3Pᙩ�3� �A�=����j/��}H�� ���\8��ؗ��{�
��,�i8](W�K�y@з�q�f0��j�(�i,����==�X�멺DX\�ۚN��j� B�tǊ�'՛	��Z�L>�3�T���1p�J�e3�_���ݴӱ�}M������ƪ��5w� �]_j���|z���[H��$G��f�˦�3�t	�f���U�n�M$]�n�E��� ��Ǝ"�����]ZdT�	23���5��_�r�j�kdW�	fAL�Km��C1�"\C��> "�e��暪�+QqkmMNm4v�K�\����Q|MaTeN����ӎ�(����ʢ6�~��A��~y�	J��Ԗ�uy\���R�[ �E��X���yHt�0�A�� �\L�f�S��M�7��u�==�d��w4y�-���M�0ɋ���Z$1{;�t'�d�k�k��G��ax��A��:�� �3���+8b�����?��!$�>�6�B�Gy0�������w?��w�S����+G_B=�S�,e =K���c9޲�Vmq�G��Fq�(��e�%os�	:��A��"�^fy�A�PX��Њ3�J�J�eW�f}rWx4�jE;�5m)��x�kr���Y8g�Z#C�Œƽ��\�6c��N]-f�/�i����O�NA ��VYFe�-P'yzLڑ���vD�����C8��3��� K,�>��N�"�Tϖ�B޵������ګ�0�Y��d������e)�;����_j��I�
3 ��R⫼y~��Sfq�������w�p���W��NZ��=�������('^Cs�S2��8L�٣�p�Qh��-�Or�I[�#�j�:���Q}[��!����s(yu�cL|�<��_�<'H���	�6���b��CY Ko�e��a�cHa���B��L�,۾���J�~1�_��j��m�<���3<'�����ph���I��u�0����� y���s�N����.���4}su�ρX�a%s�(3����?�~Ia�p���%';=���#��B��-��(kճ	����1ԫm��K�y�,��È]/4*��9�u��?���>��w�f¤�y&vJ~j" �@�\sfD'́�#�;c-�Ūq�pS�X��u��uJ�J�n����"�ajR�¹ʵ�f�U������Ԓ6����W�7�v7v�,J2��n�Ȋ>2ӹ�?VkG��/?������ln���G_]}B�\ld�w�^�5j���RWf�-�^�ƞ�[U��j�'��C���W����.M?�F�y	h:�^�:��*�'����+�	t~������$�ɗ8��@b�c������Y=�����E�T26�"{�e��Uf#{�~����yʔ��/����92p'@t��i�t}���Z)e�&ц�"f��Wv����^ͮ會�k�&�]���tvs=�w����?s}��`g��|C�\g?n�r���_N_�JLle�wn��QZ��m (��&͍�뿶�5�>�:�JD74� �8LMr�C&�"�5��Ԥ�1��q�j�!O��'�-+�q����ikC���0�A�Za�A���lnV�{��+k�M�+B�t���{hD=9C�f�܊8��ܲ����y*et���ZE2a�Ԯ���76�HhO�.��eG��[%����q�C���TD�3��Ӫ�o�+i������v�:�1���F��O�A�(�҅`��Y��+��m5��N��[�-a�42���(����Q>M��'�ޢ�{�'���gU-+/K��y��0��C)\�o]R�f���C}GPC��7�)PKV��BɚE�@R� �j$�]7rF�b-*DP���|X:f��{�f���R�]al�}1�f�i[��y29lCa��n���VںQDOB>��Y\)%�	��|�����C[9���+���E����GjB`!����o
�������.F 1Q?��!X�k'q�Xrv�Zf���d�b�XmrL�AZ������GO�<�V�&%���,�QB�X�<S"e��gT�9**:h)i�s~Dٍp�޿Ö�����I�?ߵVTd�y��/,��&��a��@��x�� �n�df�LG�r���0h�,����Wǌé,�s�Jvs2lo<`t��I��U�ҤɃ��OZ�f�W&�K�D��Sŝx\���,�L���J��3c�,;A	Z"8ڄ�1�����՛�&>6�!6�_k�O]ϑ�ǡ����gb��|�8"1�|�L>&�>i�S��(�]1f;d=�Ѿ�!�h�RzV�s���	1�L����Al�U�ZL��	�Ĥ̑�N��|��P��nJ��d*�����v���
skm�W���p�Xr�hq|M��Gw��c�k�,R�CJ�f�?]F�u\j*̟�o���N% 0��i�|~�K��v�jY�6]�1e�%���xgʊ�uq��w;�ԕ�;Մ�/��s�}����M���X�H�_AH D�?l)������"��rסWd�&vK:�`m-7��P��'D�Ձ&�>>w�nڬ�����ְ�⨩i���({v���
�^�-�͹�j�呼��f���<�NI����j�ٴw��h�Wo�̀�٬rt�����$�毠j}tqͶ{�@��rc�Vn�l���pט���|D.�oQ9y����=e#��F�����x����=�!��A�g����>������.���Hh�'緖���D�˝M��b[��O�_+_6�z&Y��Ⱦ�wc�����v�oý��V�W�L+��~bK�:��@A�8Q���vH�	���������^��C4ف�Fo>2�B�]`��D��1g��ԷCj�
`#�K���:��%��o~�̓��kD6r��P��0�N,���)��
��&'����1�(��1���e���߲e�^1Q
�P.���
�����Fҫ҈�^�-��]�`��C�}�o�/�7**@\�xTrttZ��-�Z)~�ԕ��M<�9�xX�����3Y�r�;G��14���S
D�h���Z�Χ���)I��l��<�18���DH̣�G��Gf� ����Z�w�n|� Kt�����b��j`�������ɮ�^6;J��� ��R+|�OU���~bm�n�N%����~e���"��Nި�!�m����S��B��'
�<fk�u�kUK�a�&-f8����H�^A�ֿ{=V�fi>���B��t��ԉ�.qa��?/�X�1L���L����Zמ!��Z2ZWRF�`�޺�"3E]��b��:Ɲ�I�8[�P��H��"L��G+n�D%,����^�U?XK����ř}Q4���
�$�̣l��dA�n��9�N�I^z�{�7���v?��5��|�S��cxxd &<G)>�* �)��=xwιY�v�=o�R[h|h���j,W(m�7�4��`��(��怅:��D�X�N�YX'+��Y���;�Av3�7��EK��by\*�_=�t�	w�ъFm��|z���� s�tk�9̊���G��/� �8ł��]qǏ�p�1qx��9��.V�,�����H������������P��.A@*������?�2� ��$7�y9���|������M�kw����I��[�V����^��`����qkF0px���d�AZcu҃I�����ו��I���jMl*�,�SEr��ӎ���+~���L���U�XVЇ��f0f#s�EE�~C���������g i6>C-$�� ÅhV���L �'N��i�Q���a�T$mK�f�:�4{�ՠ6�xm��|t^����%rDY���Fd �66}{�ې?1�wgd����H&A�'߿��S)���e!Q�3X�?9<��O|������\[�\*L�C��J�_��p�S]�/�Q����æ\ _0s��GNHM$�� �>�r��3�����~ч	�~TWև&�}st�/-}�[��)���o��`������6�x���^=�|}v���G�("pcA6>wpc!�e����L�g���#30
%�]�O��1$DŀW`���9���V:s�L���*7,蹔��b��^ �߲h�����Ar�����B�`�F���|o2@e�xQ۝{��sx:v^�0�c�w���N.�`�QO-����uy��ڤ
���*iE�S�0-��^H0�Gb|��ca��B�m�m��W��s����]�a$��T��}�A'%x{՛�5Q<o�!�L�;������I�{�2)��J�:(�R�b"1k^c$d���5٧����o�Q�����/rB�f��@hJ�J�����XC�ug(p!(���{�h�ϲ�U�F�OZQ��Km@wR.���Z�q�ʂ��:���?���Ҽ�e^�3ī40�´�L<x���EK˭�ּ�:�3Ș�S`C���� ����[-������ڽq<��mcfM��Q��UhY�\Yy�@�?��{��K���
�y4;}��ȑj:�%��	�ƽҼ����BD�f2�'O�0�����+�:j���^�� ��f�������(atǡ��>�����ܘ^�˝���P�R?�^6��;9���}����uGZ5-.7n�Ss�[Oya#�6�a�E��q��IŞk%21�=d��0�C\����0HL��$S���X�[Jȏ��������ʠ�&t
���mF��X	A����Y�Pe�ye��p���	�����_7#�ˁn/S4qm����:�ͬ`_$9�3�m9��1�9�览�BwY<��V.G����`W��r�2Y��?K���64翸1���;��'�:�G5�b$Eib.#�@�A��$Z�U]���,���G]�r,��[��Ǵkh�d%龚2I+����:�si�����-�QɊ�vsZN�j�Q�>��"�Mw.2���Y<�]�w�tٞ�jf�:M!��!�Oj�`�ܙ�I!h�\��Ͽ��x��x��I�	�bk�ǐ�b�R��1�Fe'f�]$y7\6e���[��$���t;��@�J%z�&P19~ '�mX,`e8ޥ^'m}?"�	��Ͷ}4j���u�����&4�t<��O8���nN3xk�[��;Km��$��'�:�U� x����Am� ގ*]iJ���/yx@��cB1ޕL����	;U���Ӫ�Dg �uZ�Nn���$�΍mU^U,LЌ%�l�n;m��]蝒ڮ�탚w�?b���G�!T�w�F��
�����мb�2�)t�C�x�ŶdW<�:G,��wH@��=�f�K��s7(���L�������(!UV.ș��S����*Tw�/����
�2����_�
�ӿrn��=@><u:�oV]*�}��n[������C��祇	޺z)z;�|��8�7[G��e鷔2�Cn�9�|KdΈ�Rn�o�C']�.:K�ᗊ�
�0$���'��pQ>D���đc���/<C"��6q-8�T��`˓�F�)�Ɛh�|Bڳ�m��}���BWC\�ު�%�&�Q�t^���������l��T���ik�_	G�g�� ��4��`��kM/���KO|	12�caL�o#�7f�	�9Y�U慨�i���{Jഐ-~�����C���n���9�xr�~�[�@[��^Dwz�s�� 3���*�h�	y�G�v%���@��@��̰�J�kR��]��m��Ʌ� u(�i65�V#'�%�ڪ;Ȭv�۷qD��#2�Vp'���+����*��Ć��gjQ]6
N����~hUЉ��Nٍ�B'|{��g��*��3g�7gG��_w��:.K�':�O�i��>����a�釬�WYr� "� �y�Y,��hJ�Нב�h~եs���Z�	�Xi��|qx�lΓ�r��De.��M��Wط ���a&�p����iKl��������"�qlH�X�d�Om#^1��Qe��h.����ڭ��M��]E��n5Pjb>�`]F�ś�9a��t%U�6 !�9��RLG3!�.w�� C:�[���݇	��\��v�ix:_�ؒ	��,ҡ��v1�欸}�\����!��$Z�\M��jP�}3�n8��ЖյC�%���Bn�68ˆW���E�&}K�������,�iU�D����R?EWꍳ�3�/�G�Q�Qt�7���a��]�j��W�a+�$D";�n��<W�NTqӔf)�>�7x4��]o�������ZRNl��Y�s��v�F_�E��?Tf�Ӌ	�X�4q�6��վ7u�Wf����U��.�d�_���"�C��|�AM�2�6~F+(g�eڄC�jݬw7�9�RO���f�3�xg��䶤zk�-}Kƃm��4�����:�=|�Յ�{cs�đ��B(��;�����T�Ȉd~�Ltۊ��V���l�Jb��`kƕb��#)�
\Dn#��.~�Q'~ Ʉ>���FV�.��&Ɖ�p�ɍ��̴gQL����cH��)�|�2T��<�	���U�𺶶	��k�[���w^]'�BA�7�q��.3JB�C3?���l�&X$�5��AZ�P��w�n#�Px�6�:�c��	�qK���{�[�ݞZ��i*��J<��]�]zb&�-	��S~H'����X��(��{Y��WC�h�_0�|��&�y.���R�ؓ�
F��'�<�-̦`�������=�$<:-	#:Z��4�@�����i��a��������������"�Ry~�4��p�*bJ����iڄ��Ԏf� �����ɸ����uz&A�ھ�q����w2J��B�v�C�gl� �à�A&�0���o�4v���7�V��
���FA���&H��c����QnB%�1���W#/�!��köyZ����4��-��^;<� ��|�|/�R�B,��E�	N4���[��ަ�g
�\@,��62B��%����������X�Kb���Q\��8o��'�h��YGv$��3x�l�J�IQ�ۡ{���!��P8Z���#_�ѢC�^�'tg�b���������NQ�\��7���.��mb�PF���}�/'��t@\o(����I@ �o����+�f�k�O]bֻJld��E�
�U8�(�c[�p�F��2��1��6r��H69��UP�KniusI�C<�&�#�|"#���$l�K,F�,Cz�	���Z�x/�e��0�
��Y�p����*܄��t{|�aB�Ј�'�w�*����Eʁ��DfK���h����O�h��(�Ɉ�"gi�-�e�|�?`���#�#��(��=�u��~X"���n��l�gn%�m��=G��o
RX�c���%�^<`�ϴ��5�A���7��%«�	�G#�S�g�+����?�![�>�'-�,"ׯ�bB;!k0����:���E詤�F�wЗv�My�XT���^}��5&x���r7�<�p=����u�8�RX��D��Y�uC��D�f�t�%��٬�5���:2�t����	ރ<�p��҇|�{<*��
�/��Z�.�9.կ��lG=s��R/�}"�o�U+aŜ�>A=�{O��g�;�\����l��M�.VOAG����j"��7���Bd�E�ߣm�qٝ�B�QwL@!;�鎱
���1o��������i
��Idjl��]mz�6o��m=)����dI6����c���CP��Y3����0��?"���娣u'��i߂&sjF'%��فO��Θ��Bz�&�7�4m�-���~��%Ӑ�c~Y�o� Eג����q�ʕ����_=�:[����|G�������|⠠_�<O��0��9�c�u���ͅ1#w5e\���-e���io�p1�(�zL��l��Yl�eµ�=�<���K�f%?ʍZT?#��֨����6���bO1x*�S_wM�tb]�/Ѫ_�o�R8�ǹ�/�/��NGCI���ɣ�%s�O	�����(DH���ښEN_�W���ZW�Y`E���z� ~��cd��VZl95�c�?(�6@S
}��f�����~��%f+�^�O����z.$�o9�Dl�3�ʉ�p:���9o��k[��%}�3�$����n�1��"�.\��D���)�A�h>�n!���� w���z'���"�&�,���[��f��TdݷM�-�[�Gҧ��=��چ�+�;2֬������쫱]յ`<��>Lr�U��n�Ƀ_c�bΜ�;)�k��B�Bi�:�)���Wޙk�Ӝ��*��2SA��+
�0$�)d�&-���r��!.-s��[�G�:��Z��/h Qnh����r]���A��ذ�F$$Rȳ���a����>T^�?-(�i���>ݟ.�r��p�cc32V�b��P����[ T��iT4́VpE���x��]3�L�vIb�e9GA�/��^�G�������b�Q�E�^e)ۻ�l'h�a�sج�?(f��yi��0-)��Sn�`8����:�y��g���m�M�B�Q+�qpO���ϱ��ſ�"�Ӽ��kc��b�1�.<5��"��# �aa���Ƞ�3������� :L�fɛ�Z�m��COhutpF�w���]:^*esg�Jfy�$b*8x���݀\��Q/{R��Z�PfE��l���֬F�'۟�I�KЊ��Р8@l �X����G/�*�9���(H�����]*N%�6��I�g�G��/P,��S#*`-�҅�5��v�?�UQ�r]� �[�1�'0[�V�8f`��'.TX9RBJ_��
�pi0�p��hk!���b2��x�M}
r�X��7�	y��MS���+1 �x�v����|@c�� ��[��G�4=�^���\�s�tBV�ĞR��睚�;�jQ}ꖘ4���Nzh2wFM�Ř�"+��w�j����['.����ĦwC�B�W�Pua�059X��=��W��M��6/�V_a�x�h�kt��)g`�5I�,k�����wB��T�o�d���ղ�ƣ-B?�}��9��88��;)���;��j��ij^k7&;��>G��l�9���T�Pμ�ac�փMo�9��� ���<�����;��dջ��]I�z�����,�`�Z=m�BӮ�����&�ή$��b��w8���	γ�T�ه�7&�G�M)O
��i�d�I�B��|Lu�hh��C��?�٦ςn�Ͷ��b	[�Ѣ[>1�4��̑؋�����*�X�m��m�6v��;�z��~)�mA��\�Ɇ�����)�W[���\=)����XxHƀ�KRM��c��P�����j�`�r\��\�N_i���ήx�m�3���&����{�G �ۯ�-�d4[�`���ǿ��QgK�2K�'��ӑ��J�$5�qm@-�۔�~���g�Ω��fI�(D�sF=.X��UnP_�˸��k?�	p�� �7�-B1~,&������3�_>�gJ���)�C@�n���F{ԵBс��z'��ڭ�����1%x
1f�9���c0Y��p���fĵ��k�|iw [F?P~|;�6�"�l��w=3;��O�� 5?=7�^�]�U��(̨z���,1����H����ơyzJ� k�R���al�Bm�3�*@f�>��\뤺���S��J���*
����*���]ם2�HðU�-�ĴK��V�I�.(����+�	 ��IǶ'%��*j+s�t���%����rEt�Hץ ����?Q�Q�J|r��锷�sTCu�KXAh4��N�5�V#C�k�ö�y��7Dj��>��!�TΫ�tٴ!Ԡ��T �+����]��ժ;�>ƾi~_D��)��ʸ�Ր8�8�x�Uf�����J�8�o405��ԭ���GeA|�#���<�I��8bh ��E� #x�-���M�sA�6��{Z����MԽ�G���֥'f�f4�nHِ��|���f�OΫq�d+-
��Sr�ш@mPǛ^Ki�}�x~
�'�Jcr�V����$՝� ��l2�#Ӝ�b�E���MB�}�T���	���[C�#I�������T;G��A�7>���IǗ1�e�a �A���~b�uiX�C!ş�p��o��	�]�y�� <j�n���M<��v�/�euZ���� ��*�}�Ɉ��.��K�����h�����+I,D���-�L<.+��ŷ"K�g��#�t������	rǨ�Z�d�*!���7|���Ӹd�;SNWBE+�g�Ez�q�U?gAp��j����kV���RR��� M��K��9[�-��v�`��I]W�>'S<���y!�<��6�+�uØ��a�8g��Հ>��a�$D�>�A�Ay*���4�2;��L�����I��Eb&S�v��Q�`�:&gs�pBmBO���MP�x#N�{�`�b��oEua��
+uKx{�hL?}����)P[��dG�D��o�*����짖�N������R<U)�A'|S����դ�u'&���ߠ8ܣ"e�>�q��U6Z�����`�T(6_����Z�'�0<���
.%���}<��]!���k�C��w*�2�hsڠ+��Ż�����?��bF���e�h9Ȓ T�3� [�IK�{.$�/��j���Z�2M���d�C�\�X�[��OQ�.�����<�ł�!�s�Ĩ���w�|�
��,�E��wW�s�d�F��@�+_,ui̸����Zw'BeD	���F�b�����'6�E���!�>�H�c̟�"u%Q�o���q�p���o��ɔ��Ҥ�\�SM:R��-��K����B�o:Z����ʜbN�Vy1��Q$0�P���'b�m��=۴N�(���+i�n���V� -Y���L��7�bA�������"G�CkN*�I+�+H�RdY�_-���_�V�&���J�x-ƕp��l�y������Wޚ�2F&V��D_��1-/Wd���� ���?ɲ[%�-���q_@���d�ѵ�+��bP�ݘf�^eNgB0v&�$��F��&�K���%����%]�����?U���q����ģ�Yj(䬹P�\iI� q���J�v�������@���H����w�+/�t�Ui��S�������<� ����� E�f��wc|3�#�!н�^ ��6y�yk��v�6�]B�*�4��0��E�u�,09�ZC��G�h�j�e=����|�e�U����j��2���s�U�jth�`�,��납��41%�5b����^�s�k�NJ�����R;��$/�]Ȥ���� 6�z�8Jo��.����cc���ʹ6���o\f=��@`E��b�"�<a�y�>h=�	��>��ҡ�:�9_6��|�y*N�Ppe�$^��AL�e����٣R�۬�X���e*���D���V��$&2tW�~�Y��ʘ���pR�KXʴzǝ�$�jU���S��0[2V��[��K�3���F�k ~�T�a���ʩx���\����fK"�w��#��� ��<-4k�ow������}�3��Je��) }ql�UNz6O�j5�,�p���g�$JT�Q������? �XSi0J�d@%g��I�����1�7�|��fM���r^c��~�E�`��\
ާ�%��{���c|�0���N�r�^	���l��x��v����1�{
����M�#�0�k�'%2T��\�!��� ��k�M<_��X
��y�c'��m?>쿨�+n;a �X�z!��<p�G��N�O�/��w2��ґkSKJR	L��A�h�f���Mѱ�W���Z�w�J�I]��2(�|��̉����V������=���4L�+Ⱥ.������$y���5�م�c���bbp!��7�I(8tB����[���΀F���D��dP��Љ�C�z�o��x�'k�
�ǖ��k����Z
9:�z�o^v��Lz�Z�m�8�B���M�ڞ��Mv�4��
*�A�*T�hm��9?%z�Е�z�-��<K���l4\Z'�E̋�4ce7�(E:S¡�P���#R��3��ȅʖ+�����{���>�@I֊�ʗCy ܙ��-i�e�]����X�hY"C�27h:�PR��$�.���\vs�%�8�q�l�k��4�4�@a���I�A�^�� �a��U};���8 ����9��Ҡ�xmy��N�ki�;C*΢�0���x�h��p�V�ΐ�ka["Fm�H���9��`��"G� ��R3��.q�u�J�O>J@m�.Ήfd�VV���y̞�f�X9t����o����/�sv�<��2홽�gI���/���g3�B�b��R>8��pg�P�s��i�Ӓ�C$s�__H��Mt�n�G����E�NEy�h{���tpƍ�O0�9,�n�6�T�\E�B��U'��[�,�N�3�aa�m���?�q<�i`i�\^p��WW਻�͘�d�>��{�%ұ�x�Ɍ�=�'^�K��(����h��:����]� �2|A�u�:�H�������9�1�w�h$��-Eݎ3T�.s�4,����O��9�)6�j�!��tM��A�*���9V]��1���Ǿ?xdf5�3ع|޻n8�\�E>K}/ə�{?�͗�����	����$B���/��\mݚ5j��������0#�&�qH�ю������2G����~:]����9C�A����n�G��Y:��j�^�"B>05=�mE����͞B�r5���ϙ5�9E2��ZpZ�ѐjZ��3i�|V���"p������`3n���~i{�j5�*�1�'����v�1@�"�v��
�CN`�h˧$�� ����.yv#��ʔ���
M�o���M��1kZ�&������t�HلR��m9G*�nCk�m$�T��>���Q]��^�J`� ��q!�??,XU�0Wr��!�U��u5�p������aM~ �4�c�q}�|��V���v��Y�dr�׼X�����f�2�"}F�X�G�{VJ�ZӸZ��d-��;��:��ו{d��˄�-S�E�y^!\�&Z��܃��;�)å"02
��M�%�64P}{iL�%�@����*�,���7��D9�{�ȚLZɮ����t�b��s��_Y���˿�tS���9G�:t`} ��Ft�Usw��I���������Ǳ���{$��h�juHc0��yoGY2t��o̚c�d��e���OY��&+��@p�tJS�����;]���H*�wv�`:c�-�3�)UP� �'m�ݭ��[�������ra���A��2~ͭl�]��� ��������0���ژ�2|�����@6L���+�[\�cbe��I::�3�w&$���"ڿ@��D����.�|WF>��t}�GV�m�sN�  �6���a�E�!â8U�A�=���Á��tCf���n|��S�҃F ��w����pWG�P��&8��A6=�X� �5q�zV
>��ln줞�sj�ޖ�2���!�'{G�8��9qu(^�Y��t��^1{��4��
H��?�y�ٟ`���D'������`6JC+2ߥ���4�X��j�?���,�F��m�˵9�WE#��,Pf2R}/0�1�vPɉ��z�x�%-R��n�Zo�ڇ�_�������Vj(x냴4P�98�[b-{*�߀ٴ�9n�SCG��'[I��`�1�ؕaՉ��`X�&���^��	����ԐO<���"�bI����v�b炭����\m
�[I��xD/�p.���jwv�(�I�/�Gr{��X��d��d����S��0�f��㳲�tܛ�5�C{�rOS�[�ヒcdi-��n�6�.������0gP��^�6��'��븴BҰ�(NJ���칣�O����PH8��m�s��Z	"�2��'@:�2��� ��'�K
?�1v�Lo+U%�\_8�n���b2�A�],�k���A�����Vf�>:>{SԺ� <�����E�v��PF�}����-H���j��_���Ö(�y�z�WX��Mg��V@�-9��;}(3��������.fX�4��n�ԔLd;���+ !(�I�`�ר�=oٔ�ի��_�m�_�f�wx�����L�z��	=�q\���L���m{P@pl��=���G�]����Χ��S&���������8G~��*�.n���q�����y�EN5a\@b�CF2@�'�&�>w�=�X2f(�8��&���0�e�|�6�l׏(	�_ݕ�5�[>w�2Q��i���B'�z��� mQd�]�U,P�R)�p)nA\���(J�!A��ޯ�*��=�XX}<�0R�6��h���b���g�[�_)MQ+���x�]#d��_�u\�>�ہ;,Wm9�k?A�7�U�9���U^y�������)�@��ۃ�`4|a�G���=�Trv���
�_[R�)���%2�f"ޔ�B9��$Q��_� r+�E���Ԋ�gD��X��.�A�/�d�n�jJ��Փ�!7%5�k%.��,�C<[��WN�
���R�p
�p����_`O���m-���J;d�Ӆ�@C�����v�g�'=/r��,8�Kѝ��� �R!� [|QF"Ip�J����C[�z���PۍO/}ڇ���!T�F	�٩�"�H�Ga0����oܷ���Y�S�悸m[\�]���t6
����9I���聽��S���3#��=�N$1Q��0�+q����"�䁗��v�~8&Tn��#0�EC�/.���5:#�����c��[
���U�h�����I�W8}�;w8��1��e}-���0��=�t�൉/;U����"b�K���6�7�J&]-(=x4J-���UL[�@���
���e�����$gE[ Z��pC"=J�,KZ��DNU%@>�u�(�ͳ�Uz�Iל�`GB�v��J��Sj;�!���:��O� E��Amw�M��T.u}(����sú��6��4g�S[����ދ�"�����^W3	*��֛�<Ȑ_z�p=����|?N'�g|y,�����fa�/�����DX�q, �_��'����cĄ�n�^���f�#�w/����g�?����BYה�X��1B�dt�G����7��,/ ����d4;�����x�)R,�+�S��!̷v���|��	���Snl#ݖ{oIC�V�
}0?r�TB��G�PF����N�����v��`$�&�m�$�ѓ�:�֒���7%R���)�A&��/�a|�$�eD,mغA���@��`?�*�V�w�֠M��c�Q�[)����8s��N��f^�j��O��Z۫ 'c �v��yБ�%ӭ8;�+ԦP��T�AU�s�#vW�D7=7Xn¦��dR)�*��D_�m�Gb�"B�����7ɛ\/���ˎh�Ў�DFD������f�Y��P�6�B�ZF�u��\�ֿx7���m|�&���M�M�;�ㅖ�+��C��7��H����4vrb��f~ڀ�	~��m��wJ�XC�,m+�+:�Ȧ"�u-�[3W<.���q��[�.�1#�<��O?5������2���o3d��Z^���W<�HI��gd��,n�b�Jܱ�U�<�.4*7OE�M^��9�<o���>Y~���%�PWO�ē�A��f��D�\q���P�Q9"����ݦ6%xܫ�1���Q��dF��"���8�&�9.����Og���h*����0�k�ˣ��S����v��ڑ������Q<����C�
��%SC�<H���Z��r���8q"�����C��+;�D�{���U:��ޚ���WQ$�4�oξ�����c�(@l������&&�۟ �{am������w�/��C`1��{o��\�����t�/��M����<��?�NK������7p0���}��S
�au�P��e�['̐��$���E�vf�����@rPf3��LY�~�d�Fb	���v��249s۲@�JP���-xLP�O��o�[��7�u�y�.��zۼ�$��L;��i
VTArG��+P�~ԑD��=��L��-\$<��_��~;;�~���(�~4 08OB_�%�%�'\���ab,�)����W�F�/�B�ZF��U��W��o�|�a�����B�=��7�K#����Xf�3���9��Rɑ�M����Z�6dG#M͕^l"\fg/bqґ�QK�wٚ�7b��@W$lW������0�EUm�����[s2)#Ø�;�@�s-����,�$z�w,(��#mPC�`ìN=&MXܥ	���md��s�Kt�蹭Z���J�#�܃m�l��r�y�������;�O��z�t�i���oXS���t��o�	��L�F�W���X�����}�p�y�ˈ��H��U�]�v�܏f6T�t�k	͑�Hڢ�v������� 2-�ї�������m��2�틸�D�z�-��'d]�5=b�qS�ܘ0Jml�c����J��/�Foc�MU��/��f�3	K�ڣ���?S3�#���2)a�E\ ���+2�B����	�/�<��k�����X{���h��`�O�>ruǪX�w=�W7<�N��-KeF�w�B��s7]��!R�����v'U�Es�� O'��4����E�R�3��[��/(ˈw%B>�7�h���_���g�~�(�K��~��Q���0���f{��o��ƚM�w�hh@���+�G6�Dd�����
y%_#P�L�e��p���C�i<�[����G��-�K����ք>�V��ř��l�DfG���n���l{�.� Y��ğ����P;��(�i��lk�J4�_0�p���1��,(:�&���j�li�g��eN�rmp�u����)r5y+��I�p�SL�Օ�L	,́��'��5a��V�K]YV\�ʹ�~f�,�ae^(�<K�.[�~}���������ঠY)׶�]-
TT9��<U5L��_�8b7tS�Iip�Tr'��ՠD]�h�R�R �,(�w�˱J�-	h��G�:z��v�<��Y�{�F.K�QBH��V�o_ٜǯ<&) �u���<C�{q�u.�0]�.�-��q ��6��2N8��ի�ϝ��/k�T��H�MtB�Ku����#}�뛅��(vp��J�tK@n����N��xO�2���\U�q�0��s��|���̈́g���@M�M�ʔ� �E�s���_���m�v-^�����l��o�<w�m
#th�~���@0�%�?[&��"���i��-�^kd�X��=~��9/�����Wӫ��D.	�g�s�t���b�%܄71pѢ�f���W���P[$8�"�T�
�n�����XE1c�g)ؚĖ�JĴ9�B�y�;g���ж0ż����\��Gh+|+��U�L�e�H�5���s�+�Cڹ��ʁȠ�d��67���� ������n�9l�0�1�����~��p���3Ȭ�\�}��t#�6��@��ՃܠGn� nI���s���ϧO[U�h������6n}~��"+H�@W�2KB	��Zҿ-�0�MBg��p�7�3D�*C���6��O+��֫�&G�t��ٲ��4i=E�q����?(�� n�q�ta������Ń�d�p���nN�/�^ �O�C\@���Y��KIa�����	&v�J[t��@5�)�^��!F�Aς sE}�\�����]C��#��}�!�]NKWY�Ʋ��O�g�g`9}�oU�����K�Mf�H�3%�uF�W&*T�N���R�hK{���+$Tqÿ�ܶ�­�ZrW'2��8Sg��މ9�xa����ran����hR;���#�������Հ{ثgw�e�<i������/~���͈�4!��oJ����y��-�7��"5=:�
�#�P��>���@����N����C�6 ,��N����&}$l}�2�R?�W[�Q��X�kO��H�h���v�da�7�т��q/�Gٰ
T�q�-���T�����w�fY�����\�8;�g<$������%��v���-�m⦒X"��Xâ�����m%$Æڜ	�I_��Z/d3R���Кl��r�v��}pI��sV�����ӆ�׫�rw9�t�"E��D���o&@�7T����?�縬�J��G�t/���UZ�+�1N}ӣ,愃�W�<�E}!<'��8l��B��KC�j-3��r���������ɀyP������9'b�g2tHE��|U'5B7�K{����I+!����[c.���3y�"�D�/|�2�	@�ȗR)�|g�t���=x{��)Em	�}Rh�E�y�$���>��=2�r!�OF�E��fuiT��bg���F�C�4~#���mW&Ӷ�Q������Wp"Iq����o�Z��֚E.�DHJ�h�7�*_�tyUAki�������q��&Jb���ٙ[���t�;���*���F+�X�]���?�G�Q��VoCQ���.z22
��j?�� ��:�ck���z��^�� ��M4Y٩��Ӷ�d��F[���,O� �.➋�Tu 'T{i,�x�e
.V�I�þ��򰟸�"�� ��x����f~C~��/�R+��Q,~Z�p�B�z��$���x��R\�R���_m�F����Lk�"��NǶ�nw��9��v`���P^�r�=���k?e��.)��b�%�R:�B���Q1uJ�	���՞{3���I�Hg����f,|�����0lB��a0rF[{�����y0�/��{�Ӡ��^�c8&�%�$-D_�ˏd�E���O��"~��y3{�>E`xV�dc��5!-��8-�M��n+���/zUO����d���'���|Q$Tk���Y�*P�� �uc�yR����C�ޠ�Քqh�9��P��Z)���'��������X�m��O R��?�;�<���3[܉�$�0�!e��Ȩ���%`0�.�\KHL�t*j���A���	qac��E8�o�[]& 6�(�^4Սw@�Ρ���ݞ�����c�U���ߦ)�������8W�G�]eH��/f�*�ٗ��3�N�B�!��%i&敧[<�\g�.�N���.|����l:�$���c�Lٻ_kQM:�ҳ�}o$	q<�ŷ@�r�6��Wkr%l��j�� 1~7���q�*lń�E�Ă��Xגa}2�b�����4"�*�3�³R�Ń(ҹ�����19��B�c�t.&�.��G� !��t�"}���
�&��fn�0����]����U%�e�l����&3��k�_r������%3��J�7A�K��"��2���d����#�7����x8JT)1xT����zm� 1e��B�ܼc�v��o[v��u��QJ��S*_yi�o��p��"G��Jĭ��@X�ϥcu��CΕ�gm����=2#�Ao�1C�^r�̊������Y�Uv��QWg&�d*�q�|c�a�Oz[EI����uf��ܞ�]��	Ѽ�k֫���"6cN�)4� ���EHdP24�����7I�Q��]!y>�hu|�#W�m�Y$�tv\e�-�i�O�V/�g��U����/���T7��_�l������?cU4��{��$��*��b�k�,M��N�T/,�w���훲q}Ҟ}���=��H{��s!�g�<K�6TCeZVj��:�-@I�8h�<~�ܫ�Rh��?x&s8Zz���m�e��ؙw�`nr3�緾	WE9nm�� �����A�>U1�]�v��^EQg����L5���_��[��7�2s0Hv"�
�ڎ��f���ݢoy	�o�QӠz皴~!ޡ��֝��ְ=cͰ��:!�}��=�g�ż�/� ��6�Z�)pb_'������p��[��TOT���n�M-�]B*���\S���V����� f��<�9^�0��㧵?�~Nk	`w�E�߄Ŏ���}�|�Y�u���w#�W�}8�Ef��7�$�����oe	�	��ay��NY�K/Qu�/X�-��(�����naK#9_��Y}Y�B�� �p���!C�(6�S�>LQU=���'��]:;yBn���j�+H�)���4i�[���/h��q����Qu5R��ﶷ��T_8p�"�w��<^A�Dk�Nm�C�$	��^R3Ϫg� WV���.���ٰ�>R�)aI��O���6R�@ot��AO�b�-c�T�)PC���z�0Y_��ꍩ�Q\n�����2��'/���
 �z��g��N�b�66��sM��e.P�a/eG�F���CՊׁ�~\��u>A3����"��V�߅d,��Ǥ��.OS�����k��ˀ@�)�o��x�L�������s����B��e��i1�5������l�XK�+41��_���	�>!w��w�r�@=|�|�ײdL�xag$�GH��ne`;�;��r�i������Br嘹��[(����i"�A���Jf��q����`+\`&�`�|$B4%8��N�⶝~k�/c\�'k���F|�<c��=�ڥ�4�
�~q���<���͍f.xIֈ0�[(G��zQܹK|��A��*
GɎ�wgϏL���^$c�b%��h'���6ܰ�1���v,�W�#�=Qb�j�Jo�ۖi�Z�h,�@�"sY!~97:��+����喎e���Z^���uY�8d�u����D�=����+!�� �a��g��.�S�u�_��K�Y��?1ptu��݅ſ�݌����vd3���+�3$Y#h�i�m��Y�k"Ƴ�/&"��(я���/d��q�S��%�OSww��[\��`O(�?k��9b�*1���'��>�[��T�!B/�"}X��k�����ξ���+׌=�=���4/�����6Q7J�$X���������r9ֆ�5H���ȬtqfJ�ߖh>\"�9�������2X�� >�მޔ2��f��� ��逄섙��`y��z��n�$��~W��XYH��d�5C�.�[�/�&����Nf���|}���(�����\8z��l{���%6mٰ��,�Ӳulے�&2�q�dn|c��7�@?|)Ȥ�)`�ҏ�'Y�:�G���Ż�J�}���j�r+"gB|iKD$:t��N�Q�C
Gk4[�}�K�A�J�7��z.�.�>|d;��ƒ��h��cu��7{o�GQ��n̗UƑ�5K��$�"O�t���籗�d+�'��l �}U�@Ժ]OذT�S�D} >1m���>P�����!���0~�^rȅ�ˎ���K(��8óo�君518�"��]I�3Xx�>�f~�1ː�:��Ơ,��{fv�]�aÇ����nٛxC-�%�|8_c��5n�9	c9��j��7�q=lt�N�-C���Y�8� ӚT|�̾���R�|���X૴~a�ނ ݘ�����1��ο�D�lA1����3��|�/��@��!���们O�gڶ�����<Pq6��P$�.b��˼�\I��������,yH�*�/�,a���r�@�ħ��6�����������Ṽ�r?iɅՀ���8��+T�i]��xM^b!�.�\W;׽x|Δ��gkuI%l+�"�D�\ �yWcpC�l	7���%�/��Y3��O�وF���N[LK��u��l`�Ŭ�-�Mo��%JyKk%���T]������G0��y��H��t���EjsK�O|��Z\�p~E@���8�·�����!��5��Ey�����pQW��>K�a�!�IL���>h�� @���w<���l1�'��-�)���@
�'w���D�5�G���s�N0�/��Y]F\ܜ�[�g��γm��a*�k�>�n߆'�޻���������.
>�����Y����66�LA�~4e�M�u�u^�qYVQ�e�8!]�/�C�:� (���L9l�LO�<���sb"���㔦l����'��d:��)�tL~=>H*��2ެ�ԓ�O�s4�0�pm4�P��!�4ǧ�	*p��َ��4:�f�أ�׷��]���|�U6� q9j�'�/�Edzg�sw�q?~��������Aܧvc����P�'�^�%K<GF^	����eD'xnx�Z�'.�@$=�<������g�����Ib��U:�~���>� �e�^��elw���j���)T���1�QH��]��j2����Z2�ŀ��2�p=P(p��š����5 |"A�������*�_s��q��=�S	>@;���p���A\��ѣ�Kˬ����c�D�ft��
�?�%Dn��i9����k4�{%���Ĝ�fhk��l���r2������Ö3��;!B$�.����DA�y-�NJM��#����4m=au\ �_L�+��G�!P�O��K����b�/8³�[@91���7]�C6&,¨���^�- ����%'�p�^���i�RzHy&XΖ�Q{��1�(�d-!ZP��Pʋ{u<=x
M�p�!��<f��갋w�T���FH���'��XG��d�9�D�+@���הe�H�����{�� �/��j��1����_�^@,ѿ�~_�!7?	o�}�m7O��%�8�̒�A�ԥ����d�\�_r�M�a65�](B Q�j��]gm��Թ�ʘ��Ifm�D;�3�)��gzv�!B3��V5J�޲��!��l���bP)��݅&�?�N*��?

���>u��Cq!�V�w<;=�%<���>�YM֠Z��	���O��z*�
?�]�9p�r?��9ʸFlg�t܌S	�rp�CH��5�pa݌��c�{'�+(�N�Di�|(��=����)5ڿJ:�)ZzC��'��#�ܮS��a���wk�D����{_{0:$
B$��4ب�����%�ԃ�hŪ��?� !Ն=�c����I}��R�*��
������]�f�)��#�-f�_$qU��Vک�0C�ݻkQ��u�Y�σ���x��mWם�e/�R����d(��D�s\l<'�Ȁ2�Bմ�\sѺi����;�f�eS�x =g?�����\���+E^(�)������]����h§y�Y�^�|��$]\�Vgc2#��>(��!w:�C�1h�������ٶ���P��Q/bO'���O���O�/�+���h�D/	����ՑB��j��8��p�#��?��C���!M�&Z2�k&�r�I����O�ٗ��-�۲�t���w�ŔS�M���0����c,�%P����ߴpcx��S�+B������Y�����
	ް����L��zg'8��0��.!�!�f6+3�����vPVh��߅U�X���h~���X��oG�Z.�c�xc��uSA� ��4�r/�������$�>�����A� �3�B�������j�l���j��O�&�w�
eH�REhP�ʶ Ue�T�y3l�&�#�}Q\0>��g�����/@Q�D_&$�arlGO�k{�S�I��h�'���� �QRV�b��Cl&�u,��j���9���"�H�1������$ɎBSk�d��A�[��T5	ڭ��e�\p��������|����bNb�Hma�!�t��Q�����_,�Z���`��]ovt����1�͗GEn��ʆ��3m�ER݄\,G��Qh�J����$���<r�cx.ZgM�FE\������9��yo�\����%3Dm�����g���~V{���T�4ui�lv�;�v�A#�#+��B}�P`7.�O.�sH��&����8)QǇ-8��;Y� Jf���	l.�i�:�7���	�n a���@5s�P�
����U���k*���1*��G�GYrh����{�&q���e�����YQ��0KS��宐eE����+C
��ղz����	�J�I|E^@/%��ď>�r �N�y���F��k�y:�U2�b�,�O*wm���%�:���^�m}�����ܸ��'Ftɡ����kY��cTpOH�iK�<S 'p�q��[�q�us�.7B�E4�r}���`M�2��^��L���OSaӃ��;?K�p����i��&p`�?��9[2��j�<�țn
�h��-�{��^a��U�O��ƘD7fJ)��t�i�$W�G��� ���2aNh)�p.Z�=Y��ss �UV^������kk�B
wJΌC����U�~�%���Į���iQ��2�������v�.V��V�,<�	�?������>��`P|R�)8�LP1R����d�rh�}	�f��A����Z����=¡� T���܅�w��0E�RK4kW`�W ��׋mw�_Xj��es�;w�`���ʕ�o���-�.*5�4c�"#�I��~l�b-�"G�TQyA~�:����gw��x$*��)�or�-��X�6�e+�%���A K6&v���������X ��I�|Z̅�8��4ǂ�>��_�$}�����mz�\���)���.�N�wME��us	���p�X<_]z��,��)��Cg5W�YC/�%�}�_���GW����
�^-5)����D^.m�P��z��a�r)W�?b����ۜC��ZT���n�y�IVe��ӭ����P9q�����w�6J�=S���&��w����tmy��X���S�S����U�b-e�`�{�r��q�Ǟ����
KucQ����%���S �yU��Ǩ_�AoҘ������O�t#u���ޠYm�:����2�B�{��nAo��G#cf���L�m@�eG��U�*�o�v��U�!��㪾Y|Q�$���c@OQ�i��a���۫a�f��E��H�Q`���G`x�O�R������h���;O+��8&>��+��?��S�7q̴��N�<o&��?5��~G}&�M&^>��2D�e�_��*�A
}q�8L��[N�Oa�w(9��*�O.ü~i{���%?����X�2�Z��H�3�{�l��mϫ}1������D�>a����vÿ�d��PUK�������֪�(��W7˖���Ҩ���^}k����P-# s�h�n>�����<D�U�
!0uW��/"+g(7�hiZ��x�O�Y��ð��P"o9$aR��TQ�d�j��� I6�ir���l��:��X�	�=ޤ��v�m�j%Dh����'�c��[w����O[�1��7@��9�o�?��J��nUB{ΆU~@�������B���\d Zn�^���"���=:�Ƚ�YUi�-#�/�*M�l˦���C���_�8 ��~P�@��Yt��׾������� 4�M�C��pݸ����c'[R��`���f�:I�M����2�+6�헆�OJ�U\����h>)�V�{��A2-߄?8ɋ!��T �"n�̹öK�hː�Wy�l���p��{���7���3�l�p��Uda7������`������/�J ��K�{.2j_�o�v��]?>;h�yxD���վE$~ׄ��Ũ<F�I�y#��*P-��o��^��=�(���+��L�p�j|�l��9q(jض`��yG8a�Y�d�[c�.��4[���9�	p0a�+���ALE��<wu}����X�I�Z���[�����eW��4��~*��Z��z-����ÚY�W�*�,cA���?�9	r��wSh�^膴�o�lb=�8���U�:&�$7��9�3*SW[�L������'�f8DN�nOgt�sy�z36	r������q�%J^1݅e��|i��5	��|�j'K=
 4os�SxQ�J��j:2P35~o̼��� G�5k����7&u���^�

x���{N�ؖ��G,0����*�sm1nt�w�?6D��){��Ć%b�G�
���mW�"�l����Y�At�Ee��mW�s�L2�-�{�;��
�&�1Y,fF�-1�z^7f�G6���:��֤���\���K2f���ȯ7�q~��?0RBWG�1I3+
_��� �Q��J�.�^�St�N2�T�iA�i�vv���2z��&U	��m�x��"��X�F\;�w>���xNx񍢏q�'� ӓ	i߲Rr���B��υ6����w�}���� ��z�4�T��s�LS��uX��P
@Ě^��E��9��H57ۇ<>_'vp��SE ���E~q��$azDSzt\HH�\>�(M�"�������j`�[ph2��!�+����O��g�&tyJ�~�˰q�d��M��V�����8=�eLL��.�w�x'����K��#o�3���6Sg��@�X$r�֏$&���N�Ͻ��C��>�J_F�;����7��A�:s��ତ���SosR
���4�n�$�:`ú^&��X� �$"���rk9�`9$�EJ�G���~g�m�8.�1��K 9Ԃ�	�����.�T	�@�Ѭ UC��B�l�Gb-�n����s���v ��/_MnC#�@�ʣ=Ow�����=Jk^��j
m�~�����=��l"S
ܲ� ����Ytu�̠�s�]��a2���*b���1����O�b��?�}�@�l� U�P��[t�u��Ъ��)|݀1	�/�Y� ��;�̹r��9�!�<fd;1a��ZD���?�"�k�`��l#���)���^c��adg{2`�~�\"k<��NV�����#@b���b�L��Ʈ��j�F�N P�	���_�9�F
�������n��B�1ۿ3x�;6<��W,]��͸q�2����]۝�P;��� �9��7[
�"^^�-�E�˕��� K���OM���vyk�:����!����{�m��u���9�t�3��8�M4��5�:�IX������4�'� �>"�	XZ�9���3e�  2��aC���t�Akע�Z�#T��o��Yf�|FX_mn����j%�*���x�0%� "��뻬��_�O %��4!29��wk��,ȚaE�e�Gl����I랶�9��GU������Ο��S�i�5[�ךC�b��Wzax�*1>�.\��ܳe��C��<K/��:�Q�	w�Z7���9�^�	.�<Y�@<	�v�@�bb(��M��E�BRXx\�?�Khh9�g+qM�q��>U��{M�L
�wV��S�;����Os.B��>yW��~���f�?Z��VO�jݸ�Ҷ/�2@ ��#�(���ϵ,���\�~���Aq�s�B���z�<�i�:��� ;OS݈Uq�3��?�uí�B�� � ��L�2W�:�Ҿ�bD�%��(�WI��@����K��s;D'��Us���+�_��R(0cy��õ�=J�������G*�;�H�G u�+р�	34��T>����*�5$�lԱ\ó�(�&��٩�?�䐖�zx��Ӂ0�V1e���y�`�Bf֌hn�֨�xD�x�\Yʚ[g�@�����%����*�HGC���q&��$����f)!�RT�=��!	g��c"/���O��Kk�n�j&|��W1FH���sv�>���3�W�z���#N�d��5��t3�m�����)�κ�x�O�qB�*�/EC�`D9��	�0~��w2}�XK-����y���LV���˯'�X�p��
�6��hk&��Z��	qeMf�*�o���pC�ydsf6M��bҺ?���qW�lV��IB�M�#��G��Ϊt���i�'M�x!��[(}�Ⱥ,I��R�p�3Ĭ��ld7�)׈�f���R�m� ����@K�-|�oý�-�5K� �9B��6L������{��q���W�֬b �o�����9>.�{A҆�V#��C�ٵ�U_����t��28>�����
�1j^:b�-��5e�wR`"J�
�.�iz}��
�[j/6�Ɖ�a��� hO��(	k.S}L��̮Uc�HN.�;�e�����?r�/I���YN"m�pF⴬o���<|�L�N�N�������#�%*�L1e�2�����R��^p�wb(�d�=�a��ޥ,��]���|v�`���}�=�������x�u(�+��n�$�0��	&I�z$�Ȅ�i�r����� ��-ĳ$kq�������M�sJe���B�J��]H���ZКu�r��1�.M��p�pC{��qh'\������&�ʹݧ5����|�� �z��6�~�U{��2�?h�C֡��Z�i�F�� �_��AW��W�q��y�6���a^k�$�ޭ��~Ж��ME^C���xP�_&�mU���a;]�Wo���u`����O~������gda�qOrۀ�5���i�x�)�&����U'T�X�$}Ԡ:,�{�3`;�B7�n_A(���=������#:����Սyg¿���c��F�7�v��%�a�NqHCa=��5�p����*U���'������0�U�$��r䙮��ԩ,��<t<Q0��3�蛶Tz>^�t�K؇�#\�G:;��2��� yp ������q��ԣ"T��!�����!B�V�:G��֫�2/�5Mh�?�����@	��[(O��j�r|�t⴯�| =Sږ��F��Bq�Nw����l����E�dHz�����i���-��10U�{ti$�p����|�QH�h�&ԋ~Hup�6G�b3K�����ͰQ<'55�Qn�%�߷$1���������e9�m�'ɀ������%��,xVeHi��E�񺁚f�2=�X#�i Ȕ�ܒF�M���Ή6�� V����\��xr�Ԭ� 1˃�L������jY�����x��dS]e,��mM��j��Ζkn���Y���x�Fb{�+{t�j$H�8�3\�_�=�+��:ΆLk����p����)l��@�r�Z����M�Nv�~ �={�>�*O�Ta�g+iĚ���	�~��d���jT��&���x��CJ��C�s�[ѯS�_Ŵ�AϬ@ߺ��>��+6������4�	 sB[�d2)�=M��4#��[��wg�5���%5i�4�-K#X�uk��ub_�(Z��h���ҜL;%a���~Q�dk^�Vm� ��^'��sl�A��4��\ܑs�Z��pJn�����Z�Uc�	!������b���nm#B���� �Z��+��$;��;r�_0//:r����tN��ߚ>���o��rl�kv������TR�rg�e&���#���f��scĈb�o���|����RIyT�:[����+�MUƟdk�]Ɵ+����R��ZkN��k��j�<tg+�xw�er�%NX|X��C���(,������i��6n���13d��P�p���0��҅�`(�0�qv�и�j�RB+��_��y/ԕJ���-w����y�H˄�?$4��Y��;��:�|<�`š����_]vgξ	��Y������E	��ֆ��e =Q��V�؞;P�x��� L(��ү|͆4K�*�3ɷ~�;k^[foe���lI��B_��2����A��|�&���lx}��K�h]��:���h�-ml����l�R�� 3�⢇�.ag�>
����]\�} ��l[��'K$J5O��{�-�nK֯ķ��^e�m4��>53�����;J���a| �z4-u+�?]g0���T��<�ļ�� ����묨�ey��NsH�6���l�R5Pɏ��0�6� � ����{{��~B'G1��""�T7���:��m8��_!��\M1#����\�J$!J55!}(� ��WriRw��D���"x�a/W��j3͝��F��]�a.&r��i�v-oxG����l�����\,�NF�S7q5y(C�~Hύ2�		=߬1k:�w���E7p^�]_������/Xd�����h����W�����db��e�	\5H��;^�����f���Y�@�iIs��G�J���aMg�bq�_���aة�����Y��pu�1�t�&S�h�5�b)M6}cs��C���0�/���f�{lBQ~/��~�C}4�����RLF����J`Ż�'��y�EX�|k\~\|6�\��\�Į����^��L6@D��rm�hd:�za��wy���͑,�꤯So�4cS�qi�|�j7̢]X^ſ9�_��dƃៀ��}]�,�.�j4���mCj�O5��o��H̓9@^%T���ZG`���Ӛ�)����J\�P0�::a�5Y߬P���]�׻�����<��Hq�	���O���z���l��c���L
!�n�PQ�E�A�]B�u,Mc��F*�2J��6us�P�\�]�f{o�9�IT [�vf��������ES��e	Av0vcmb��Z�}֬Z���\)���f�7�Ӹǘ��*�:���kC��C�^��Eujex㚛.¤	�����=�d��ĝ+�g���1>a�+y�I��X<�b�γ#{�Q<9����i�x�j�q5�ќ��iYx������[�[��<]�f��d��Ğ��z�C�\���/�J�pJ��,,;�#�E���Y���[)%6@��f��I��Tv7�ˏ�s��ȼ3����o��,V. h�ѳ�b6d�?��axU{���yGF�� Y��x���Sqq��{X��`Wf��X�J�U�$,�)n�Z�!S��q����Z��i���C0�Dt��7�� qE4��	"ʣU�c���Cqͧ�z����Z��n�L��7�eZ�)qt�hi����#f���T�^]��oQ�ʈ� ���WZ��`����A��4|i]b�v�!Hk�t^k�F��w�MfY�Ƨ���}*鋋r&���-�����/�Ѻ�#�o�aq�"����>����g�w�x3��\��We��O�9\�X��$A1�K��:l�_���쌐��`E��Τ�	]Z��@;� ���	﩮a�y����I�k0�R�E͙�����ߗ6Ĉ��i&K��EF_���t~��db�53>t��Ob���/4`�ۖf�N�@Z���(~o�ͅ�����j�����[���>�ɢ��ZK�G�������O���˛5vӾۊ�'�2�[hݴ:硣�V�-S��q������}!7H
��Z7���6�m��0�{�S�L9W�~�2#�~�Z���0�#r��Qwo8������$�F��Cvh��T��.N���N��l���*l�j��Vr*�T��Vt�S|mi�@
 �����f��H��L��HN�ܡOst�Rq�9�����N1���¿�a~rS��`Wl�|Z$L�c��f���bh;���]��uR��Q�tWsҷ6�j:�ŧҜ�e�l3{�j�FϦ&a�Y��+M���UV!�g1���V������}�d��P�kk\Ee����x�.]�� &F#�+kd~����N�G�mY����f	C�Z��#:=[E�a�Сcv��=:]A���7
�]6�_��X�DX��o3��G���N��fJ5
�ybw�@�۶i����]�����ƮI�u�x���R��b$�zDbG���ʅ�o�G;k�Q���s�����mӺ�h��"i�`�ؗ{=���;��|M*�в��K�7��jh���O2"�܄� ���N1�w�ezr4d�A�^��7�)8��l{f�O�����T��s4�P�z� �fRY�\�"-n�pL���D��/%a]�"�dwc��q6
y��g&)���{��fg����fRd����i)�G�o{���}<'���&KBډ��acޟu�S����cˊ����t�/P6o���(�dA�疻�$����=1ڦ]c��T���:Ւ�`n�7��qŔ��x`�����c�'�bI��B����30�i��`{�����gl�s����
�^d�9�P_Z�[FZ2(q�r@���&�-V!���6�Q��y�߈�<�f�_����J�;��{'����jKS������J��
G[ͻ`�F�&��":��-Y��7��_�Q���Ȋ�"B+��5�c���
�.�[�]�2]�m,��{��AE�*/�5v�^�qUPH����D�������`���]b��a
�o�]N&��8x�|����&�eIgB��pPU��w��D�{i���ox��{F^������XB|[���{Q�����z��|�i0�5��d���A�,-�eNd�|58�� =!�`2b��=a�V�=ʣ��J~�m ���K���a� r��������ڰ��ց�?Q�d��xஔV��x4��L)Uɹm`c�IYL�dt�\&	r�zC3��i�n��R(}�=��;��eka�?�T`�Q:d��8�"=����>�̃lۨv۴�����=0'�ԯ����ŀf�� &������.U���k�G_�);�L�r�8�����J'JY@����b�� ����,��kAm�4P.U���T���l?�W�Sy93�vȦ���m�V�^��3�~d����V���ɥ�4C[�Y,�u(�E+Y5�W�[cS�Cs�U4o�<��d�Ϥv��-�����09Rّa��'��$� �5��]%����A��҂���n����ֱ�Ĕ�3`PlO؆����]t���R�O��e��ro��.A�b��{v���o5&�/CN��<�c:��/nm��:N��<�Z�s/�C�:����^��V�5��,��TQ��˳(�%��A� ��E��t���W���71|�ZG��jR�`K���UR-B ǁ��(D�PF7��Y���h�5�&��Mr͆�=�Nv4N)h+���iJ8-U�S����� ��L.�_I�)T��~=�LN�qXp�R�
|�53oADD���};�	W�9HQZ�MK��sϚ#хЮ�p�zMU��8�J��֗�+k�w$niճ�\�!�W5�sC����Y����Q]����43D���O�Z&I�o����������Q��#�h���V���`H[ݘ�ӟ���=Re��F��s��	c��z�3�g���t-g�����z������6\0ϲ�=���Ft�r�SD0�b��;U)��*p��p*�y�����,����`3���&��ƻ��RZ������o|�o�d�UOb^�0?]`��Ec�r�L�4/�0첡Ϟ�L�GN )5��<��3��X%Z6���]�rEY o ���sE�����E���u��}H��	������+��Mb,�b����_��Ǩ��ip] ��_��������=�}��p��C7��-���eƪ���~%�z)���(�|�����@����DE������9�s�21_WC�H�n�e����?m�]`����<��8���	��
e�O>֮�*� ��~��1���f=W,�ͷ���h֧�H?bO��Z�)�M=���4BȘ�m�'��yZ�� ��TOl]�%�[v`�&�aB�3����}{���[�#�8B���E%˼a���ϑ߃i�-pϪ>ƤA���Q�h`%�c�,Gl�jl�u�S�S��W�-u����î_��g�X��D[1���DJv+s���^��$��̿�>��çuK�}����p��5��Ӑ_��ϼ1�]gx�uD�S���0o=(̧���R�8�-X-��h�ϙ�J5	����js�K��C_��V��bt�fBq���k���(C����w=]-,�R���5��P�gФ�Z/�˾N�,���3���a�n�YHϡW�	p�z�;���Dcy�|���r(�A��"��3MH��_c�)�`�%pC���Y_4���g�mz����L ����T��!���;��4�EVA:�*tK�>P�u��+�k��Y.�"p�I���{��ܙXI+�e���R�xZ�^_��0��[�2,7?��)f#�(%l��~5Yl��#�Ҫ�p��r �NY怗&��ߤ����n�{_<R��"� ���o����'uզL_��N�2�]�\���
_�Ze$Ư��v��1�W}�E��i�Bkv�6��g���+6�ꅷ��ȭ���'�Z頻]���e��&��C Lv>[��"��8G%f.h��$ܘk�fg�ƃ7��vzћT�߄6i����B����~���Ny1�g$a�Unع��Sԩ��&ׅ��C���G��i��]4*b>��F��M ��i���|B�6)Չ<T�M�XKl.���_�L��T���v�&i���~%u�X�@�F�)O���ؤI��ܿ���������Ԛ2)N׌�=O�C5�)г����_�r���	�)l�x�D�I{+T@��y��MfЕ���b�� �o��H0���s��Tk]�E~�'��2�p&[���˿�"f^�Y;��g�573���vk+���/���ִ�(n�~ՙ�a���}i�R.
�{��n����X��T;�E���B��(摴�+��8�K��Rs%�#e�즪�(��e��)��ؕK�3��z���bM���K��)��|Tz'��pc�;��ӯT��nY��Y�M�N�Kj���I�)q�J�;E�� �o��8�q�� f�[i���D9��O��a����>u��(Ĵ��V^�&#�������J'�Ā���1�����F���1��5��v�T�껨��h�a?���������M�Ǵ��2�3�7���c�p�@=��&��b�cxQ%5�n�)����L�WX�S!�濒��COy�*Z(?<e��-�����8oW� �g�sY������>~���Ux��� ����s���I�י�x�� ����HS�9�X�A����/��]e�t
�!9�>�9>l�zDŅ��W�4���BV���J�A�۴2̱���$��C�#��ϼn�>�¼���������b��ʝ���Az��?���)�ũ���o ����(C�!�a7tȔL��J��(˨eqkԧ��G-�r|��p�����s�u|�O�_x<��(�d�z��mΤ�!T��m���;�������	[qo���֜tKYp�)B�&�^�t֌^��i�Ef-I����2�q�lK��ױ$
�01�#�p8�l(��}%�P�~�Xo���s�]��21de1c[�⧭!���;ߡ ��k���=$�@�|�_aP�1ml!�@a���ob�$�s`_��9���6ʢQ�%��8�d 6��.?�ݔ�a~��P\������h]`Z"��K*��o�Gu�7)E��%���;�	N[�`�"9�^��`����~��"| �O�^��h�>X�hr�F�`{����H/�OQ�|hi�(��lHoN���5Kɞhh&}��7U��|wqK2&��n#C��u�������>H�rg��u~�.�KQ��6y�;�h�T\J�`�><_�~�6����˧$T���V-?'�q�٢T��4:E<�x�� �f�ܯ&5¸ΊQhbx�Z�?X�l��m�&K���hmD����f�3s���8�A��r���Z��J%I�;�"1`^m<�`~��|s��6�g�m�*���������+xi�
��t��4�Cc�L���*�4��ŦWʜ�C���%!���@'K�rsC���&��N��k=��1L,�@K�+�h�n,�J_q������x ��
Ž�|EwJ���!"X=å��O^�P���pz;��{L�=�"Q��8��[_V�*���ܐ����V|/i�8r�g*�D=��8T��,��{F���9�����p�4�곐g�ީzj�D-�e4��Z��l�l���vh4k����i�.59d��:+b
����$Qg�� NuT�c�$����.������B�{���	K9��(7��1+�År����t����x����b��.Ya�tiK�,�م���*�b]<�c҄����w^��~8!n��\M�o�V��NQ�ѩ>s�(_Xk��a��k'3�pl�F-�V�����UY�5p��yA~<Jw��TD�A8���W�A2fŰ���c��#ߚ�s|X`���:J&j���Z8	.�[���5-8d��3���t�ҫnq��1��$�`���6ZK"�c�����H������A�(ŕ֪��dpM�@���J�6�C
�%ɮ�aᅘ�Њi�>�>�m���G��_!e��{�X�'�z>���{V3��_8��$ɀ����7w<v@�a��`��������i��݁y�4IזJ���vo�y��b�7^�cN����;����N!�"-���t�.\>z�������*�wӏ�An�^�����m�W�a{=x�}�cF��Ruo��W=[����d�z���}Cg��V��*0	b�N5��S'X��qV�R:�n����c�vR�)�����,�3� �x�[g��?�]Y�r�+1Ǽ�A�P�*��B#���CϏ	�nY\
�Z��4�
���C��:9�]`�i�ҿ�#�B�m&��Z�J�8& k�Cw��ML��=;PB������Y����ǥ��`� ;�GsBk�H8*2BrA���S��.uz��E8�頺%� �bqi�!|���ӓR�R�ep?��j#t�B?�AF/m��;{@�~����B�|O1���]�������4"o@��'��#:��23{��k9��(68_������Ԡ�?���S�AR��֖���E2�%�U]Tޫ����#�[��W츨K5�R����d�o�<)�ϯ_��g;IaEtQ�/<�j�$i�L)��������m�����w�n�o#X��FMS�ܭĽ����4��ڻf��5��y�r�@�P��P鳰'���z��t���^G�C(x���9@h�F\A�}��4���ϺYⓣ�E��P����1W������Kl�)��z��i#9���F)�5+Oy�sk-�Q���p��3�9����wTR�S����B8R�r�_�؃�MR�*�^%A�Y��D�1G뽢�Q����a�"d�y%��U���`*�,��e�܇F{<5c����c���4�_�W�Wr� 8&Tt��N�C�,�Z	��o� P��e�ՙ�n��w��?	�&�Ccܬ��E�:C�+S�wf�U��A��@0�~�EL���ԅ0C<��f\Ғgȟ���w�҈�_�cb���Q5W9�oo_�Nc�����=��js?�@8�r�xřIɟ��<���MU��c���wc~� m�1P��`��φڼ��-��{�xP_�$Q�>U��"��dH��oS1�t�5	��BK[�F}��ZaQ�����9H��V\eG�`QS$'_.b}���7] <����ai��k�n`�0芗nh�`M��,���3�I����X���Ҿ�1��	:l;�(Y��{��b��Y��Q�r�2�?''��=��K.c��YϼG��!����d˛Mb|�AA���&�l�=
�H��!`�}�5���ӽKݽ�����'}& ���|˰S�F����PU\2��AK����T��I��;�����ʿnOH��k @���i���K����0@����_�O����yJW��޾��^d ���N����H
���A�B��4�_�k�H���D��QI�w �iˇZfuF>�zU���vS�#��L�ԏ����d�*K�L�,U|���e��f�a}T��^m�z����G����:P����r\Kk�},n�Q�����*Ɇ�b�� J�B+:��L��f����j�sV����ړ�F1�Uo�LwߒR͉� >ۣ�O0�zX����}������t�G{��]T��@��P�Bi{c���s'�W˼%�3nU=aC�zY�v4�[�O��0CJ$�>lk���5���Lˏ(�,WS�w09�$O�si����~�	4+hAR�:�͉����j��������céM�����g9�6Lf� ����b�wRY8oQ�;��w1�㩼��:<!���W�3
���4�Jb^<���W¹�γ�լ��-��g�@��^ck�.T��/e$�#w�5`��9�DK��Fz�ZeC�@��w�̋�px�,a���ō$���@�PΨ���Zz�M�Op����W�!ѫm�&ЛUfR��?���8K�ìwO�M��=%}�Yu�����L��Z�ݭ_.]���%�*�I�1�� �82B`�t��c�[���u�Ss����C=��Ʈ�V59�	�aq�{b7A�)�n����k�bd�n��"�{v{�'��ų��#H�ߓ	n���@X��9��$\�W;@�p6?�<�i
&܄P�Ż�������[,�����Fvj�(�U\���.F%���\���k(��fU���Vߜ�02-��D�¬P��O�����*��ԋ��O��[y�t43e:>H�T��z��R��|ޥp{Ѧ�f�`G2g��)�Y+;��r�D�B���Zs_�kN��S���	�\����_� ߾R�0�.k9D,���8��cV�cϤ+�2�=����Wh����i_�jW�4�5R�"1����(�Jz�!C&���Uq������6���a+<���L��䤝���0��_�('���W뀚�4�J)�=u��;3���m��rR.��ib��[ ������&�D؈ud����kf��m�j�su�����0��ѿ��Ҙ�J�~����o靏�}�h竐�PS5c0���!���ӎ�/�S�Y}at��-\fN�d����4�� �n����i��w�L�Es��ا������a
�RCөx��b8�"�Gz=��|����,�׫e2�>n�O���*� ѤM.��ӏ�$C榻��D��>�6E��5�������4>��M=C9h��4��gpX���Vx!?�<"Yk�Y� ��z�T>��y[K{Q@=�A\�����NoaZ5�����D�X��`��(�z� LRv��`_椣��Ы`
3�z���ˣ����A?E��";n�:��\"&C��/PX�k�e�&�����2��yI��+�J�#���.5��5d���|�14���;c��7s�H��Ƞ����.a>�����v��3i���Q'�d��S��=���ਜ਼`�#c7Xˉp@���1���o}vB��?* �J���a�:���9��|�\�e���%x�~0, ��|�sţapj�CD�Z��X�N�����z"z��</��tɢ´.���j�Kq�9�ܳ_�@U��� PJb�KB�;�t91I2���BWtây��I�d�3S��[�V��m��X7�նbÂ�OG�N����j�P��d�ڍt��}�.��� 0�W۪_���JN��q
$����(*������� ��-���ӟ��ֶ�k2d��({&���ⓟ��nw�O����,����V=(A�W�˘���r[��$��z���G���B�8t�?e)aH*�<�6���'�[��sWxJ
'6���o6rw��3$K�
^�T�t���f-0:��g��
�8�7��P��RR8�_��j1�av�o�~�����E`�(	e�����P8��M��=7`pa�;�ԙ!�r%�����c��+hNn�y����WؕH����K�1ܴY�}]�g�,����.zˣt�~��Υl�0V#�R5_	9���.�{y�t�z�����&��u�-���Ձ��J����8���dG�C�d~'e�'�S�A�[�;5y�+��'A��葯q
8?��K4��iBe%5��T �u��z^���#�Y��v-��MM�p�"�s��%gYwf_��F�)��Y!����o&�JX��e�����nG��^�˅��/�@.����+��B5���}X��Ho�a]DO��M��g̢Z��>������k�5�ｽ)~�
�=��S0�b��tZG���[t>�w��-�(�în��o�Z�cU���z�,�s�ZP"��������w9y�@J���(Z
:����Oy���q r��F��>�h��L�b�[Y�PH�0��k=�D��ᓮ���e-5��S1��!��Y�Y���+���x:f5H,SwQb��X�#�n��j��N�Ls� �hNYwM��ԫ/v�b�6��D���R~pP�]Y�����]s�H=L�Z^ϯ.r!������g�}z!`'\�źJ�����v�h�gPҐM�_��^����
+ܞC��
�OV+��.���H�oe�S\�[� ��y�Q����D2��y����h�{�j�W�;9JM4)��:�r�`��{]8˺�o�hڳ�����L�[kZ
1[��CUa���s�QٴR�+q#}���������f���7��E=�L���O�DՑ�d_5.��B�.����n�_!���D7�X�.]��?K*�Kײ�\��)���u0S���U���mq,'�y׸itf��#�\�<V�Y�n�/k�I�- Zjy��~�$>Q��b`�ld$euu�s��7Ch,���@��~}���#�!g�x�֨o��sq
��C�UǍ��=���
����q!
�h�\� y�g����e�ׂGL}5�P����ur&_(���
�>����C��D�i��T��mP���i������S���Y�MĭՔ�eZ_Ai/<v������Ay(A/�o� ž���Y�������EUs��#w��{�e6��sV~&�E!�n�2b�8�C>M��
��WΈF������K����t��A�� ��14�W_�w��a?�=���l��w�]��4e�b����M��Yx][ȣ/��CH}T�@ɳ�(��C��XD�{����oCU��r�m�fɝ$�|����6����c�l��np���*e �}�l�3_]��Y�sG�p�fB!Z�S�io7�r����3���Rԯ�����9��F�z��H�	� ��kȽ��P���{��|�͇����߸�T뢕���X�	!?�H�7)(+��zQCwl��=T�J�ͫ!�#Q�X����o���s�rR�S/h��Ne�Ek�*�����F�8DU:؉�Tg� "�b5#�3?��.d�n6I[FH|�zp`ƨ���E��ZO������T��IWR���ﻌ���B��gX~�Q9���	,+���#{g��p1�R�s"��b^��hJ�>��a-���>
�|�Z��Pq����y���>�É���tݭb�i�M^<����UC�=m�2��Y��q��(e�~�6G�#LH{mϷ����l�>U������'ɖԆ����in�����WB��۾�s]\bDD��+�%`52�o�g�Ts�F}��m�&���4�JHqD����oH��a�fƦ��(�g�Ζ����K��b6��*Μ��+\ZM!S�/f�
h��Z�9�O/�x,�ymcP��Q���l7;哰g{���	s�~̸n�i�,�Ø)�8ʏ���QN����F�A5���n8��Wd ���6q���5bEs0�_������@^��i� =�aM��C����Ԍ�X$p��n�$�x�U���N:����ɋ<����.�H{!�<j�Y�D{�B��r�|����I3����&��4������(���[<�"��l.���F�̱� <g5�[>���kQ���d�tR�"��ӬzI}��̩6�ӵ\�g�T�*e��)p��i
oU(y1[v)��r�w(�xT2���7�W{��+O7D�}�I�{4>���S�:�%�VR��I�Mܓɂ��&a��뢣�]��S $�NK|D�����?�R�<���� ��a��b�Fδ�a�A�U�	H�Ir@�_tF������1��O$�t#w������3���{���[(����g�ZWBR�TY�4d�}�ǉ��P�<c�����,.<� �V��m�9�b(0نE��ĩ�S���(k<jS4��	XU28���^۵��H�d.�pB���QB|X)':x���P
L}<�X��W=X�h�ֻkД~�dpcE�3¼�T}q����roSuN�U{�@���m|*�$Үe��.�̈�!�Ha��I��n�}{/�ϲc<L��	4Hq�1)GĐ	:?�TQ74�����=l7�+9T����.xe�VF\f�-B� �_}���@(�ۏ�Wb��hܷ��H���<��p���\+���;sT_ ��v�2���x!���v�����U;��Gʈ�(�!f��+lDD¬m3��M�YZݫL_��l*�`u9�q�4h�fb��i��*,�oe�����Ѱ���ٌ����tH!�����X��ٙ&.��X$�NT�(���ǎw%�
sz���^��O~�$،<��i�w��;k�ju����n�~,���&�[j+�]⤃��!(����gkkQQ��O���y��$m�r,G�J32�ͣ"�V<�����8�׺�G�i	������M��,5�~�dZ�{�՘���<F-ǎ�KԠֵ���<1p�	6q�F-!G��6��e�zt
� �V,�׹K�5���5`�&[M@o�!��\F~Z�:�A��Tf3�S����4�k(���/+��qˁO�7r�-�@��s���˦�{�������]b�֍��9�6:l���C�t|5DR��ՀW&��	H�qK��
9�!�s$c��H� ��R�Q��|Mkt�cr�HX�6���ؕKY��S1�Hz��%�j�������paAI���s��F�����f\E�e5y����������t��I!�;z�V9OD^��_��C�
��DA&�9rYTM�oг��>�@`�;W@2L�]7A���n��]��Ό>����h��b	_�BX�����
NRA�Uk����Sj���Yj�>?�юuJ��UI˰4��rDWI�(�d^�}@�a�af5l�������(iŊ�H6�Z$H
p��+���l�K��!̩T)�Dԝ�Ӕ��P��l��k��x|�V�1��q���jeݯ��O^TS0/�~ٮ���uV��h�ڵ�%��5_�"l���R�v�e�X�=�!���\�
��֘�t�Z:�R�a	�cM���2�����Aoܿh�"k�F�S��Fyq�`��o�;-��*�"},��]S�)w�%kJ���2P�ըW7j�"ہ{e�	�	��� >j��yr�����Tp�k���@�� ���̑��e&����x��*�9���a�hS���E�tέȡ^_�3���.��pV���o��06R������QZ���Zؚ=eպ��d��}�3�ϑ���a%�[e�WE M`�j�y�f��{��u2�VU�`hoT.��qX	��\�5h2�֟�����v5|�=Q�ֱ�>*���A%�;���eu`�p��h�f,�(q�?gn_�ܳ�#�h�|�M�������𬜞��.��7����(�1,bg%��:k�� :�CZu�����b� P��F�&9g�&��ysE2&�f����@~�>NO{�>P�t��p�t!�%9����6P+<��t��� ��@Mޣ�}����2.�9��y�2Q�4�U�x��{�>�-V��%9���Y�Ȳ�3xv� wo�����~c�S]g�60-�����n8�(�6<v�f�� �u4^#*d�0z��w>�ג�H�Ju %�]7f�������=�
�q%��n�r�]c/\7k��qx	���ZQ��T��D���~p�nX���+�Bx�&,3㙪(���\���{~B�uѝ�19���Yab���3�����Q�:hr�� �Γ���0�7@
{я?%_Y�$��>�AZ�[번�4FYm�]�A\m���N���% ��us+L�9<�L������/m`�D	%�Κ:�M���*�|!�{�t���>ǣ���ۇ�&-|��]N�`}w�����/js��X+�`�*��b�[z�]������xB�>8�OK�]j�P���4zo�ڶZ��U�S�FUN��De�������r6���2)��Bo�T����|�mW*�EX��k�k�������ݜ�\�c1^�<uA�QKv� �S��@���(F���v
�.ER�n"hE���)�B�q�R�Ʊ"H0W���������n�Y�a?�1,���=��<S�SozO��&�S��{G4��#�[A��ӵL�BX�����00�n}2��g��^�x�g{�.���Xg�X�`�E}�$�2�7At�^�TxJX�%��Ȧ���!*"�)K��k(oT��&D7����QEX�v8j��W;\-f��Ez�aBH��'#5�=���V��ɇem}>'}�i�_��ن�Õ+�(�hk�W	Gn};
*Y��ŮC�[��/!bB	��Á�'�Qs�w@X�E<vX2�W�bA�1�z��d�&Y0߱E+�0F6�貳"�n�m����P���Ē������&|{ ��\�C	�)u��t�ď[���B����b{�&%�-�ER��d��ptGw�s��`Vą�x��F0�8��+
��U�Rx��mOoM¹['^.A| �`EQ�8b�t�~��`���Ds`ѧ�WZN����H�Y �3�9.�xÝ;�6�g��q��+����1(�!!�B+���Eϔ�����R*���~�c��ζ�R�i_x4o��{��n9����Cդ�!j��x��uz��'}�d�!�ꂵ]G�ra(�c���yr�Fu���D��3Y�؃n�[�7��Hg�Jm!酥����n���N�h�S-V���g,���=�A��M�P_o����x/v��w�c��Jϱ�E���Y�K�{���[�y�`�c
�����pDQ���x[V�fH&��&^_�('G�H��|%���8R�ާ�����=��<��w@#�Uc=B���m� �p+�$k��]�Z@�m�ж-�9,xWk�U�PKaX_�F ����P5՟�RĈ`)��)!kDP~n�1^;���ʒI׸�_Ahda���6;vHeF���FO\~�1tHN��P9'/�����=x���i:`;)Ow+`,\ؙ����Wx�c�͝T��a^���򃑃6C����
#��_�m�@�K�̟ɥ'�F��+�'n�u��[��m�_|;RsF����s#�"�ۻG�q��=��z���p� C�#�֮����>��h���+���L��R�֜�F?.фP�c�����J���V֗ǥg�3/�U�T5���8|�!
�D���������l�.P�{�eʵ6�i-����nn��,�r��`�|�R���s�I�u�eSCN%��r��;	&�+b7��ì��5~>�W�~/ ۷1��V��N��Uꭓ��!o
���K�+�0�oq�c���I����$��m@�h�[y�C-�|������֜��⭊>8�8���j>�{��NլI�o���po�(�f�紱TC�
Uc�����R�?�Y<F�s����2?n�x�/�Y�����)���x-�.00���/�
�Ϫ�I�H�4��}~w ��ă_�Q�t���+5�H���SR��ۣ̘��2Q��&9�G8/�v޸�|�A�^ڄT���{DvC��̧�үǜW{���f±`ҳa
�P�ݧ��,���)��M֐C尋�t<jPf<�A�'��18������	R?	�=��3c̫����Ie޹�Hx��G�����y��O��'�|�D�bi�uE.�90�v�O�2>;,Ay�炳N:fdp�Cq`ĭ�u�A�v�!38����{�,�#9��m�6g�F���JU�$[�;U�7��B�I�!;p���R���� �=���Eqy�U-�U�������=@پA8b?+�Mwܻ�p�Z[�Uƕ��P���𹮀�!���4J�J� v�9��� w�&��t��ȹ��"�?o<��}<��tm]���<"�Z����� �"������}2�xq{�1�ONt!�|��Ӓ��+�,� ���#$l��=� �g���Q%�[���=W-S4C���������t�������M ��_���1'��\h���<hpp�fm8�why�\�d�u;��(�J�m:�	W姲�5G�+0�}�4fe�$������h��P����6ʽ�e�����9� a��P\�����S 4�5@�j]F����Gꀗc,v �5�Sx!��J��K�[|=��5WfO�k�z��?8U�n�
G�PKAY<R�#z~vF�n�O
^ԙ�F��./�w�E-����t	_֧Uv����U����N����cCtn)ѫ�GdU=�c����a�Z�]��џ���܊��T���nV��@l]rH�=����Uk=@��y��Z�^�m#�i)f��#Z��LCKk�.wlf��������d?Q�ga�+��ͻb�?��ԝ��V��{c4��35�cd�s����<P�����
g�+ԭaY�8K��T���3�؎����\��0Ʈ���=�wzIߩ֌ ,�3�]���j�Be)�Cd!v���0�=�Ж�� �@��)�����yD%:a��Q�5���o8���6��7N��T!ױ�P0F�NeJ�ϋ?R�A��ݡc-�ҩ.8?5U�_�w7e?����a �v����U��\�v����m K���ke��E�<3]�jɒ�%��^sI�CHG����&B��N�tO���h�J�)��~M=��{������PRˆ�u¡)$�tdG��-m��J/LX3��=7S�x�t��v&�ƯKw{��>�&Ϸ�"��A��h�]�i�_���"�!��t��t���Ii�.M�@13[�ze�p^_i���3��'�7�x��`zc27�/����~�pfM	� >�ل���'R���#��˦�&$�3P{�t�]�R��2�CM�Rt(��-n�ٸ�YË�N��}h`����[��T�1���J��'�`S=T� )��LNv8�r�ubNc��еTwU��>lݗ�{�p��	����;�7���(���q!�ZI�L�����r��T{ �R��|5�|-ɭ�Z�`G;w�Yb��.��ӥ�`�{�1�y�l�-iW��~���o��ςs.��5O�_�3��4u���q*qC��)��d�ژ����A�nT�#���ǳ��U��N���d��#f��h��pm#��&����F%{W]s�1j*Idf�Qe�ɈJ�g�݀�D��!�~vZO�Hh+<�i��V%:p�^��Jn����,P�qX�^��P�խg���W���r��AU�4q���	� ~��Տ��6���k��j��y�(�8Ѹ5>�δ�E���Q��)7p�1a$^����P�� r�2g�oF����u�c'�9�Qݜ��ߠ��p6�mn�3L4�Ӂ�VB���^�t+-���i'eE�k�R3}�q�	�۫7��O,b1M"������%&W��|O��Qnƀ��72����;mjX�n8&���B�dK9�8����)Z��1_�#���KB����Y������I����"�����Sj�g�V��<��]c
�M�m��u�����Yd�ď��ҿk]Xu��1�FK��K
�Ԯx�� &QP���wE&�����G��Ui$�|�$Q��)m��Qr��:u��������aѯ�#=@b�d�m��kq� /ú��Qs�1@�0���7��T
�*E;"���Wqy� *��͉-���R6ቱ!�h@%�Mw8��w�-h3Ț�p�	X
*>�?w���zH�f�e3=�2��_c5j	�*9�>{ 2t��8��Դu�AV�:����.|<1��O�P���1�ò�f���7|�f�g'p<�����㴕gt;<��I��;h=7ξ]�wLU�F;�O(�8( ���	�sê�Qe}pz�}���g�
 �-���Oz�(��O���6b}���ڔ���c��χՆo���\��u�Ü�N��qt�R��4�������	�[C��ZW��7I��Zf�uM���[�/zO�A6�M�o�<�4q@`k��41��R +��~`?�FK�eIy|��ߓ 5^�q��/���)e=�"���&�T��<�p\Xr|�;�4������#�ß�Q_�z�Q��m#�������7֗}�� �w1��Lxs.���M���P��;@���Y´!	 �/lc�y%��b'�|�R&�a|k�&��l*�,x�'�R7�[ &j�M�U9���3�k�������t����5�h5��Y��7��l�#�3��e7<@�V9�{\�>-+�߿�,y{�QO���vs�h��=$t�����,�aA$�Dv��'���� )�g�?�Ȑ<��w+�b�=�7�����I2/r$�%�]sw�S� YI���'��/ч�J��6�zDरAq^<=��{�B1�^���֟��瀺�j���ŁD�4␒�ag������L��\$y����4
�	-耼�60�����ݫ�U �.v�T��MP��;�
���:�D, x����Jδqz��V��U5�$����nm��ZS1�g�]x5u�q"|P���͜��_��[��!u��K�t@Շ��z���U6��^~�n��}�u�o?��#��W�n-�C������ �c�@�`��.<��4@� "4=���t<6_*�[6��m�3gD�t���`A�Iڡ�8��i�Y0R�-k����F�m��%1�a�T�:L����`>6<�Ƹ�5J��u�E�u����1]]_u����ae������_'��+��m���I��,�HD�t�C�/t��י`�i�+8ݚ78|\�!�n5b�re���u�/�����;SBɈ��r60s�>�����m��4�����^�:��]�vk�W�>Np��s��]#�i���dfIP�-��	����+�|�~�N$$4E�$�K-��d�3���)x���6��m;}�����7+Nz�ޱF��=�3/[k�j�0�U�<v�_�wH�Y�A�`M�����<2�[���כ��8�h�i����t�8�H��I�ڙU��(n,����e�@��d��h��L�s�����vm��e,��;TD_��>�]�Un��P@�Ǒ@����wl�F� ���2���t�n��X/Z}��#&�d�%M�e�һh/( R�Q�BX5/@��r�9�^HH��N"�p��ܾ�20͏KC�
����y{�[c����D+�����DPّ����-���"&G�>��4�,!�p�N�U,��^a�3]�5R����'%-).�xh����\���:�/��hi��N#�G�(�P�@�� 䊋P�*���$(J�s3�`�ƈ���]"J�c̫	Ɍ¹��3�a�&���}S�JFYq0xD�uUv�>���4�w��KuЖi� b$U����L^���|�y�"����i �<�8��� ֦�^���Ox({����ڈ<��h�$��:tHh+D��oB��U1�G9�|:0~?n�I�[�UB\���N؟%C��`:sU�ꀎ��^.I�{����uXSp��t���d��D���Nm�RCF4�ѝ}��~���S�6ڒA�D뜲���ѵ��T)�'s��J�����*b���)�Z�4�R�~���~��ҷ��O���e��mBꮑin)f�0C�Ϫw��>g)�u�� �m���k�W.�cLp�:o�9�m]�1y���TzWL.K������9���T�h�eJ|�گ��~Xѯ�B�>'��N`��e�+�v�����Q3��@3�D�����&p��o���c��KB π��'|�y_��V=;M��)��k*�R����s
��j��Kv�5��rס	��RDr�
���P��� ?�fv�.ʭn�BEw�^��I��[M�`$m��mU��B�te���\���bqJ�x��
v��;�ƴ��,��a�nW7�y=�-�=�>(��� �C5C���0E&b��Mu�G�ڭ��F���8��5�ƀOvt��	�t�r�ok���4Ff_S������?M`�>�2�p��OV���ݹ��{w���L_�s)e���4�{.DAۘId������+"�
	����͞����9Ĳp�ss&�q��{�8��f��9˾�E��7Qߓ�o� ������܇�?�)~N
0;�v�_������q`�4���'��:��7��f,L�7�Ԭ6�l�=w��*�'�[�SW���t��
<��P�%=5�$C�6�Q�5AT�œ�|�T����`*��o���9F��k��!^s[d�w�z����h�g�C/զ�*�'S��=VȞ]�5�u��.�{�Np#Z{>�G�c��R�^uh[o�%���,AE��i���+����N�^,�)�qh��:��8�]<�>��&X ��ձ˶���Z7��ʍ*���*�k��4��/@�V�{{��	c��32�!2���e��Ti�y�>4r:���LF�%_{8�h�E�܅m�����������91{Ϲq!`y%T)�.b����S`R���Lnx��|�z5�HMmz�y$墼R\/NĔ��n03�c:@���k9�5�"��m<T؄�S��U�WT�6�b˽�qo(���b��d2%uO&Tf��4t�6���@�J|�Ռ4��z)l�V��z&�Ą�1��V����6Z�1��G�tA�U��%�~KM��wH~8�ϝ ��f�*��o��s���=��",���v�bY�A�<��pɕ�8,6��W"�h�!�� g��8�M�-�ы�l
ɡ�,�N�>�U;ӽ#�lˊ1[�j��F�����m�����.��/�s�2w">OM�����z�Ÿ�xEh�>Q��l�k����p�=+,�[a���+�����=�� ���#^8/T�0�?�k���<�.+�C��`9jȓ�J�0��]�`d��X�M忒��ص�>vo�X�<�O0zD�~[:�~s<6*A*gOY�_�KƖj��!ӻ�iQ;f��0Tܳ��Mֵ�,�ݧ�7�*�ܪ����tZ�0Fy�D�9s%'թ���~a��7跮����%�v��I�-�zY�D�ڽ�r��{ЀJ���{z��n.3@p��)8a����aVae�!y{b}���̯NKܓ�qEpLϽ�0���5x"+������zy#s��)K{��$�`����{Q%=�ܘ��2���#\A��P��b!����#�!AB�;�p�%�]O�$�9�b����a5�PF�����H��&N(NH
��d�
�F�gO��MҜ�=�%�f�ǵhل���/]ǜ���t��~�=o,����l���A��v�5}��{|}���ciG�w�
FAI)[�*��@��𸩔��n��Rm��f`'��Z>Gi��O�,?�H;X��UD�R���c\9<-��������3���<:�鳸��٫��6��$����Ȝ��%W(�oȈ�����qw�᫹��流��<9u�N���Ϋ\E�6�!�ip��R�Z[w�f�oMt2mg$Ȉ�?�-��	!�r%13��k������S1|��a����o�����Ĵ�&B��]`k�@�P��OG<}
Y"|}���\(�[�6�B�
���$��"�
��L��Q{g*����z84�u@���q�,a��A���_�*,��W�)���3�L�@�ar*4�\�s��@ޱ���I{��vv[�Sg�Q��`�!�7|wz�h�oVD�`�2e��������S��~to�ր�y9~�|�Ӂ�U�Δ*�"R�l�|K�>����]B<d��e�CX����mS+��ףʭt^��|������#Pƴ��Ռ1�W#�i��P�H5p�e:��r~��IS��\�$H-�fXf~v{�p��L5��@`j���9x	
�e�H�h�27��0j�E�W�����
fy�Ub� ch����B6�@l?Fs�$\��a�"�j�-�<FX� ـ͐Cmoq����q��'><iQ�,���*�`���?-�L0�ڟ�WO}��/5Ne�t��(6�ꑦ"�d��7�N�$�$�s�.P?�=:���` !C;�����S瑱}N�paN�g\�!$��ΞMs���g������:�7�R���6l�E-���?�R��޽6Yy�n-Hɿ�A�YA�z`�熹�\D�����F�j���b�Ӽ%@�@YQ�3��{Z�������,C,1��i��L4�����^e�1�ur�A���	I�4`��L͹X�9��.����s�7ƻ�R���WO��&q�J�c����2�ʚ��������o&���V�C[��ꇉ�eܢ�^˃A)���_�̱T��khyQ�a0�Zͷ3r�|޽*e�lU��.s�h|�*��¨�"��$��)7�B]&��;/��g��li_5����e-N� ��%�t�Fi����)<��B�̕٢䀜���\9��+����Y�l<�<ٛ#?`�� �z=�d�nB㲒���.7v˛�u���:3��C���:�Jv�|^!�}^�*f�M(Zm�<���u��H%�{��]���ycy����s����Hy�	�o2���,�_L��C0��E�K�����0���0��atg����Qg�W�oS�~�8��c���T��kܼZ�L/kFS.�L/%Ǹ~P=���Z?�
�w�{�yҊE���P76?�Ow�YbSBw�9�H�3��@�6a�b������3�Tz	O*�3�݇���z��64IG{C�fW��s�П�(�2�=8-q�7��Y��7O��+Oq�R�G�+�e�Zn#Qs2���?�֪{Nh�;a �s��~n�:.+�WЂ���"�2ٴ��JBY�6�KX%���c7�ϮNt=-�9\ʹ��A��P`�q�f�Rt��)F�|�[��tM����0s����6i4�hkT)&�p�����	��"��hm&ҙs�QrS[�`��(G`��@�?��6������ҥ��u]=����w�M����gf�կ<}}AI(�E���3tp)�G�'�0�!m����H���#��آ��f�������P�a����-�t0֓��A��h�m�j�
K�47Qk�(0I��oT%�1R26����i%����"8��[��(��nOT��Ԛr�@�<�
��f��j�w��|�==8Փ�j�b��(�
0����l���Ғ��=4l).0<�P���c o؀=5W���V4uUg�;���ICYF{8��귻�G+9�A�ö���bX�)�3�K�� ��F��L?�\i���}
�b��ܭ9����vc ���a���
����
�q ��^w��4��xa����Iѿ�N�Z��>w$��70ֺ�LV����#������밨��{0bƙy���a�������"�ܧ�'$a�1d�Pe*��լ��{�޴�E�ņ�:�O���TZK��	�o�?�>��'�<�`ʢ��P��K|�i����d^}��𨮹���ӭR'}Rf`�p�I��xݻ|�����]��EpNDs!�Ǯ$�^=�p�n�����_�a��t�`���4���3����φ�_2!%�^Ұ������)�t*��P�7�x�l�fr(�]%�k3�<ͭ�ZU��g������ɏ��������#������%URX��D�,wm��b#�9q8\�/��"�d!��F�i	�Y���ug[r��Q�$��H�%�@�)&�؄nRe:�G)e��&���e-����;yBP
�&/?�%��*���_����fSC���l�,V_e.��?#xv����z����e��Һ�X��)��Bҝ,�l��,9�P������11)�,��?���(��u_��(��D�ʡ)�#V��~��I݋a�s[z�*h����Fǆ�g�j���v���#zj'5	�/����)u
;�X��O��a���I������E���c��?�PnD/�'�͘ز��c��� v�ˈ;��:��V�~I0~@/��'�K��2��No�����`iK��	n�aD�yq�j%��[��H�ףG<pB�c͑-X��U�=��3@�K���T�8Y�&������!:_������D���W�V��G���)�t�����ꅡW�h�]���̸0+�o��y�Gl�
�܀�Q+؉YE���ؿ�����E1�n�#�I�v3ׄv1����g��u�Ӣ�R��{�2e�(�{ɩ\��`[ ����+��� �%qd�w$b|�;#���|q> "O%y���F�|����ӽ�:'uWSz-L�E�y���k��}��a��A�`;�PĔ���yK�I����몙+A���sMSY�ߕVTxMKgk_��oB�ίy�B-�;j��pWIw|� ��������ޒ�-��-#KJ��l����"��\8m3�����פX��5�D�[�6�9p�l��0ə�WYYl�f�|�����������H@e�>mM�[w+��y�Lv�v��o��4~�s,�� -`W�l�4ض���!5>��J�q��]8�y��w�@��C�k��}��.�6T}{&/w�_�'K��Ӭh���;b��uY�1��kݽ�&��h��HR-I�S��i��*���)�+�H��S�e5q9Y0�1o��&����G��}w�����:%NׁN����: ռW������i�� W��i��`��ߥ��R��*i���־�y�/��J�k���e�F�}����O��ڗ�}_�o|2g�d��D�g�%��v,gh+�,�����.Ei]Rܒ�����6n���1A��x��j�-�v��:�k��Ìj-t8��%Y� �r�uRi?�q��O��x��5�� �zɕ��P��U����5� ����c0&�=d��P�#
rs@-]J���L%���z�x��؞G2�����k�UF�,|�(�j�"w�#��X����:�=c����Ux�s���Y'd���Й̔n屆�gp���|�hZ�(�
=�6q�������e��<
Dm�!4�����#S��r9;��u��A]/�v%�µ}�-��+@#�S���4a��g�b�>R}674_�d�/�oF�� f���=7S<���x����+��:��>�1p|_%m���/H[?��	���<a���sG5A��reв!��N�W���5*V榽i�$���a���6�2qG�3� u=�s�al!��R��ʉ��
�H[�'�e#R�^��|~۾O�����qJ���e��� Ѷ�޺Q
/�!U�:���8�brXt�����*[x�:��6ha�=\���`��AY��7�6/׬�rK:�P��x�1��]ȃ�c`8=�Rz�i�cש�0y�w��1� �,��M�g��*�!��9̣s_"%
0�h� �~���H�Q��RkhU%lq��!W��:�~%cDƿ��4������ǃ�ƣ�0v�#6�SQW�=�Tȴ�F�qvV#E>>U����
�)�܋����;����$5L� �D�r�@?-q�X���<޸��	�ߪ���}�X��2.PU����9U��\MIN�5�ni+G�֮s=m�����Q��^�'����`�	zM蔷>���s��FW���h.X���qw�u�G/�2)�r�$�Tf�x�1�4��9�������#C�û��{�����M�h��Z��u�͜�@vЂ���Lrj�� +�Y��US���S��:��3viXiB���5���n�0�����!}�b�>��"ɕ�e#��T���>�*�XE����Ҡ��O 5��71DX��g��'�N�m%�KK���)�h�=�����be�Φ�z���&'�����ۣ��P#��rBD@H�<�r�c�����ĳ���C�rN��+�]]
�A���?��w�M���D��a���Q�sC63��K�JO���H��R��aa��l��8W��ך?����L[,7���|*�!W*�J�`r-��bt*��E'��3id���
������)?�^�f�n٥�|՗���m�R�u:�;>���}�V�
�m��e�^"@��_�k5�_[�*�K������N��Y��-1�B0ݹw��6��2����8I%���f3���!�ِ���/Hk��np�8�ulq��X~�U��w��|2'�2\�L��0{�@�Hs{���f�{8^,RZP�W�I�:si�k���Mc�(}�A�?��/�+�6���)��מ����ł����R��j��|�s^T2�F,޼��*�� b�]-��@Ύ�)�4]�	?�����v������U$�~=��$zlKMWe����jq����o�������F����:��݂	��#C�¥Ҏ��a���\1�|l$��B-l-��в;�@D;E�����0������o��-�|F���G�qe&0�(�/)���Ӏh�|o�{���h�d[�C/�ʚg����1Tz��P�^��`&�����^!U�.ͬ(k�o��n<V�d4��&���Js斕A�m��H��� ׋8����˹��4�t��V��(������(��&�x�j�T��m��nЂ�e<�g|J
���Qk�+2�t�ֻYR��qߌ�Z�!���(���s�����\H'@�)|��$�51����BT@Ȧ�(ԷA�(_V}v��ʝssr�H��Qx�#F���.�W"���7Z��c��|�؟\�7(MT���3�JʦD@ԃ�p��s*�=��C�
�	.ȀBX7I�Mn�Nȕ�ĭ?tƶ�*��|a�ڼ$�n4���;6Fjo�#�Z�y�HXO���4q�ƌ*��hjl���d ��Q��b]�/�R��1�H�Zs}��0����Hx"Y	J��V9�3��ׄ���fRq"��|;��ϯ�k�W���d���1� �O��K!�a�ԋ��@�e�;E����!��D��&~�Sҵ�kcz�=�ėG��;�>Z��-��\vOh�y����*��)�8h���S9>���q�'��쌸m���}�(�����LA׻�Ϭ-~.�u�S ob.�� � �(y/6�q$��h��+O��㝉�Kl�F�E�%����?�$���C0<w��4>9��m9���J�b!�P��X���Ss��/���I�t�#�RA`�P#����4o��\�dS�|��\�������={z��sybafd<[�� �1m��B ��2x*�H�	K$&�$��t���}8੦�F��)�n�4��`1k#�ӏS6i=�DH�cMr�EY{i�w8҃d�8�+x$�+�6���2��sK��#�g�c�}�G�?��^9�R�	%�Lf}^x0�47��?�'5J�p�:8c���|����6�����6������ǫ�k�V~̆�6�� ���.�F.o���ǻ�d�q�_�<�x����/�^',S����a�Քc�q�j���	�?G�?g���T���u����l�A�{G���6ja�.��n��O��d��a}0tV����;c�R���K���0�=���r�֧����T7T�Sv`F�F7.C��/8��>�ȱ����rb�"w��Y���ܳ�r����VH�-_?��$�̴����޳6CC!�s M������3:0c�A��*�w��~�s��yW�`]F��n� ��O)�$e6���BqwP��ξ���G��m!aJp���<�;-�R(�����-��FW�Ֆc�q{��y�YW,��8tɽ������x�a��GM�8����xR��*q<��W�>�g����/�b�3��j;?\�Ǝt����6����E:IY�W�RWs��N�U���m�?p�(m�0d����k��4���� �ԝ� ���Ǫ�*L;P+��z���V]�����'2�ȅ���5�R�膃B
��'d,��-y����W�9YA53���NU�w4��\b��Q_Y�#'�D�)�kK�L���J8�w��ć����{+�,?+���զ�X��	������^_��8��D�6n��8L�i��&~A7x�:[�������h ˆ�cN����^���]r��V��	�ɉ�u��^5��VךY�t�C~�ji ��*a�%�+n��_hE;���)��{O����/�]�T��;"r��8yx���W�A+�u[����rm�1�QT@%zf�퍈��q5Յ�!�%�½�x��n�k�Wb	�1�e��/2�ij�i$���G`�G��c!���>==3��	e�m�9�F�Sp�x�V�����7��Vt�Up���'p�&��s��b�$H���F�Gak�1ix[��3�k���B�m�n�������In+�s!�{� ��a4�4#�*�q7ҧf���'z����3��8�A�F�ę���'�X�C����n��`Q��9��*����J��W޷&���p��xd��p���k��0�[�3���t��3��X�(h�@>����{}zj��@q2�r��>�e�x>�
�XQ,n�.&�Ef�����	(���3�x�s��61���0+�ޗF����b�D+�|�MSSFE�n��c�ڦ
3�װC�tↀ���	�F�}#e����A�_�D�6q$�����8��[���ʶM��x��cw�aBsnֱ�w�Ae|����EAl�����H��b������J\S���t8��.�0���c}��@3�8�+L8���],�`�}�z�C�gf8�{ 8��)Z��:�f���W�MB ���R���r��4�1�(��&��1l��L�!�gJ^kq�����>]�n�h�X�p��3g�d%~�o%,y%Ky���Rp,�U^��|��smi@�h�!���?�ۨ�t/��d��ܮ/�"��;n��$M�~Q�f	6�D���^�`�W�{������V'J�� �K��J��яi��EM��^"�vL���_*>>��bB
�9���e�y?��nKr^R��߾���P_�1��?�Ï��Ӹ�C0�9�) h�3I�0��lX#�v��NM�D�%Z����tE���@���	7$H	'�pY�Ew���R���z�����P���}��t�<W+
�}�>�
�zP�T�	��}`{��`�9���Ƶֲ0�tnO$��Тf�=������T�Yȵ�T����u�{��cH���1}�w�_���/$W��"��!]Z�#�ַ��p�I2e�ݰ�lXX+B��;�[/=��U�g��������c��
 �w�~��[u��'�9/����F;T�Ԥ�5�F���ӽr�_1��koH�÷o����Q �-X���g�ۙʲ!�"�� �oI?؆&u��I��Ó�n%L�q����+��W��+��4��ϥ� �3F5�[�����sW������Hܸ����p�H��_���9��Es����!���YN�ZdV`5ʹ�M�n�e����Ɍ��o��D��0&������Q,'�'R�,�S�ZU�=@������
Qm��H� �;�t�w�w��_�9:,.hk��[E5�9�[�m2 Yc�k2�'v�n0�����	��7%GK-Q���P«����(���_ο���Zv������e��34o �q�[dna�ݩ뼬xLX'>`��b����t��G���g�������M(\QF�����������v��L*��q'��m�{�r�U�H�t��*�1��(������b�Z2)��@���g(���R�����ӆ�Rh�+ŗ�Ëpp�w77��a<�GҒ�x,� +�,���+�qIA��!�{����e�E־�ʴ�}��IE�͡ �DPs$�����j�
�Tzx5��Z�T�-@��� �U`R�;�Х&0�2�XKPQ=��K�om���G�
x��C5y5�֚EO�j��K^�m�R��Y�.a@Y.�w!�mL���H����I��^D��`������Cu�����TP�}j��2O%��&�q��cA����{*­-���j��*i����K���G� p�Hڈ�*/@�;Nc��ry��U��:�0<��y�i�>��fS�����?���G$ʒ���!u�s:6�����o�M�c�(�XW�lt�2R��1�����������>�s0P�Ʌn����-��	%���DG=L��0��E����@�	���P6,��v&<l1����S@�hn�� �&��q77Q����� %���r~�ge߈���;"s�U��5�D�������Hp��f��D!riL_=�[.%�S;:��&��:�I|?��1ιg��L�"J����9��L��O�������p�Ҿo:��)���`�x�Kf����LێP���OY��/23$�*#��!��XU8��kow5f��]@_y-Z��D��!7g��䉯~�������;J%A�D C$Z��w�,8���N�f�YۿR�od�ਹFX0�
��M�-�~4�*���Z |��a�9.Tl�+1l٧n�2�,�P��m�w��k_�S��&�>�U<���f�����32�����<�����3�O�@;+��l+S��D�J���4c��{��/b�oPB�۲���B%�����-rx���S`J��ؒ�;�r+S�ol08�?�j���w���D�7��
�;+F���@�Ͳ�0��S3]F�����89��[ǹT��-�}�#��
3���$gH�d�)An�-�-�C�o��q����D6w���	j�$z��C�cXe^��}#�6#���s���o�R�{$��ڳ��:��>T;�:�-�t<�y}O]Y����&eFʧ]�#��>��<���Ad�����#��H�*��h[Q��(�h����ٗ����v����6�`�c7�WZD���úr?�\���"��[������B����!�U�"J��c��ct��q�ULb�1n����)uĵ�EM nP��-�����ϸ�T�����u��R�#�o�jc
r,�R3������ n��@�me =���Z���&��2�����z���M~Z���n�hK���\!�-����R!G���v|�}����#�Ǉ>�-[�%��������3����z���z�������C��H �4�����"����2���M�a�P�,׷�~��%�b&�/U$��P�_�L#SS�O�c��-������HZo���R���+�IB7nk㉶xyXt�}�z!QE�$QAYq8_�JT� I�O�j=�}������ڹtj��7���D[U<<cJ,�A�#$eB��RC���f���+dl�f2�W���-\��#źT�E�
��� l�I�;�f�x���o(�I�; ���.�Lb7��y�F����Ct\	��%oь�;�,��A���3�΂�w'�,�e�\Ӷ�ߵ�n;:���U�pև�׵:�<�+X��q�@��v#�<x3����[�&-���J A5,���}���eQP�H6�v61L�b�-/rJ�c
~�
I���H2��3�IJ����y�M7�#~��6"�{��΃���W|���q��XRIb>�����yў�`4�'�^�)������wM�U<L�N���~�턿E���ydwHܸʳ�����N.+��0��}��ț��;崶��8�u�S�֗�<˝�L�ő陬U��ib��� X;��}b����1J�&p����k:yňٿ��Y`�ܵg	Xa {a_�<|�5�6���ku9��X�_�|����i=a\{�2��>N��B�{�����4�9�)�eZ�!k�;,�U�뙉L`��9"�1a��(f����4�_f�8�[o� �� �c��k��BbE���)T�Pe��0�z&���q�?�N~���(���I��3w��`�T�Ю4/,4��(,�N �v��͎��X	@AE�9�S��5c�F����G�@#ͼ .0���jDW�[蕽���	6��Px"$���t{����F ��-�nܲQ�=ۮwR~b������u�G�]( Z)$!vh=mg&��� $V)=�)����ݻ߀���0��&?��{	�ڕ�7�$��"�|�"{J�4�I��p�Nh�*xTh�� ��!<��V.p�P��g�@`:����I�[�7���-�|c��O]�\���N;<n
.Oc@�I���%!n��
;j�y��r;�Å��H7���yqʋ?�8�2�Q�ڒ��X��7D������h�|)��W���x�~4R\�x���C]�.c����21���j7ea����i~Ֆ0]�F9�)�ʯ���;��@� ����y�CNFo��ȴ�Bu�}�G�P��W����y�E��l��Nb�߹�rz�Ίu��j!�Hɴ(#�*@�=��"�r���~�|&
6m[�rN�H����>0KFʈ⫼�Y
�������J�_#�փF�߫���Ưï2��v<���������D6԰�B�}i^��	�i��j���RK��AO�:�f�1��M��E���V+-�-d�\�Fo����OMf�XE\�s�
�O��]Vņ����Y����G��3ƸF��WJ��o��NSe`$8�9�)Lw���u��st�`��V�G����Մ}/Q�?!��v��-|�wR=V�
��|5�ofzBi�jdF�
�qŭ�u�܈������p����s���?o 7�a��,�}\��B��j`�%�.-�I\�x�M%�~�02]V
�6ԫ�2���6�v3t���y���hU���G�t-��.�|T\�% �AΩӵ��\�[�JS�!`!X�8�z����8�m����U|B�k�r�%����$�4���2�~�wQ̎k�<C�^�0�*�\ɕJ��r��"�x+��C�i>������j��_�O�r���v��|����+�i��Dݜ=��~s�����,i��7�Ʈ)@�s�����yd���~�J�����}�D�+�-q��쮤J��|���dMM���;"q���9��?�FDB�� xE�#_K9z;�haV�+��UP�៬p�Z���~2�H;�24�C�p��q�cxo�!]n��m�x5ǫ[|<�s�@9���2__zn��40���l~KH>wEc���d�r�E�=c�zʏ߇�g}."-Cs�v9�Ll�rI�TX�f�'�ۺ��
$�r��Ɩ�Le�b�(K���ƅ����@2s��v�I�����c�(�!t�[��y��qDp��J��8i<����K����2 �����<��B�oaaf��%%h�yj �uu�d�p����7b��0@����;���;��I��k�@�(.B�`_��Y�ⳜY˾��m��`�+���Љ�BV�"[V�l2�*3ish
�:�x�ђ�$���0q���,p����x3����n&`p�:�����Ȝ��zlԷ*��x���{����ϔ�L����ƛ$���_>٘�!�5����KT�*"�;'��(�pfׁKS��vd����PȒv�`6쭆���A�S�d���p��L�9�_����
b*��%�ɀ���~�V$R�ū�x��� 0�����J���|��1�U !�z��Zvr�C
/����и��A:�7O�E����Ųv�*tzc_��@����qD�DXEC��K4�Ҷ�t\ �)J����h�dr�K��	��i���u�|䃈�6'{HX�H�q�S�%�1p��z�3�G$�&��UӘ�hz�t/����{ò���s~���:I[�,r��$��%���e���Z< � qA�`�>������R-�2���&}ÛY���k �_8	�O��SP��b,;�-ܾ|�E���bJSq(L�9B�v�|a�rE��I��z�5��+��I�����e�_��9J�N:���pKy�3�����h���[p
��(�-|sK˓J�4���͚/"I�1P6y�O�V_׿g^�29aM|��~Кe��âj�w.��}'���|,}�N�;o�5B�R�ԁ�.�1�R�-��/I[�j	+�v�;���Ȃ-;c��J�h���ۡB=�_3E'#�}�Y[o
�S�d� jEv�]�Z�C���Eު�raz��c�o�cy�l��t�x N�|{'�5��P�D�^h����O�4YT�:�A��@އ���j�a�e����x�
de�sAw����JF�q:� )5�4y^��Hj*ci"���9b�Nv��P���{[�i*>a/�M8�TO_��w ��n�Q$L�X��{�-}+�����{X�ۭV-�GXd�83("1�,�X���"�Z/Ml�a�>#�UOЧ�����o�n:�B���8I���@-	1�ԍ�l����Z_t��'�:�:�ܳ���~r�ǜʂ���xq�~��&�[���G���6����'�������NjIm�o����lѹ�Á�أ������ws}�=e��epQQ��c����No����9������|��A�n�~�\�S�A�q®ȩr�����|�}[R:`��;�N�Y�a�9��H��9�O�K�{�d�p�?����C��뀺�%׾�l�-�b�����Z�g�g̒eV�?���:���y_T�&��QlAs��Vv=�`�Όv�0e{Û�	hO�P�L�����qH�Z����I�E���6���h�w�&��R�A(�WM���C9w��U��>�����1��7��l�	��������H�KgN�7���F�W��ޣ���e.���Y�m�o��ʑ�f�Aމ�'�����l���}�ԧ�*=��F��~�3J�������"�!Ii2�JyE�F?I�Y�u�%Ԉ&τ��R�Q�Rd��r�)3}F��2m����?5����3�̶�F`->t`�[x�3~������(���X�yτ=�J��~<b�Vc���]"
QR��A����v�ڽ>�'�]���}OY���DM3(�/c��(Lr����7�H��+�@�]���IY���;V6f�;�ɾ��#�v��'�k������-�2��5��oЙ��D�~S�}�U��F�e����x��^0�zG��IB���j[��W��(hƭ�lmtF�T�
��g|�ž~���^a}�2�
�Gk�5Eķ	~���W�l�������1N�B<�JW Ns-4���;l�����;�W�zi��,7��<��(ě��DV�.��S䪁�E�$��y���d����X��4�Z:��,��V�:(�֊~����g�^�x����}��,�	��_��6ݷ�[�u�f"~��l�����Z蝅����4�%�E��
������y3���G:F�`��s���z_�QҾiW^ޭ8s�����|�J���uV}Q�8=�Q�R�r�+�a����ћܼv�a�������^�g�������M�T4�<�5a~F��O=����/f�7���
Y]j�à�Wvx�V��S��ͪ����hsB	�J��/5aYN	��P��M��9��t� ��_�}��5�\Ҵ�/҄�ARŰIc�kb%�8p���
������_�WO/�P<,�Iҿ��55�Bu�!�3�|5h;�d��X�:hL��	*��ë���������Q���b�K_��kHU3�7���.�y���\�N�����J�}m[㝑����03h)�}G ���������2�>��A?P���H_<;$pgvm�?e��V�<8��2�'�T�_yΎ�7pwiI���]thKP�Ne/Ǒ��7�.eU��1��]�쯿�Y
v�JZ�x2P����[�@�L�R����(���Y]2�s=\V�So���z/��I,����uN�b V�d�x��G��E!y��ę��|VWP�t�j�g�{-�ܞ �\}�-c�<ko��s��Ј��ځty_sᾶ{�>�"�1C��\��gگJ��LZ(r�T���i�������!�uee�Ua�>�vfz'�K=�	�\߹!'s4Xv!qe��Y������>O4��=ܙ��X���D,΍r�����q�{���D��`isJ bշQo}3�vd��1
n���gdz7|L����tɮi��g�	L�[�~�����b�o�5�Aԃ�+<1r�K��!����q���D�,���E�����|���G��g�C���ԙ�������4���8�L1^�ѻ��\�}�^��/���´R����.*��"i8K�THQ>���@|˒s{D�fi�LE���L���"�$a���k�e<+?e�5�v����BscX�x���f��&YG�?����:-؄0Uv/@g��]��)����Ģ�}����?ĆI.P%�q��v�٨�c_�Ot$�)��(�|[9O°40`Xϒ�A\#"�[�`�V�/��;ܝ�<{}%����i����1���z��W9m�s���_qɔ�j�$ؒ3![�L�X�0�0H]9�M�h� k��E~7���\�3���A1�)u<� �;����ՙ^��CͿ����iɲĠX����@;���ԩ���F���t� ��	�Eq-u]�4oK<�T�V�48J`t.$K!�>}$�γ^Rp.���z�S��R�]W�5��O�L"B&�(�N�U�8t��t�=��G�'�;m��8�i%λl5�Sj@� j*�g0R�U]e*�/�� xP����:a�����5ߐ=�ru�dv���i��m�_�D(w�� ��>V�-�g7m<b�?�2��뾂C�m-l!�z��tDG�`�U�p<�%�`y�m��g��÷d�i�81i��c�NE[��I���ay��������!a���IEE-L~͒��^U�X8ծ��i�gXy����ָ�h�?{c��葯r&k��RO�u�^Э*�ܽ޹o�1 �OB65Ow��sDX��Լ��� '��o�:�h�4�Wf�/�D�葜�q-0�v�9[k{öL�a��OIzNk:��h<�G����9��3LV�ch
��h�go�CS��n�����s,�f=9��RFA�?s>�c���kA���U���8�ָ[|�l�Zvh\I+/����ԃ4��|�s?�
j�֧h�����]��S��<�i��:T��dg�\���8R��W|w�A�� ��D�M���we���=������Y�l���u|H�TR@�d�|Ӄ~Y�Hv��v��%i��^Vqg;�t�F�+��r�2�jd��ܸ�e
kI�x$^�i�.�D&�kz�z�ױ��àn���A���&�g�������f\�������f�!�,�tc�T�u���3�$0 m�J��mMk��ry�5� wd����Z�@�?�Gˑާk�r&E�l�Z�W48�a��̜��H��]r[��K���x�U!1`�bm��v��̝���Z�+8�mk_���";v&�~}/:l9AC����(�*� u�	:�7^��m8N����4j�%�[��PA̦��`g'�>�9�s����p�nT*[�	�w���m	9ų+Y�@@T�o�K?�S�)�T>��8�>�(#��m^}�w��˭�(�"k;	Z9CŜ��:
<qn,�)I/�0�'�-A,<� j�n#U3^Ѷz��KnF.�Z���r	��1��증�<�f&X�Q�_�2�0ӟ��	ʫ(a-E�T���8�= s5X��_M�arC)�������A�O��۾j���A�I 6�� v���q���k�)otէ#ue�2~R
��q��i�Z���%p {+e[���kݽm�� Ѕ�.����,g�ee�^��-$t�E�M����aUa�Է.�8>;�Uֹ,�-���󎓖$�
�
F�����J�`3���vD��f�@�ؚ^r��n�3>=�a9X�O.�
���r���?LZr�aQ��^�nX�L�n(�WH�M�e+`��9B�U�}+�ۭ�1:����T�0 ��T$|R�"�#��8\Z�3��
�4$�߲�VU����q�Q'ϒ�V�oųc^M���Λ`*!�F����>���S����&�wP��rkY�Gf��g�����{���+�޲���Bc�ި�ÓE�#E���`���[o~8��ج��������{��T(jځ(�D�6�[\��6]>����뉢��ɚ���\��W�a���
L�҂^~1��<W�<�����j��pmd~o脓,�1H���u�m������LVqJ��--a,4�����}��Y�� P-E�(J�+����/n:�V�#
��!f��!��4W=��SJ�:ɺ_��p�s�E�"�J�]��YP/���B�<�n rg n&��E�4�f�f���f{��:z-�D�#�U<�d�Z~�(��30|��=�Nߛ�x��i�2�pP�K^ҿ�˛��+�5b��8F��p���̬�G&Ο�:����Ϣ���1�Z��d|���$�mǺ�o��{��,��-�g��s�s�r:�j���9��� s*Z����{Ё"6G9�x�S�f��V#ms8}��;ᐶ=E�$���d-6��8�P9�Äs�c��ޒ�]|"��ԃKnaװ�ek|#�+�����xǠ�S���Aj���{��Q��hgO�.�1Z�l���2ڲT4"��ɫ��0�=]� %Q#z�0��Z[AC��*�$R�y�s��.w��е������dU�/UNA��^�����A04����?I#Ac�[��I��>uФ�:�&0�]��X=�~����B�D����su���Ks]T���|�֙����(r%�b��x�ۼ�Gf�y�a##Z_�����U�D�/'�  #F���>�]���s�1�r�L0�E���/'V��P�ZVۜ
�̔�rϨ��YO`v��RR�d���D
a�v�!ɴQw��5��q�D�T�xC)���+���-a1Wa�05�kQ9�2Ao�Z��L�N8��˚)GE?��cP��?c��l%�D��ɁG��wB67YOYu�����-�Gp������o*"��I�y=gDL�aݼ��@,]��	����鼸��b��V ��f��������� �.�C�����r �����(U�BUR]#����U0����/� �od�_�����b$� H���V-�fڱ���ErD8SC��p��<ޟa0n�5)ϐ��ګ�i�o���mѿ�z�Avm�'N�#V���(��Y�lF��ǩ�(�F?	%�=R�R��N�Gg�=(��+��*�t1��?(����e3W�[vj�Ҙu�.6�Og�ܝQO�������\Q��P%�C��M&�~�c�������kư���e�|�%!��^O�q�kY��L�mүю7�
��WU�"&� ��v\ŉ�,v�',���~ BƚAx�SVO�_�L\��y�A��}z�����R	ܶ�as_�˞+X�4=,k	�Ԓya̂�H��;�]/W3x~ہ�Q8}��Z��#޾��ҷ=M���`��~ѪL�Z�zU�J�t��CD���;��b�=F��=�t�?��*�,L�^��;%�%Q������^4�l�'qܿ2�����x*����ua��B�!������+��+��p��|![d%W��������$V1��>764�=�q,�M���B��fN[���E��` �f�cc|M��R�<Z1c��֦0Ï���nY�]�[�c��N�<�W���G?F���u�<p]$���'�|Ǫ�8#>�6p��+\�'�h�a	�?>��0y"!G`uE���Pċc��fU����>��^�a4.?l\����!���*�*N�V^:Ơ��m��.���Ŕת7.��"	�y�{���Dv^�#�5�5��g8Rϰ��n�j�	<���L���]��(���B����ѹ�g�c���V��Nł�j.RP���X]��Ah�P��
�~2o_�m":q�+�Q2�[XdH'��.�V���Q�� �x(?uXSUR�s�˰0@���F)E�	��]:������~ag����Ah���-K�5ڼG'��Rg(�;aJDY~Ħ��qo���p���3�;��}y)k����?u񎴧s�]�MW�ҽ���Yf]NĬ:I�y�ϐ
˹"Ϙ0�y<��%Xt��'��As����=m^�ᨯ~ ��V��ǽLs�dz� ��UK{�)��P��mW��Ǳ��':���X��`� 22)�Yvs�sg��dY�E#��ǀP������b#I�ż܉إ��8[�\4�q��Ug7)�t�J��oPxC�yV�3+3��g?ϖ��F��^�/G�ȱƝ!ӂ8x��Ύ������guϖ@�s���Z+���W�4BS6�D0��$4�'%�l�E�����Gbf�?"������~Z�/aD����}�98k�5���!��p�g�e��#>��0�������{a��-������;4����Jk\�؁�X��|<c���/k�zAMT�z:Sғٛߚ��i;.;!��ctu��	W�@�Ԅ��.�Ev�n�^��FP�\���	���z6K-�L�Y|Wt��B�BY�
2d��uH�T/��O�X���E���u����c@�L,���7.+U&���i�g������rA'F�)0=@��d��p�QoG��:�+	��t��i
����^��O�ɱz��~u��x]�uI�[�_B�\�9G��1�k�C�_V�"�}�|d�����[�����:(��1�6������ۢϽvt��aȦ}e��;�쏚�A(�s?W[K
�"�:�jV�G�E���8f�3��f����⧢)���*#�@\��^A"�����Z���j�ɯ�Gm����,}�ǧRiuB�wt��
􈯄/��Ϸ�@����U��L�tv&�-z� �����	��V�?�W��x!qw��ml]K/���-\a���5C���\�f�RhAR��>HV�ع6�Ͼ����AȤ�%�W�� P�w�I3RR���$�}� ����L�>`�p5�$y	�/���G�،���
)"X�qh��uז̞\�	9<X_RQL�M��TF����#��= �k�t���7��ġ�ߔ��f�k&� a8��:���2��Ƈ�Q�����18㬤���Ff+IJ�71Jz�ͱ��<�H\˲�<�4�P��B��4l��{8>سi��?Y��j<[B{����(떊B�\��J��&�$�6Gwq�)��$O4 C��,�b�:X,���L��<.�Fq�x��k��`̠j�m�����
���f<�H)�o��zk��`��C�dX�8���4��)Ȋ��8�W�	�鏖@7is2iC�������cr\k5Y�$^�����b��?K��؛.ҝ���y�2،��Z(��p��A��3�ë϶�H�W�h���l�*k��D`�+qPx��`W�wŤ�A�T�3��m��4��"k�n��>��O���X.;g���w�b�r{�1�o��pH�ֆ��"�
x��Tn�DfV���[��R����)��k�"iu0��8�����r�l]YE�%�8]��sg(x�צ�77�W�p���kF��ꦗ��_��A��R��^�.������I���Zs{�/�PBron)&��,TK��*�E��Gq^�`7����u�ޅ�Q���Ts^6`:����g8��֪������>D�yue���V`21N�c[jO�9��o�2��u?8�&:F�V6FN:J�����A��jcx�f~!q[��$�5I?s�pU1)���	�w@�9g�-�s6C���r�����%b�F,R�p���I�=ݕ��V@�Z����y����A`*���b��8N���iaI	���.�@/Ow���_�*S�����$T��i� [4���"��vs���jz���~��Xs� ��Tx�ru(��9"p?ݣ�שg�P�PM������^F@=��b�U6���79#'��g5w#=$��][@���L)�WC�Gh,|�Zе��� \ώ��(��unnP����	��/y&$(Uy �2E��'.���+���M��6��O��*��}���>C8�d��ӄ��|�����Y��ȩ)���0��w&�hP�c���Zg2L�P샖^��}"K�j{y�������\�Hh�g���YVR�ɢRCU�9/����ɑ�pv%@������
\��H�&�F2,�U%�c
j�ȸ����;��3 �S��DA~T�o�$1Q[�?�Z@�@,����F��WwT3�hB�PS����F4{�כ�����0��HL�C�`�-7�mΜ����>�3�,o���]�#BC�V�M[Wf�7	ْ��I��ז�� q8��y���p;zH����2�u���3i�A�~��[\+�q �M6`(�U|P։����St��ѱ��a�*B9`�X�F"���<"(�o4_j?i�o�r�e�6��!�8ʢØ��B`b�Y�Պ�-'��+0��הG֞�����]X�V����*��qcH�%���u��?��T*ix����jID��_.�0R�j���.�/���,6�;��'��v�;�<��Gt� ,�ҫ.k������F��*�MD�5n�g H�`*��/�>�Ӎ�� ��!_r{.��0��n-^Z����T���5Tc��u�^=-��6�nQt���H`x�Mm���qd�vgl�K��nIBݵ�)���^~O�0@����H�ʃW.��Ex�HM%TI����l��u�S�s�(y���pY�y������r}d��R�Ò�s��)	���Ohж���;�1�"V��F�IEd7���F��+�p�J�ͩ�����Tgl�F�K�\ ͕"�Z(��2��<p��⊢�&� �_�X5���&����[V��y1B{s$r~�F-9�+��Z���[P�x]�%@,�BeT:�ׄŰR��2��u%���|>���V*ːء��̼v��4�-��H-�`b��w@����ս8m�܅w�����O
[rǾΌl�̓ݼ[iݗ�YR��ud�F,����qT�Y�׾4:�\�jw��}x?��OFL�i��9`���`�c����ic��$ɈɘT�S�3��w	K�|�rF1��H�u=o,d�vk��(�c>h��z<�u�o����7�N�|�cD��N��{/+�~T��`-}������nc��bV��5��@�c�B$�]��-ߞ'v�F�*��Eo�SC���6G˔ߦ�!�]O9�M��[�E��q����Xh(�唳�~Sx���zl��q��l�Bk)��{ʤ�Y~�ZX@��2�B��QUvط9|m��7=GZ���6��W��<��LV�Ԍ!H��wB�RJ�34���
�e��n�Lԫh�2���"��E�E��	�7��!K�b��y#��|W��R5:
�M��n�.�����i�I��D�zL���&Rj)N�B�"Q�n{���fa*VQG�
?�Z�F������&��f�����h�Q�6/"M��t(4A�t:���V��;+�Qur~h��?	�nğ�bd�p��\",˪�p43G�g&��6I�!������);��c4t��f2'��ah���<\��B-�%�SC��}~�e���K�zVΖ�4��ma�,�7��n�����	��3ҿ�?��A�7�?f!��#�[x?rE��V���\���� �w�F�c.��l������t
 �L��8yX�gݩ	��%ǹ3�J�7��4���7y���r����yP�R�߾�x�z2hDQZ
C�I�.L��#���(�B�i��/аO��0U)LZ��=`�ͬPܯ�g������������6B���w~����*�����\OJ�nk������"�+�[�Z'U�;�S4�U��[�xu��%,JEZ�Y�-^lo�-)'�&oiϰ�X6���o�zy��r<�M�`3��G�%ͽ�;����j� �;4�N5���3�iBX+E}WSP���x}�|��Z�7+r����[mS9�)���3��)���߲M����LLV��G��N.��d�0H�q�(���qX��pk8��+G4���	x�ΡQ�1�I�(Y̧���xwJv堩/h�<���+� U�⤙��({~�*�UV�� Km��2͟>P݄{G��A��$��aa¹�]:=�t�J�y�Z��^�PU�9��|��յ��jA�[��"?��,� )�������/��M���:ɧp�C��8U~�5ӝ �j�+�g��B�CO������t�v��U)5DKG�&� jӚR�\佡�A�����}�2�,�<0��17*ߩ�pC�Y�����n�V� ����V��׻�	`�w��^�"}D�+�8� ԛm-�2/I���Ȯ5_
Bg�< :�f�8�5\�ɋ[TP��#����?v��i� ��g������[��(�B帕�����h��O9��;AJ����9�F�f�GVL�\�ąɣ��EC1��4C`�y�)+���Yx�>%k�c��T�7�Hl�f|Y5eѪ2E��ox�q�v+^������6߸"�	DyB��I���.��h8bWQ�1|�	֕#��������-�z,�P��9�,:c���W��8� U�宔� �!\��	t��L؄s��Kí�:��߹�C�n�y��} ��@ �˗i��/j�:�2��tW˦̼��X�R�<od�#��39/�t�%��|/���Ů��n]4�.�>�7f���v$�z�����������8L�r� ��0�镁������C>sH�80��eu��3��K���������9dtL?������eI���F5�i?��_�&�����j�H.4U��4�G���C�k�3^�=���m���X.O� FQ��qȝ��N��Jos�S�PQ�^�����6��4H�+�KJ�'��_�(��h\��?��Lf���v֣���/JQ?6GC�Rf|��]=�$~,Spld�h4�?ؠ��J	�2tP�!694�P��G��J����4SDͳ8�m����=B%��DV�������M�I�^����y/��0U1�XL������<��2E�a��iж�GHl��Iu�t"G�zk�Wg+>�UY�Y#�V��L���K��?�	C|[.w�]�[eZ��_ �&�
i^	�dD��*�<�e3Q,��P֏�8��C�'C�/��`��zo%�[�K�M��vd��	�W��<<k3ID9UQ��rS�����Y�.V��O�C�u�8�T��F߫Ҭ�}����F&�]G�V?n��҇	���B΋��|�� ��̞�,������0e��i����}`2��^��D�[*xsl��v��g�$�H�sV��f'![}��&׮	�wF$�{eK��ڵ�Ə���Ɇ�����WX��m�v�!E�I�c`n�V�~:�����+�A�J�������+Eϗi���枛�u��c���}�>�����KG��6�r&~�МZ��<7���wu������6k����ģ2�	��ukY[�wk���Є�ŎM���b/q�u0��c�w��r���{l��%�?AG��G�"���e���J�D��eF�;��\##����*tO��t�q�xA�Ӧ���pxR_�3����q|f��������Ț��i.��i��>k�";K�$�6��>����������<���-�dv$H����ھ[��d8X�=�8�d�%�i�Z�+�#�q9�@��~rSه�����+�YF��c���c�;��Y�b��	�#Q�/S�6鞙����A��Ñ�>��V��Tg�d��}u���0.
M{d�3��E{z��[����:����cM�)�q�2�؈AZ�^j����������.GD���#���I�a�Z��D�o�a��=BO�迊3M�7?�z ȡ�tde��5��f=Uݕ!/(#�7o��V�]Z�t�LU,�h쥼z]y0m�������]Xn#����u1OI�m9u�Q�U�`>��s渉$2�PY�W����+�!ݜ�'����ߍ���mq�d�]��;hf�=j{���ay�{�������"�e��ɇڬ�|�2�&g!왿]��ص;��D������X��g�t��9+A��=K�Y�/�����ls������ɔ)C�X��}U��!\���{���9tɏ��?�Q�v��kjE�(�j�d#H��*`�>ED�g�q����@ˬ�)��@V���m�S��oT��_[c���]����o8�~YT DBd��4�:��a�L�l���2
����<�U8}oX�����AK��H�f���� 0'������lZ!��٪���	J�b6q|Os2.�!�����FXm�ۺ�����{�Z=]����k5c�G�"^d��>���.�h�A@�2�$�I9F�����_G�hi�(�����AN�v8q����wt��qK��W[u�/��]Dּ�m�.���jY)�H�c��
b:�r���Sꫥ�nU��Hx��D�t�̿���K
�y8�2HM��
�`�M��g<MO�����x;�s�����}�g��N�u�C�&�)q��W.C�2:�7�	�����^L�fO�����]�!� �X(��![�a�鐚
��b�%Ӱ�\f�q��򬂳i����b_�7��,r��J�����"
j����E�"2���S��6Qŵ� B��t�f��
@��ϸL���L�2L9>�&Y��(~h��̆dw��e�ةŋŮl3���ӅCp��r$LT���rU1��8xi�fދ�Dޤ��I'0�>�s�<��c�<]��r�a1�7���Ŷ��F
�[�r*���NJF~�{�ǳ�W��.��d��X�R�k�tˍ��ӼP��ȻY�3�'��L�$鱹�,>h��|Vj�w�s���R��/���P]���D}l�T�N[�u�(>�x�:E}�H�=��O~�|���H�̿�.E�|���A�� 9ǩ� �;��3%���Ü�D)��Ng�T8�f��FS6מN���:(�$�#�!���x=��Y��!=hP�5y���.��gy�"5=B�I,�D���,���) ��:\������/1�9����	6�d�*�� |�֬��밅a��B�J֖�/�ӯ�7����Q����
e�~�w��v8��![��F�'��ϖ]���cE56X�%�����\ϫ{J�8o�R)g�} ��@�����W�(�Kx��0�I؃�$�zR�\Ra�b7� ����������'B��Yt�Cj�Rq�[V��K��Ȥ�LY���w'�:�(��)�������㪘 �RgV=ˣ�V]�"��uJ��!&*��DGC=� ��ʚ~�I��lblT9�[��DP��Ry�n�!R5Y�;�R�3 �Q-�"��<�r�P����:�S�Cn�ؑ��Ҏ�.���R��&z��A"<䣒ph��i;�NG�Y���>�`��բEb};�,�r	��iB�7�Q�Ķ&a�� ���p��c�BC@����?�mjZ�����4c�H.���@/1��E;���A����1Z�ʀ�'dv�d1���#̏}2��sp��#����O�5|��SB��^>��g��SU�yi�W��K��>iF�ఱ�5��L��^�2n+V��9���	��Q�s��$g`��m)[oi�1`-۩#�]4�)k���@���������A�f<t��^����V��q�-��M&���O�O���R�&�i`��0�{�$I�H�f�5	+=��ͷ�r3k�Ҿ�.X^pt+�Q����9\F��_����<�4M����젞�V�Kl�p��kxp�!(���_*�uˡ�jRe�����-���Q�qs�|F�Š�پVMC�As�(Sۡ��?�*.;5)F��Jgd�O5W-o8U�rǹs=A$�ߑL�(�d5�h%Գ�w�DY���M;į��q�ǢH�a������G���[v�(��u��'��&y:^ȴ�HD��Cd<͚�Wf���)m��_w��G���'�+12Mw��caR����Y!#ǽD�%F���������$T���8Nsg88��򦚛U���w����!��-g0q�Q�ڱ�]mse>�H�L�/��}&�?��ԭ��Rlz�p�~�)}/�h��������!=�~�*���Z؃05σO�걩���դ�Y{\>���]B���-�e5�y\��1�Wv�)��Ϝw�z�4t���(����EC�M�'��8���� f?À#���5��¿� M�����&ɾ������J��P���9;0}羲$��n����Կ������>��q��5>%���W�NM�F���s,7�т|�A�9A�Frj���Vg��$R_hd�FŸ��x�/�,#T�{� ��]-�>c�ۄ�����݄!�ET&bi��2��d��:��p�91�������\��P�6�&D����fL�j�kYZ����p��{�T0=���_�� 32VyG�Z���I�~�+o8Rq�5�N�U�O���rG������eݫ�;��OSQH�rL��m1�9��I�5�/�Ё����<�h��� �g��8W�'z�����R�7�kE����`t7����ېEd�yms���H-����l�|D�\jtJ4o���qOI�_xs�F�,VAo8�\3��;e-�FB�8htX'�����%�ƴ����1&]�T�sr119�!�9~�A�P��&Ǒ��We�BM�h��"5ĕW0�c��Z�"</D�
���Z��\�����F��mK�R�FX�ߔ���s���^��!�����]�*�� 5��՝
��|(C���.9Vm����9�*+�^2T��`���7�Y��qp[ᠯ)^顱��o��K��JB�I#>��j�>�G �*>ðd����'Z���ᝑލ�vBzLG��ϕ�z[O��CnJ7/Ώ$|>�ېQB��jz�	�~4�KYІ�����x#ۆ�1��/��?��Z�ϩ�5�ŀ1�L���[�(h�W���4-�HyaI<o�f���R"^
�aV��G�^�ߔBے#u������=�ȵ��I+v`OHڰ���֑:���s��5��}����F����>_�S3%�b��+ܼ�5�y���ߞ�
��f�G�����9Z��TKb�״}����\����8�7lV�=����L����P�x�r�r����g}0 �"&@6��ё,j���m1�|��0�$��� k*�����\�\��E)5�:*�v����k��2��!���̚x�A.�/��X�i�A 0��ZV�v��&�z�pwpͿà��b��3��L��A+�y��Ԙ��&^`�&���b|�K[l�/v�J�iK�_��m��H�3�vq��"V��p����W�w�#{Z��]o2do�J���l��M�$m��y^
�.T��䟌 �������~���$�X&�ϫrC�4��J�ݘ�X(�:_�_���w�'*�<���-q`���)I!�6���x v�B[\zA�d�B���tP-����;�/rK+��$�������[�v	���i�/͇*�{�d j=n�{��wu���K.����t�b1�P%�0f �k��x�fpN_�U����8���c�3���XeL����V���cϔ	�;?����4/��l�;�1=V��Y7�N��F�����y��`�%`��I�h⮩��R,�-��U�U�`�j7Дde����J������m'j�ǒ6���4}�(��
��h�Kd �G�ʏ��)	ъ-����`��R���"�ʹ�p�q�Y�m���DAt�@��F���8��j	A:�G�A�ݵ�Q�/TR.�L� ��͉�Ԡ�(�at��Q�'������0e��>�8Ի-7"�Lf!)o�3��G�&[n�nhl�z��Bٌ�_�Ϸ����򆆢�����.��#�ll_Zd'���b��������i��W�@�]J�C݄�/�,��+�)^�}л�n�n�?6@%T�փN��n�|-�I��n2���Ή�`m�*�6�d�"~��g)��Rm�a@y��Ը�:�-�Q�zv�_�$n�1xx�t��3,�>)�~��sǫ-�����t����g��9��Y^��1O���H�M��a9��wY�=Gy�d	��ₖB/�EI�p�9��n�WQWǩ肆�l��ǡ�y�J��K��4���]Er��$^*�ժ���@�,
�u�iҀId���d���K��r��F��Ҭ���v�np��#ͳ���e��������\�c�AƐ��#�^���;���bş����r2��S�.	ܕ�#JIB���?��z��w����@-0����,�n!����$iH��:.�oJm#�K��8y�Z�v��mBH<�:��>�wEt��*zȋ���((��?k�,��``�R������^w�D� �*6RW�pҟo���w����R� �d��!����2��������If�zgEap�D���R1W��=��d���@��lC���N%z��!83�	�����5���O�D��ʈ�#vR�n�e��؉?�_T��6����3�l�fy|+�����.��4rg �P���?�2���I�@��}~կjS��I$�SDE��#q�C�lQ�v�fLݣ
�0��01#N�&-7��l���{ߩ���ٻ�\l�NB�&��'����F^gƟ��)�GXz4��9���܎�v�#�LOh���`�Z�IL~$<��"k�yx���վ	��oj��'�/�>/7�:ˑ����[��i��*�1K��Z���I���
�\w�X.2*���Et�h_�P� �)瘢[�pGG�aJ�/h݃��M��i,�u���7�;>N�Ż�=�FI��E��Y�-pɳ�e�r*P����f��V�f)0B�Wĺa~NG��E�1;+"�a�1u|���9,`�(�J~���:&s
����@���������RI�HD��
�K�6L{�����C5���.$e�dn\�8�!��s	
Y��2�D���
u{u�oz�a��F�]���ॻ��@хܐ����-m�}��i�&|��	@�r��;*�r�N���W\Cir���K`kXm׷�Ѫ��}�!�3\t	��
�
g5���L��}�G�g7׉�!���0Ӣ���w���ۮ�����Ί�!�K���t�<�lR�>�"����՛L�l	 ��[T����3C�T�D-a���d{OCC8�u�S�� �{�PR�<Ӟ��|���k�	@�t�,'/�u�X�w�b_"�Z�Rd�LH	rG��nR&e�$OqG@��}X��R_�N	ݳ��'�r4�d �B���~}��u����a�o��`��,*���/���|W4�� 4\:�H��H�7�S��Jn��m����K^�w���C�rἈ���S�U�GAN��Ǐ$���p��Na{�Q]+GJ��QaR4�7�*�٧N9�j!�鵯�A����7t�*�v��	��s��8٦����1|/�+�����S��q�.?c��P��3Q����'�OR�P�`���#� �'H�4�w�RJ�,n"�ϐR"Y��i��܉�Gyw:�8�����I%��]?[WeE�X�� �{��m$���~��`
�^�jN�u�n��[m7P��!���b�/!*e�����U5Q�2^�\W����@{����(O�Pw�#>�8�9>*���1��S�}`��
}� _Z�.�5�K��0$�Z��ޚ�G瑊o U�7�@�kT�"I��Wk��3�+� '�C���	?f�W����[#�y�>��ZY������f��e@3�f$�	��#���	�<Թ�Ksˣ��ht�k���C���XBƓҦ�(����~����^���u ����E�:
���B����x�O7�hَ�X�Z��f̲�ى�Au\����;�c ��>�^E/$�\ܞ����[a�6�V�]�]�>��t�AT����O(+D�JIχ��B��}������u��}i�\���PR�K+-#s4���]>�nH�)PU�ZpH��U9E���f��I��e�w�מp_��/E4F����[<�=��H1)c�:�2<�����͇a�u<��̓[~�|�0���78�}k?��g!�F��O��b��h�_�ͷ���Sj��T+���A��󫇻�4�g2!�,�bLd�G>P�1-���<pqf�H1�G���
��ܞrf��3�:���V=E����W�|/������kw��b�CQ
`��^Xspa�+��f9�@�r�Aj�Z+��5�ʓ�mٿ�%�%a!;j��햩\�G)]]�ӥJ��P��Y�L����ָ��ߥ�5	U_"��F%S��}�F�Ϡio]<�I��q��ZET)O1�<����ܗ�������%�*�6K~�:��1X<[�������c|1����~��/( 5��mc��!YW��:����`"�С��tQ�<���(r�0m�#&��:_�XQ�)a6���=woꭽ)=o�5��|lF�dp�D׀�۵G����P8i��xM����x�ç��4ti<q�i��� �#L�o��0�R!A�P��J��?*��n�r��iR�{k���p���
�'���|]���?%���+~
Al��V� >.	�$b�L�2A��@�/^���y���[������3�^�C-��g�F"a�0A������h�$�V�8�FC��
�9"�?{v&���@g��C����n��]+��DRP��`�H�o��y�[/��Ƚ�*q�!�3����V\�3N\}'�{�*�"��#�6B`+WR�P�y���[��'"�L�h�]};�*.��p^e;�l]ȴ�����}�$��UC[�7�iw0pcy���/�ݤ!��-&P�^�ћK�k���i<�m��<��g�vml�Z`�N����w9��!�,���wx5�^�͇0�5;I�0���'��2������S�Z.o��]?��ʐ`�_l����jF͠[w�Udw=�6���0T��T�:aR��޽����::�m7s@�^Yiu.�����z k�`���\W��Cvc�P�<��vH�=�@aH�	AT~����cz��^g�+��
����2:����ϔ�a��'������`��]������)�ȁ��U��&���}���}�Znf��&� �K10��a@ �!=�c�fm[-�q����Q�N���?(�,|6gms��<f��<t���V��r����Zϯk��4�!`>��.|�vg,W�O�:���>E�-6^kr�e��y�Bp�p��^rQa�D�QXf�Z���9%����F�1�%]��4�Dgм<��ȥۧ�["��L��U* �KG�v��q�&��*'\{߄,�������6�FR����'m��;�&R&A����R2�P�xJ��O⟱�(�b*�8S�.s��_D(��x�F�uNɬa@U��k�9H\(���>�Pِ��:��9���O���h�Z٨��.�,sɋ�i$>.@�u�ꪘ%�KN!��O+��9���(l�͔7�jArlv�qՔ�al-{l%
�v�})�`��Du@�U-V�|'���O)�4�������(O��о��7��ui'�sMC��"'����ޣ��F���	c�n���$~�Yе�4�r�'e��4e��k;�I`�Ni���@���<�^'�E�� I'Q� :6���;��OO?�v�=���?d�ZAr���ha'4 ���@g��_O������I����5x ���M��&6�#:/�����1"��{.S�Ҁ��8��AO5��2�u|�*�+.��>�8�B�Zj��
�b���Ʋ�OVO1��&E���eu����YQɢ~&��3�@�f[�R�>��$���c[�mz~�i���"4��Π0Q�R�[	�;��[Ą�|�`�u��[��݂��� �#���~� jt>:��Cc��p���)�L�7�a�ގ�!%Gc�=��/X2�bŷ����f�4+�N�A'�0�Kg���>5�9zq�H�'d�����ߪ�,�I#���#k�1J�_����q�T��o�ϳ�@�!�;��
�5sB���:)��}�4PU���G�v���m(=��+���� ��syVfm��B�<�U_˨h\{z��4*�q���I-�Bcgt���_V���?�m��urr��
��k��ۈ��� �x7��@�zv��iK�1"�W(5E;�v�Å�kUA�ҞrT���F��I_H�4M��OT*�zxϚC�(-��oo����'���Ĳ�g�la.��Y�/I�UG���Dn�W�̐�#C���~s�����3唏�y.n�/�B�d0s��$�&:1\؉�=����� �
��;�շ<?�@� Go+㟏x/j��}ѧ�m��ۭ����/��^%���5����ms{�t��Q�<t���\Z����6�X]E/�]�a��y֪~��n�{#��{0`�8i�~+�~Nңs�  W	�y�Ӿ�<�Ķ�I��a��͍�z->#�1���Av7O���05M�������]��sO��ȇ��([��z��%"�,L�18�B$Ü�
3 �4a��!/���0�X��d�9k�c���p��nߕ�~�'�����dz����G�$Y�R��E[�TV�T��~|�,x�I�;rp���uVs�(��=���\*u~9$?y
;_(ެ<���g��Bĸ,��x����� '�8Z��t�x�k*���v/��A�c�q�Kx������ͪATh:��|�"��z�kL����,�������
���u�,�芌yཪ��f�-Ν�(�e�I�x[c���ll]��b��]��c~� �s���>7����bcJ,�v�+���S�g�u�q���W2�&��6����cy��F1��:A= ����J�6d8�����1[�?�s >�y��N�D�J|q�Tdf��|���������5�����=������X~����G�R܀ T�'��!PQ0��3D�e:S��ׂ�q�?7Th�Y�x PY-q���$9��QDE�!�c~����Z���w��^]D3�5w�^)��*�IՋ���%ܩ\ʨ��>\�~���E��q�˞F
z4�I� .eB�K�X�S���ʀhG����\z0 I�|[�����!�*�W�%rA�8!�F����D��ß�W���l�$Ce��G��0) =��GO���^�	��a�KHn��f7'�9�����#qz�9Ze�����5��)�ONn��5��������e�<��*5�Qc��ی��S�:�K�D
�\Β������
4�3s�O <������E�O��[�~V�]�3솄�-?[g�>�z�&[�
C�F�����;[�"��Ɨ�:��%C�y'�3N�_�v{V���ߨ���G����_��X��w�.�l#U�g�*�J�`3+��X�+�K)�:�o�\�� �X!�Q���s�L�K�p`��i귶�Y�%��U�H�NL��.,V/���Db���ɋ�L~kfy����۳��ԉ6ݼeߓ9�$v�e���Q�f�E�-غ7&����g`�%�nm��D���zL��7֠����M��C�w���$o�S_Ш��[!jx�xuK�yctR�p8�a���R�FͰ���Z�F��l����>L*�񇹟��y8����>O ܥ7cw���T��ғ!i@	jߋԢ.g�in��~�`s�L��O�Z��������Q'o�R%�G�bE�ީ�����Ȭ�E�Z��K��[x��w�����a����y��:jR�K�y�7��������x��|W�����D�+?�2�ՆMV},:T�/��Xp�7Ζ�M���qn.j1X���t}E��(�h�,WY��/9/�J8@��:��a=���AN�e,�Q�ѹ�,C�����"�؄�B*Ź����g4��˺L����ņ��e�醭��Y�yț��{n��g��,-PC���:&�c�Ӿ)��q9��R�����8�(��7���*�h�ѩ�������*+Os \����ڒ��j���ڑ�Pc����f��H�z>1��a�	Y�B��?�9��*l����Y3�'7�K`;7.d�2T[ �s�k����I 6���5�+	Zxo%*���-q5p�h`�S���!��ο9~�D�(Jۻ>������v�͵ʕ6d�N<0㖤����rz?y�+����b��>�+��d!�B���+�)^u1'��L��,<i����ND��v0�K���-Ĉ~-?l���f����mЁQ�A�M��a1���7�[��+�6��2�[#]Hbl�t�F�����R���w�� Ӈ�@�I����s�W\q���&�H���h|)	KfhRخ���/�	�A��z)l���f�W���r����?B�C0?u��U�I)c��>��;k�Yg�h$�s��%����լ�:?���I��y�we�WR��@�v�\��<�t�����n��Y����.6!�d=Be�m(�I�>E�5k\I��a�{���c�a�!!F�nora����kr|ec8㓑�'w��� ��{睪4�I1m����湲mf�)���:w�v�#~�)l��7�r�;{z�����Z��bߚ�26�Z� �,R��63e���2,�����[�������][o�+�G��iZ{L�{�J���l>�g�D�7AO�Xa����(�!�?	��I7`%sd����;��ŋ�6(X���k���c��^���
��Ի���o��aЃ�H�Y*Yy����澆����ٲ���4M��ؘ6�G�A���C��
KmW�2�9�P�_�gЗ^���]uk��.p�Ahl'B���Ú=Q_/#)ɥ�_s�d�ŇjЉ��Ճy�������������r"b.�k�G�%����eU��h�ƅLr �����mā���TL!���3c@��
g��,O[�.W+yC�~d�zI:�O�u�8p�O��ѱ'����Ͽ�L�8�*��z�=o�4�Kc�3i����m�2�և+�L��}hO�V��d��
|"����EyAє�+Q�����H.6D���lM�<�� ��p8�+�b]�((ӚKJ5"�A��]%���㤁��k���h��F����yKZ�&�z����Q�͆;E��8��2���5|�7�m*o ���Z"Ğ~K�:sۇ�n�q�I��K�<��4NEϔ�͘Wqik��%&.mо��O��Ml`ϖ�Fn�9��\OeEsfn���/.tG)Dk�o���`}B<�(��~ @�N?�L�F�=:z�?�W���Df�;�P];�d��.�������Z��0��nK���"B�d=pYN��^֧��)�y�����3����N�j٦��X�J�r����6��y��?A14f!F9`����|VmR���>5eZKۯlZ�"Ť |g'|j.�ɉtΚ"���kCd�	!�J?�C�\.��/�l�׺o�.0��o5�<=�h?m�Sva�4HU�mC�v��$_$��~��@mw������Qff�ߗA=�Ͼ�i����~���͉Ʊ��}A�e�^ E��� A���
�W�b	�ZQ���>�Z8c�'V�
[�<B|&j�J �F���f�� ���?7�^	�֠l6�����Å[�)sx��"z�����1W`Р�')�5,�\E��y���lW�[�[��J>A{�I��W�ei]�Vʉr�}�Cn' :0ZIE��yB��_W4�0�ީ5F����M+m��]:b�>8�#&�W������eD4�7��'h��U4�B =	�ٖ�勌}�|~>����G
�OE��"yhB���F?X��Q��e����T��������e��`��kc�N�hV	`<>�;�V,M���p�ä&a�j������)��=y����%��Yi��v T<�Qd�?�ۏ(����'	Ö���^��[��v"�}�~Fդ`D�����f!A�U��~Hf&g��I�<{�u�=J��>�8�׈g}�i�R�����CN扮��R��Qua��� "5�6����Ym]d�b�i��Z���X-˩�W���1M�+��ܻ��W�? �k� ^JA����u�o�jk���'�85P�Ά
���x[u��rK0��>\�ھ�Y%o6?���.w*ppsR�{5��=~�T�GFz�n�M� ���
�<�:���I�qυ�N���sb&����;|���(�wnz�'��K]:��{��cS�H!+�%�TyM�f�v[�^cA�(=��{ڎ�+t�US�k?�� "��VAG]�k�TBKB�bB�����;_�F�>)/!Aa��� ,b앓賱�0��[���9l�������
��BH�P��������j4Zi{���hv�QA�u7�ݔ[z�s	�H�͎3�`���od}���2��q���TeӴ�n��~S�3���|���%�44���X��FC��ȡ
�"��Us�X�*����7��޶����Ik��*��S�_)�]��`2���$Ik��?�>� �\+"3%���*l�Q�� �?����j�e����x�܅�ы0��]�PtP�!�p��U�'/oӖ�y��m�a�_Y���X����XY�m�vɎ�I&Qx~��օoW ټމ���=���s�O䟋8��N��t�7�c>�1�k�eڥ�M��N)���8K�ד�&GU��܇Oc'�nP/�Ĵ���5Z���q��t�����FG�7��w'Tf��*V�Y�B資�@˸ɧ۟}���5+e�޺��~(�����e���&%U��GF�'�C��:��DiH�5��maydS�K�	�T�X�O�I���	4W���EmF+�d�{Tt~&/mT,/�b����}��9g�ߪ=G���ݦ���g�e�}��VyZ}�?����S�z˅7)4c������"��%"�7����.E�k@�\��y*ț�Dϵ��kJ���fމ/�9�=X�DE��\�l�� ��K�dp�����ou���������^��"Hn�4p���cc�n�,[e�eM՛	Kb2�b�t ��dE0�o����TY$F�F|0}��+�`n�[솤�"9�:V��a{�r���;=��czh���~<~�RkC:h��Cr�Y���Q'h�����j�$5�jR�.Z�MRZ!I�Lt��kZ���M�d�
�~]��j�-�*M�fY��jP��e$7(�}��x�p~�pn��#X�_g=�������������#�o�+˒�mR�Qe�Cx�3J��2�)�M�&��k��պ=y[xa�<C	���]a��@���!f���ڋ�=%��?�u�F�2�c�W3���l�KM��7q�GD��p\�wJ��ߋ�?��5[�d��S-���P�J�����޲bW�6�p/=����_6���3q쾵�o�Z���ւ�s�04�8A���[}$��̠����!>�3���E)a�vS_��<ҕ�zkhe���+&�@F�|��*g
��Iɧt7�!�QX";���<ܽ����C!CM�Az���z3�!sq�w��b��2��
�G&��uq�Z�V�}xبW��{�l�(y5�g�e�D�vl6}A�Z�dK�#`�Y[�-*�5<-�����w�����cL'�����3s��1>�(yJu�"!�^W�³�A�P�a��t�"�s�Y��,��GJ��*���?۴�f�gĹ��si���,�h�{	O�G�~T�Wl¦�#�b�ڣ]����rT#,�!�cZ�Fש�&����#�n������!�훴.��Ɇ���t����U�l-��x�8�9FbNYz�;����0vOU�*�a������?po}��Z��9ف�	cF��Ոj�P^�c�cL���gW7�g���p��=�=�M�˖��2PeQG������ߵ��o�bV�0;/��;�MYWaF���a`Y�ju0��2�[nA��V�:���^�xH�����,�n��U�]S`4�Q�ퟞ���^v�Vy�9IB5�h�#�F��	�1j��ʬ����9���SD�C����}�5uF��P�.�+c������&(��էv@�p^���%�?����C6"�?m7��:_X�\kh%W.��r�KARi�ֿw�t�˹��gmB���mי�!i����$��~��>����?J�ބ_�Y��ÔJ��8~��սl��8�lɛ����u�$H^�ްee�Jh1rr�����Xʟ]o�b��U9<�
��O������9�~��,�B���R +�^̜Nl�5� ׍��e�F��篟�%��pϑC�n�0�9݉��n�uF�]���XQ`�b�L��sJ|�;��z�Wg^L���O��px!���9�/�N5]�Y��T` a.߉c���5`|�S�����\�]gw'��i���[��/��L������H� �*Z������>'�0F�*u��Z��J��
]��Uq Tf�N�<�ug��{�$���	��ˤ5s�8KFb�u]��������R)K:�	z��-����f�Xi@=XN!֊L�L_�̢��p��#���b�ȧy�i��]h��GyCj+ٵe���TE+ŗ)��)K�	�Gҿ:��y�����T�9$�0h�Iq���S`),��E�ց�t[�u�+@�ݮPGW�oQ�Ne��/��A�"g��q���u�U��}��T�/� ��ᅤ7�&��vO��6��^d#%��U�2�{[E 8m�v�+m��AWbP��'�Ё�Y�wm���g|O�9 ;�%���>�G��3�ԇ�Lγ���xL�� ����]R���{~9=�~Wpd��0F\���*����E�����$/�v����<�mα�z��Jo��y%�ğ+���)���GJ�3�/��>���r��'��&C�&L!�戣%Hs,r�&���ј��ʆ��M�?1�V�(��bH�%}�e�g�'9$�3>OT~���'�졙������J�gKV�h�#g<� ��\���"������ĵ�l�#fׂ`Z�s!_���q�y�$%}�9�+Ӛ3��撩���+|���=��=?Wc���}&y�3�ǭ�j �_�[�k�R����楝������x�2���ȂD�ic#iئ�1�"}��j%�徛8� y�~���p�YKss+�,mv~NN�JCz;q;���EF��������*�3+(���1�;��owDIctp<�ȅ�&��u�~�r�J3���U��G\�Kv�Lb��\��U���c��
�uЭ6�v��  B��B^�U��=
$F�ZB�G�����)v%��e�i�&]c�$�����j3��He�b��^oX��A}�Z$�8���/K�'�.H�����Jbt����)�f�0]\��q��24�օ!-pڔ�H�ewHkƍ�v1N{�[i�v+/�=�Ɯ���U-�7*U��˾@���i���J����iH��1�l�N!��:t��8wd�?�����#��C,̵�m(�9�Z�|o�Y�t��ѡu95o����0G��zGމ���s�g�jL��%�6t%m,Prה���y1�otw��@�q�$�#wg'�c3�@�,�L�	J4t��vФ�n�e�����e#�$�+C]m���ێB���G��&�hb�;k�O{���+~;���$�l���S{����)3T/���	�t�gܖl-$����xt
�n�:wvHSF���_C���^"��,2�a*���4��ٻk��v��q��AT�ճ:��@�lF��8�(�~Hh�-�;V��|��@�����jk3vHp�������%g^+R�1�ګ��0��k�h�����p����i�}�"����&���V^���%����m"KY�]�ʕ�#�jP]��1����?dGt�;d�)�|`���7DQ7nW�ϔw���d}Dm��aD�7�2A�ݕd|ܭ g~t|#�o�F��b���Nc�h/]�m|-]C�t��l\�g���:��6s�^-k�1����s�C(��V�&>�CA��
<8�����oeW��h{����~d�Daa\Y�pV!���r�����V����ơ�u�KT�?NaNп;�=V��w'Hd����G1m:(�G���K�s A�V�:��:d�ZLx�SY�[�rK�֣^՛B�a��8g�Ǵ8����X?�P�pR`&�AJ{��]Sw�O(�S~"�=�ƛ���^�o1���Z�~<qҕ��c�q�;����mΡ�y�O��n��a[b�j	'@b��B*��4*�Zm6���RH�q\�,�}�D�������" �����gga��M�d|ԳF&��� �s����`l�������n�F�p�����҉�'uկ*J���|��d	Q�a?:�QC��<��=mAlu�=�*ׁ�k��8#=f�3��ahX{<�j�.��-f2I�(�o�k�b.w��@�<-;�_;`b*�؈5���E�VO��^A��'�#ł�4����YyL�5	��+�Ǌ�2���5$�����v�!k+�c�(g,��
T L�ѡ�D�,j��f28��y��v ^Ay��KDb�~��͋�y�ʔrǉ���=��V��P�2}ah� &�&�K�5��'��C�I�H���
L����~���|���^���=�\��(ZB ���f)��2����� �i�룙�)&A�Ge�b!�z��c �@�=��lL9���}�Yt�}�<Ej�p�_{���C�!��r�j_�����3=$@�W#$�`o�/�_4� t�������q�HC�=��e��Y�*��/���%FQ&Fu�TwO�_/�^��<��1<֐�Քf�e��_I�?`�$�'%�y���H���k1���O��T}�5O�g+{VZ�})-s,��';��0���t ҟ�Z�o��v-�-�>F��P��ΰ]�h+�|`T��zb�>�� �aj�"����u�G��*�AE�%TZ; ��\:�1<��������5ܑh��!�Z�iz�M�bBI�妋Ly�X
~��� ��r�����N�� s��������Pv��k���ƿ��!�����"�50j7�J��hN��q����JP���||�f�f%b ��]��!�wRD�PT��rY�s�f�o1�ޅ!��58�]�=��n	Y�O@>YLq&z�.���IݸZ.0�z��>Ps��E�� IGz^�Բ���Lܓ�q[�j�3�o+[�4��t)��jE�C�F�oQ��������'g�X�'�bA�
�t�@O
Ȏ-6PM�F�%���x�d �M�X�� |��T�K�FC���1��FH�`|�ޖ���U��CND��<e�g�x���O�)���Vp�vi+��I���Ֆ�)Ԣ���@�DRHv<'���Y�G�y��AQ�[���|�5���|dk���� We጖?�o�簙��O�=7
�AQ�s����!���s�~ts��1�2���B�e3_�U�0��|�X�WC��%������t(��0;{�l�&gXXٓ��������ſ�p�����kλ�H��;�|)��� ��kw��/A:q���-"tG���A�(������%�4�Ɂ���}�-�>ڷC�n�EVB`5�J�$���!7\��YHP��F��J6E����H��S�����_B
��S�[E��8[}��{Q��:��Ēd��*剋xb�p^���}�0wS8��(H8R��gÐ`}*WR֕�#��*���p�L���Ԅ�#��>�<������~��+j=�Y[���y0RwL�חM�-<��;�0�|��z���;�]N�\���a���œT=B~�I��d��	0Z��t_	8�p����<���O��+��������㭸�Az@��]Q�E�&C�P3��8;��6k�6h^�D�%�+��+�*½/\S=n��n��vo���'��c%H�.z�`������D�@5ȝ��;O��������������[i�����E�%k%L6��7�6�r9����ZD.M�K�xN��a�p�x@�	.b����Kq �g7��O_�p�ӫ�`��p�L�y(%Õo�G���E��^=[_Lj���4�'2�f�Xٛ�����CHʡ,|Q�:_�h���<ݴ�<L
��g�d�]ɸG	Ϣ�w����^�i ��aU鎕
�*�<�;��8 �D���E�q�^�� q�1q��u��5\r��8�v��k
+�����Y�8������y􈾙L���̂��N������*��^1�1���z5�Ǘ�jbĴpH��=~ ��l�^%��0o�Β�Y��hQH1y���j�������YY�9'������2c��sw���M�|D.�U㜀��lE9�*#ߢ>� )τk�|�[j�{�Mg�I7$�1�H��](��?Y�mz7g%��������wd�}�6D:��	�=�����a>3�������V���рra�QY� 7�Tߡ�	Yd���dD=9= ��Y��\j> �� ���>O�{��{�Rl���??���^�ԏ:�q��Ǵ!�]����Sa�~����wl�V����(ax�Qk&iM?��)6Z��zn����=� �5�"����<[�G��i�`oi�U�C�B�����,8��qR���m'�h�3BQ�A�g;#�ݐ(� |���SG�%���N}݌�� �h�e��nqi�����(�F����n��K���jN,y�m�bt��<�c��Ϗn45��R{0��h@ C�<�v�l��֊�����2C=g&$1���<�鼗W�I�=�Q��o	r[1��HOk�N��#^٭]gD�m��^�).�0��6!���C���l��*��
NT���᫊���+l��`�o_� oQ�uG}f�֔���/cf.//=�5�V��c�|�1����4Ay��N�	B8�&���rn��I�SwP|�!e��Kdim�5q?X���q�>�A���K*���X�5
�>'�5�n��?8{ZC&%� ��K!��i��GРМ��} 
>���^_@�sc}�v]=�X"řX�C8N�W�ZI�ԩ;6�0�[��Ә�-�欇�	&(M������|.+/�-��h�cO�i�:Sv�i}P��B���>"$���>$�����^N���b��8ap�>���q'qe�$?�O��Q1��AAr�^��D;��+(�@��6cW4�%0!��.����A!��3����W��U��L ��D�p+�y,9F'a��.|Va(/$M��iêVu[��\��X��eya��L���?{��AI �	���ӠY�{b;}t��F�YN/��7|M��� ��L��\�abg�������{��lt/� �l�U��_c%�����k���Q���vKl��ט,3�D llhJ�?�	r�^㕗W�؎��B�+�ێr�K۴u�q$��4�jj��+:��{�>#�ut�L֧X��MY��,~̕�l_aW�S���)�'�x6 ��(k���:J�ı�CA@�D�0��L���[��M�>6�0�����ɐ�$\&�*�0���,89L��[mAD��ļc�uwj��ZQ���=m��'Պ�2�s+�` �k8*����_ ��Ž�9��纰c{�r���r!΂��y�?
S�����q[s�aA�E��jp��>y��o�n��p�������2I}u3p]�>�2͛�w�0�Ъx��O�෥~�"(�'Г���.�y���۳��O��@�6Hѕ=Č=q�o·4s�`ԟ�	���\Kpx����s=È��C�9��IQ�#�镀�텦`]T#G��$~O�r��X?T����,wy5ӗ5��n��#k>�vPH��7���Qc�.[�v!?�_�	yWD���%>�>�i�Ϊ[��T�eS��k�--�/X�#>�FwT2�z@���g��`��}��K>O��p�M�T3��]�ǞF<��{�b
5%ʠ�i���΢�:�>���{��R��I�,�taw��=�{�/OS���%ؑƆ��	�!x�k�&�p���S�@���:�#C����,�h��n��H1�H�F/����8{%�lȓ�3����\�)T��zz��/B9 ���W���E��mt/D�;ۆ�ǹ��"k���)�k&�T��mW�	s<pƚ�#�*�U<���%�g�,z�{��?~}DQ �T����0���";.g��/��k|?,:��2�A0Z;��C	/�&�Q<V��1��V�f����*��y�b��U�� ��Q\MYй�0<����}����v�J�j�o������dy�y2�I�I���=	3��S��dMhF{�6�+Oۭ_f�V�8(���po��Z�q�W_`�l����<����~��$/�\��:8\���}��-��?a��;燥N��� @�UYk�o���I�@gN�Y8g���7ȿvo y>�D���&o���5���Ҭ@��Бл7"�P�R�LpT�+�sC2���^(���N�R���JoZ%�AE�w�Ұ�*;=ܧk�ѻ�L�Bq���ʤ628L�kF��K�S�1���>�	�xT�}�Npض���帗 8��,�2\�59�7yę?�T� ��� >� �p�0�x}�%}vN�L��. �s��R4�n�B.j�)���+�m07�:�iĮ����9	w|��EL���_�00%TT��הIL���J��Wl�_�?)8eI�`T�`ζ��F�����T��c�+ G u��c�i�O,|9�b 6��(*5��2���q3�c�4i�m���n�����o���FO����ϒ�{U�<�=�S���s����1��3��
��K��f�Z��ȿQ�r�e#�1k�;��	�:05Z�Z�jk����;��pҍdAY2�t��AL�9 �~��D�����n3Sq)��3�dj�4J�7��pz��W;�&���Т�L�*y�N� Z�%�W�~k�G��`y7�k��$�W����`���i��U����e���8�`����+>p�X������}�����UG>O�Eb5��R	V:x�w�7�[z�С'����k�#�(�-F�I*�L�c���5�#����t�mE{�]��Ā���h'��K���F�e��5x������Mބ�����,`��L?����ci�HL}�����q_��U��6 p�����
�5rK�C���}�^��4)����� �44�Ǝ�-�2;?Ş�*	S��Ú�
�ky�2�P���?1��9���E�I�٪-��v��=� �8 �|�6ak�$�S9����,ppݧ=�����r\Ep
C	�
m����@��oMw�K���V��gO�v�dC@��>�e��5�1� ��p$�R�'�?*0���h���0����9!�a�}PPbt�N���ِ�婴>X~�~�g�kA]��q�o&��9e�ְ�?��v暍R�kd�r&ND�w&��d�&�FO��g��xp���+|�E�+�Cl��Y[�v���mQ���x�����+�)F�lhj��q
H� �J�wފ�P�dJ�ڥۺJ��'rMnw�k�>��X}������n3q���Ig��v�馴��l]�4G>�Ӊ�2�O�Z���qg=������1�*���'�" S�S6�ӭ�|��*j-I�q��MJ��ͤ�4�Пu��ۀi!L�LA�9�\9��οP�|��W����;#��#q%�"���oT�Cu��K��h�����&`3"�cI�-aPW
�4��8.����2��,\�5�i(�z�+�ƚ�R���B�'_��o+Xj��+#F���₶��;�6]��G�e\��寇a��S��yf�������=��v�X���.�w4&%۪��7׼�]��޿�/ 6	���(\����?@�������u&��G 2��,����ɺ�a�k��ذ�YE�����wLfW�y .:�P�t�w��A��'���C���7���ܔ��ߦZ�T �N�/��{�>A��>�,�pg�����ҡ=H'p�Y7�l{ ��?�b\����,ە��� {�J�P�Q����替���H-C��o|��*�>�GIO�NI8ԥ�N���𾏡�����0�=m|�ue��n�`VHDg�
�����e�e�ҁT˜OQ9���;a��6u��n�li�jÀuczw*��`�__�k�&A䯞��:��k�_�2؀����;?�[mip�~�Lm;����}@�>����M�K��K0����t�4B#�Eꏘh���Մ�B �³�C�NX�Q�O)�js*e�2v6@�yJ��/a�ɘ3�����'=�O���rҶ?L[�lX�@rOn�u�z���IAm�̏ ��K1�ھ�X�ׅ0_�8f퓞G���P�����` �()��]/�����CN�����ع[H�����ᓼ��9�oS+�q��6�"3M�h(ͅ�)0���3��H�JU��ov.�2K�c��n	�ȧn�be]������~�گ��[2G�ɔHt$n�u�z)Rw;J��'nCP������^@����%
�V�eK�hgb��]e��К֏���W!?`��{�Tg�y���dE��5	t+��,a��ơ�3�h���@�7:��9����{>������q��D?-^�f5���Z �y������z�]�a[�_�A������!&����-�Ǜ��"�E�~t.��;���b����t�L&lmٳ.92+�րh���Փϲ��0B�/���c�#I��B,�<��ӺU��p\��G��1ӡ���<�>¤�E�0���>���{���X�	�=��@PN�qn��'{�ClR�:�Y���:iٻ���9�� j0+>����g��ei�-�j?Hd~�%׌��g:X�P+ �3r����h��
���w"���Z{��qQ�dY�z�V������Ͱ\9�Xdަ-|{�
�d������S�s�I�\rݑB�(RF��$��T�{���W%b�@�_�v�@�8�g����C_���[�)Ӛl2�P�ݼ�F����0�jcL���Y6�D�-_2+�xRq��H��Us�4�azi�7������Vh�Ѡ��,��@פ�E��{ߚ���A	��1��HyJ�q��E��`Kb
���� ���!��������������kT���ڌ%�N���x�/�K~�Q�A��cE'gN�R���4��P�.�5��8���.&���:��(��s������r0��G�S��j��.�C�`'�@-p�oB�r�3�~l[��@p�xr硜FL��*sb�
��nɅ��j��4�/C��Ô�ȁ��a���0u9nQ���v �ƃi�[���-�����p�����XI>T��<f���ϻ$��~A@�J�?]�g��Ugw�/���wR�D��3iG��qF-�6ȍC�ǇS!�dv�>7�O�$�����c,��}P�0���+��_�s���_�A����g���
�>M��d  �5B3cJ^�����]�W��F&���vb��(�e2��-
&��}H4-�I�:��^)�ˠ��藉ly��&�V)x�ɰ���;�"{BIgc8��"`��o����ĥzgZ���R�h/ĳg=5��=�o:�i��>x,�+�2�Q{��-"�'������(���2}�$�Z�s��w��A����,�'M+U9�\��3���r�vt����[jv�7Բ_����G?$Ty� A�J���s�-L�6��J:ܰ�fdLxֶ�u*їʘm7�H�	ݑM;
�=�g��0|����2o�&P2�t��v�bw^�a��q0�z�%��d�C� �E*ܠ叽����E�`cb/e��H��$_����H�Mltr^9�o�}��c��#B��v6jx88��6�*�*�I�jJix�9�b������|��`��K����֢Z��^�N�:M�M�C4�'�vc��&�[��E33ro�͕`Jp�&1����`X�5$�e$"��䠯`��>���҅� ��%��j 	�d��[ߤ�v�uϤ�,V�������v���?�Q��{@�4����dl�V����7x��U�ѣ����yoL`����]��f�}�������K����1�D�}���ːw��?rW؊�pC8�����)��9_��c�H�D킴M�A<�8ǹ� ʓ�K��68����#<���~Vx�X�X$��1���0R��}�'���cqcǰ�#L�&�'X`2ʋ�"ZQ�[�vhV6#L`���P��x�V��}��^S9RK���v���b2z�F~x��nw@<pG�ɚ�_�*���g�C�6]�:֟�o��h
�j�C���f����2nY3Ss9���or(O`*p1u�?w�+���on�kX��^��b�"��PP´*��ǿ6i��?�\�,@CuF5J��S�}�X��{%<�W&�Y�)�{��gjY�A��Z�Q&���ȭ�����C[�����i������k�����|zs��{?�R����4/V!��?��턵�ȇ��Zs�_G����>?�q�nCW��Q��nX����3K�4� ��s���[�fٵĪS��
E�n`/��k���k��l���#�=ƕډ�e�t#�(	Y#��D��akF\�+	�[}��|�M?M�>��������(n���U��T��i(���|C-9�D<���ƞ�o�k��Q߅���$bEɊWDa�u���E$�":�$�*,�H��B��CrZ)�)�#����mS���e	���V�G������:�`��i�6Wc�c����QW¹���b�e��{�-�Q'�IoK����w�f�ء4^��M�4�V� ��Qp�$<yUSAR���J��Μ��^��,cn/�%g��r�~��0��	�Gx�w�N�����7�����㙒�`I�|��J�����-���狯^ՑN�.O�����%��M�K��{�b%<��˞�!Ә9r��B�3l��ƶ�>��<h��߽U�#�O|Ҡ
��jW�='�s,�$��f��o���^�=RE g6�ݧ7ݕ_��ϩ~Ě�dА�uw]r�����b&*���[�@�:�T���|�	K_�;(�Dۂ���p:�E������V<JDMX
��;�ˣ팃����'J�aB/�+���!H=%�V%�-�8�Wܘ�[E���PY���?�ḫIN{���	�t?8%+��av��G܇�v*l�~!�IY�p�
Lbtv�D.�Y�=�sh"��$C��6�i����w��V �_�t�w�j~jք��:���)9�ҳ�k��à��WI�����sqg÷b��?]ME��s�u�l���;F]���w�B�� ����������!����v�4rg���s#m8�U�O�ee�sӚ~��h����R�Α!CZX���=1�nK4��D���.	����x��ݲX:�D[4�a�t�asX�Om0;*B��;^|�j����d����	���hP-@
�Ȁ�`$?�̳Y��/B2��C�r�@il��7�f �x����]��NP\��s��X�E^H���3�e�h:
�ۀ��k��H����YFR�%�;�m�0�i �7(?��a���x�@�B���d��ՙ6������녯T*���@�p��>)�1g
U�K10����"���eڃ{X?�b�ژ�!}c����}��Ha.Nvx\��0�d9wb��;W��������츏�����\o7e��H����dBf8)�s�,�n��ϳ7-�ЦW�O�n �z��:��1�����b$���2�|��ӏ�Z���8I��qi8ҭG�JV�ͮ.�ƞC.Yמ��'���r����"O���}Z�l�\jN�	��w�菚=8���ޗ���ؗ�,1��ԱRX���&���3Ŕ��
�A�3�6z�)���uOn���ib�b+�:�	�k`)�9?����c�n�LV��g�탼!�y���{�͟�[�?ј����h�q��~���g;����D:��7�o��PV	�Hm��~.�k[�y��rS�s$�j�M�Ұ���&H��q��yvC�RyՏ7g<��g��� �@�-�� $��xPYJ{
�r~��