��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0������x3&3�����h�|*�9�bJ�����7�I�l�w�j�B�x�;x�&��9+���v*o�Z�	V	_�a���:��UL������h�w%&��b�S��?����9c���|��B���qX 3TRnCP�e���e�6в�f�Q�N�#/b'�Mr�,N��ō�p��yk�xV��&bdڿ<R�e�&k��ϑnu�)�ϱ=@512�ܔJoZ�(\j���k�y;=��%]�]��ݥ��^�~�ۨ����8�/�f�N��)k��Y���2D�e������xˀ�;�9�y�<\�`���.���l{�pt��3"��z~>�Q"��M9��."à�̾�O4182-Q�����e��58j��X��UϮ2�+M����6��T���
*N�OE��ޅ��1���Gѿ��m���`�\���M��p�*���*oW���f_w���'ȝ�����kbh��eL�i.�PdX{�K���|��[�4g��/Dg���.lv��F"�F��/�V�w5S�^'9T�3��A����(�g(��ï��JvZ��x����b`O
K�$��6.�d���Y��I;�\��_�� �>�~�!bc� �i��	�c6��H���U���g�$�WIH�O���g�&*5�wַ��s����˗�����}�c��W�F��I����`����W��/�j��ɐ3��L��N9?vj��
�qz�י綒�%��T��23D���֗\�4�zGx�(Ox�����|[4�{(�����Y�d&�<o� >ڷ�IV�x��!zdAG��HNi�p�����PAN��(��!������B��Qj_|��4ك��Y�T�놐\����ՠ�(W�R����5}_R۴�����F�\R!o�)?"0O����ʠ�'�uv�D	w�����f4 ��=��ű��d�N۸����F��j��Eҷ=pg�	rnBp�@7����2�hNNK,@�x��o���55,X��P9ⶺ�IX(�a���Q�6�sES�1��D�C!�(�ǋ�!�6�1ݖ�-��񝎒4��_jw+0n�i�1�r�s�f?�C���h"�;AO�Xw��V�`)ԋ�k���귵Ef���!�*rb��`�?ta���;F���n���O~f�b)���"�I5�q�J��2�y��X����.�
|"E�-TR����q/����V�?��^���N�2)%{��\������fQ�R	mMk�_���~�����C��s����pkJ}B��jƚ�ē�#�@r;~��E�gW�n�f��.�� �~�B�?��]a��)æW��7��>C��2�)iJ��V��)١ô%ӵ�H��:����X9ZFOG��mK3�);��[,��cd{#���S��:�np �����RH}ÀV?���@�Y�[v,Õ�����	��r���E�{P~:�S�ǆƝ���� ļ06`�7\��>��x'u.�@�(���p�O1KZ+�6ƀ�F�H�����z�������ZƮl:+Jm��d�'#�!����n�_�θ��o���ԓJ�h��j���%z�`}�c���b��B�t�;�c�=��11�D�H(�d�OZ�5:ՍU2���{0�DE ���D~&��>�neQ�Vb�؄E����b���+��� ��P/,�.ʵ�7D$�[q`��&�h�y�Y�J@tI�k�NT�0�Q��V��KbP[>b|�)�Q6h���6�i�������4�HV(ϭo���E�,�Ў�U�^�Ω�$�K6����c-F+�{��UǼ�gi9
|����z�i�F�g�\޻h<[�)-Ts_5�`Xձ�Zn�
.��`"������2:�b�G6��I��_u���	͆E��܌�}�D�x���X��G�v�C�F{<r?M�lث �4=�����Y �g��lYR��\|��]�Ý��Q��6�A]g�#�N����8��
�-��#��yT�p�ߣI(���5Zg���S�_���Wp�n̛��������H�1v�p���Ŋ[��a���*�I��Mc��Ӻ��Aժr�R���H8�*���}+�"%��7���r[�5��S����g��@d6�mGNi*��e�|����N�J(O�&3����*���x�4}b+�B�H�{ݴ�Y�-�[(�d&~�wq�-�2��I���M��J1�<��[�����&�X���HϘÁ3�<E�Pm�����G!���k���?Ż��tތ'�b~��mռp����O�c��������.�5x$h)�+�}�#�m^[�=\+�֘$_~�wXJ}-��F�t"��XV��!V3_����0��Zn��5�RzCe}^)ċ� c���7�rr&��{ -�N�h�u��I�����˓t(��75//̹e�bX(�Z��}ȩTۘ ��+�d�'��w������^.+����Yڷ��K����/I�� �P�p�@����"���{h�`�[^x��~��$P���UGK1�W�(�h������g�}����x�B�]�L_��lK�2��)\=�i7r7�G�F,��-�d� ��y��ФԨH�٣a�k��mk�\��
�l�o/�0�ݧ�LAM�Z��e�İ��<�gS �W�~��`��X�:��l:@
G֫��Ĝ��яu��9��y�ΧX���S�b����6�oH@�׷���o��Q��	���lZP�E��Y����.�S��ZUKMQl���.¸Ԗ��F!��������O�#��?a����f�f���)��������W���sr�ߵ�k�+��`c������~Z�t7q]�����4!zi���1cNQ�`��<VR$�G�HZ��;&0w};nR����z1�hx�yYFyF��;)��L��\)e��d�
��p������VqR�r���e��ZT���F���E'x/����w='���Zd�L~�~%����~�ᚒG�5(��4�,}�M
�i������$�a�x6��v��"9�kFߗk��"mn�Rpi*5����$�?Ib��Ζs�Z�:'�g-���R�S�>�bn����M�ݨ�,��X��Y�G�S�(�y��&�`���9���@�^�G���ԅQ�? a�/"[7���f��bR�iC�	F�t�9R�������5���Z�<��bYc#0���N���w��4�}�����2os�Ly.��LY����$���Z2�j�=�D��-�oJtOZE���|Ȭ12�!��g ���CrQ[��3MR�$4cw���i܍r&��vY�YִcN�O�����Vk�����\b1��a���mJ~�o	¯<j~�O��.��������J���,��B�j�gX)�Z$�������h*m�A��3�MB��&18��!}"D��6'� ���NpsݦP����!�u��_C�5�4�8�ug\R���d&~B�{�q<�
Da�����985���wGi��V���R!�9��n��o<3p����3�:�d�C��o�`�D����?��F_��ҍM�\vjta 1X���[^�G���{UrH�ZyG���}�ф1���K?2����"���D���ˉ���t�n����'��ve`���s� jO�F&/[k�~B}LZ1���p6u(F2o}�wp���X���,T���H~_�����uZr��i�\�ŮiT����{���Pf������
M%F��r�݌�8׫7�ҩ&�d��6��-�ht�� M�F3���w�w� }h���K�|��9��FEJ��EY<"��n菾�.M� ��n�][�`'3{X(��z�j�w������2`�MU�=�8s�6�{]<��B-T����o�M��zح�������(Oo���dئr`
��v� �T8�H�q����b<���,4�D��9�SX �4Em�{H���ޗ�%�L��I}Y�9�D��}���D4���-��U��C��{##�n�}�?��ab���"$���ފ~ <�>�]"�G��@y_�>�4bEF�q
�GLq;��w���~:O�HIW�F�- )d��˦U|���!/Βtv;!�w�ƾ1������U���%�a�{�t��E�f��H=7���G ��F)�T��}��r��M��1�Au?�n���C���3Y	<9�ED-��ۓ��T��d]�a�aB�p)�;�j{<��0T���uM����&p�6���;��o�2J;=s����*)�T�}�`�`�q�s?<�("S+,S�:wsL��[�Y7�ˀ�� e��Щ[��lQ�_'Y~9��'�B���A����ܖ�t�]�w��|��P��axXP�����V�����߰")��ݗx����}�_�]��������d�tDS�,����)�sK���ً��um�̚��'�0ᆍ[O ������R!_��,�����r5�!:�wD��Hxo��^#�K)F�xG'��S�	xȢ6�@L���1����Ĥ�2�*I{�6���Ԭ��ή��Q>]ҹJ�;��d90L�W�zxm���pА���:tS� }�������}[@���� j�5"��Fo��ƀ��֨��f���x�q,�!�I�' 4,�v�lV�$T,���8���	"3��/R�Ǜ0�P���]�
��<p|�:���I,"Z�F~Aj��T���@�@�|"�X1���>��0�΂H��IT�Z�@�8���m9	]u-m�*��ƌi���\����'��^-�{ٶ��`*�`��R;�q!Uz�,������v��M%m���qbk`���Z���؞< ~{�S}n�	Fi��$G��ѐ�u��ǆ��Jϱ�ܷ�50-P�z0�� ��W�{!�t�����|�z�W�����"���nWVr��#`�{A�U��H���N�"u���׻���`ܓ'׎�����ּ��%N~j}9��q3;�v�F��M�p���jo�x��s:R�ѐ&�/�Δ5���:NR�%�w>��d8�}��R��H��?�L�suP5,�Ӣ� a=>�oQkQ���!��g7u�BϽ�N@�H��@n`���'̈�uW�C���=�(+�א��6�IC���J;�C����I_c�x��9>K-�R<�1��`h\�xX`D:�ǖ���h�%�o���ѡ��zQ�}Vί�P�3�ф��i1Jq�J���J�g�ɦ�y����qcmƜ~j�Q����tp�_����/����O>89j
��g^�=�M��{���J/*��q\-���͋EK���z�L����m�����Ո#E��y
cL�:	�*�n1^�DFw������ږ.Q������՗�M��h*А�t��@2�S@���π@�@�iS�"����sM0	�X��L]��p�j�}�Ԭ�������^ԇ��T��+YV�a�'���)-������*��/�����~x=���Qũ��1��Z,TuCh+Ȑ�,��{6r�I�����n
}�Bj+k�s Cf=Jd�������U��[��P��n���6�Pnk�?3�o��l��t���l��u�x�d-�fUc�-p�=i%\"�^:j�1��[�򞩭��wo�б��)g��*N�%��m�L�P��YjUBRe2rV���w�[|��N�%Ŗ+��%�JCRm��6����얳�HkHs��t P��y��Ӹjs��A�����1K\��]�p��l �@݅�WO�G�{�:�%�N#[�ʗ'���%�W�36�ᛌ����7�0���2�o�g��XU�2k�٩�>j��霴
�)�A���B�ܻ�lL�݅(�/��s�B�8��f�0lK�r����3��'E�`���L��6�{�Q�l5� Q�RI��g*�h����{.7�g��WP��P����t{�lq�Ӎ���!�2K&�O�/��f�*19�8�h��PR�lŸ0�1u��@�<Zq45)�lgߋ0T�Aײ�t~���`��9��M�	��j5����g�F�Ίw��v�lu�v�����J�9��������i`0��ȏBd)�uJ�~Q��*�B�������sݷ�2B���v%E��_�`fUpF�'ť��@�k�s��ۻO9�f*��q ��Kɘ�qS���z̆@���J܈i�Μɻ����P4�Z}����������y��nd)���R��w���p���L�gQa h��'�̄/�/�lM��*Jn2u��qI$.q!����G�H���M�\ğ��y�Zr
A�Pg�?	��Ϊg�T��ux_�i��"�5�$��G�FzI�%9ʹX�z'���>Y��o���h��I��w*��A�{�Ϻ!n�6әce�W�S��&��� ��Q=	;�%*�o�������$��HǾ8�X0܋ zF�آQB��-�ƕ \���#���B5�*�Fd��4�ڤ�o+��ͱ4�����Y�H�@[�i�!x+���ǇԼ��Z������߀��]]��ۦKa;�5�rU�����u�����<'X���&�����0l�ð&��g��"<��0K��אL4I1�;Fx�y�M��7�� 2�D��$Go�F�NׂFz�}�ua���W$�uĊ�Z��{�N�f�\V���N�؈BFI�8I޴�wRH�=g�p"���KwԒ)�)��>���{�؝vϪ �"��.�{�U'x�hZ��~�)T�4;��rӇ$��������Wl�Xl?�wuYWf�R꧆�Ͼ�.
Y�fK��oo
���x��@��ՠs�%����/N�Az�b��s�����-S��U-�{��6�&_�'�[e��,��X�r�`D��_4� �����n�>9��&�3B�1]?u�u��p	Up(�p�Z[��C5X���'��J�rR 6i�-F@�&�x���`��=�Q�I�P};@���~�������s�G�{����(�b���}Mn���Z�WG�2-u8dD�)�W�ږf����^�k3�3���^uoM��=������(삓��W��S~2QZ�[h�E ��,<~zP��\��FYJ��jV���/W|�OL
�W��@�� kh�\�I5�r��I5	.��t�����&I��=5v:�S�]�9�*[3���<�S��S��
a4�R�~��S
P���n�K��CL(�Gȥ�{+3���i0Y�ϷP�Z��D.��K�ֱָ���2��.&�SՒ�����n��)�a�u[��>	S�+i���ٍ����y�\�<}�J-���%��+s��G5=zݵ �vT��rډϯ�,�
D/{I��a	s���hjm������pz �Wz��P61�p��ДQJ1~z���HU��ְu�}hIڊ�qBn�3g����S�x�T/AZ*�(�.O��䃛�#ģ�0�ii�D�O.$o+�:�괩�$5���g+��9�2Fν�΢M�5C�G-�{�M������:��7����H�ܫ�l:8��r���8�'��ڊ�%�Tߣ���k�[�5<����B_�04SӉߡ�mC	�^(w\���s��s�:��^��M])_ޮi��4�y��ݺ��f�
�ZOj5K��"�M�J8/�7�*�LPM�@׸2����~ўR]l<�d2o�S�(����"�a�Ĵ3a�"r&2,|T������QǸ��[�!I@���f5���Np��Pm��v��? l��p4/Ͽ��#E5��Gb3�����/��D�>�y��\�W*�]�|���n�{K����w�B�n�R�k�ja��/zL;+�s�^ôl<ƴ�uuG�x�$��oF�\�eCgD���vr~f��������ĢX�`Q��Eڅ����+%], �G����b�5���$��ld9f�d�.�p#���V�͂�� �]�_-��T�h�z�\P.��'e7pK��!��F�{�d����W��k��{��ŝ�0�h�<p�ܥ�V��?�/b�) <��\|��~EF�5~��������U	�����X��:L�{��c������e�4�?�������uB����?�e�zY>��v�jp��������))BF��&�����k3i4	C�vdXx�V��S�~ ӂX;�V��Օn��j�������2<h���cK&�Zfsr�fAHk���3�/�rd;C��8τ��T���y���F|�C�%~���o,��6E�f �q�f���Ց�6S~?� �娥Y��i�M���M7��h[�вJ&/�VV9f]P�ϣ�C��8`�Or$��w@f@A��W��a�%��)��r�;��+��{�,�C��T���乐�\��`�o��b�SMK(z��R���"o�aqP�p��k�D�r@�5l�g��%��땷�)�W$� $	e�Ö�	`̂�(҃W�W�E�lbY�|=���rc��!�Q���6�e���~��ײ!UP�-8uTT��Ϋ��z���
�>rva`J)��|���+oK�U���z�/��O_bIa��{C���>��d�v�&a8lt������Á����{'Vr��G�����[ �)��n3z��2�{ce�(X���b`7�Ig5�A��ms�	@FB�7@�?w����㫒�qLp��a��K��`���dbs��`�m�{\Tr���jD6Ϲ�i��i��zq�'8S3m 6JR|�_<��:���"�$J�s༜@�#[�a�Ob	�����}���.L,�I<-�9<L��ݢ'�X.)<�vMh�g �}��|;����!�7թ����ed*�N�s���n���� =��®��Ffj�SjV��̵�A)�%s�;�cXrw^m}����K�l�Uװ7�(��f�û�f��s����y�ܛ�Żi/-M��d������Z�}|���_���mmg����[���s^����a���S�08��0���('�C�9@���<��֗>��,R����w�+�;����eW3`V�����Kd%k���Pk.����\��#��LԵb�z�Tn�d�X)1��,�L�Sʴ���`4t�A�x�̨��LO���W��T���/$� KT����P�3�o�rᢄ�������ucƚ���o_Pԏөl���A��:�ǣ�.�7��'ްY}��4���U����^٭�?�/�\NQ�,W���~7^0�UQ��s�2^q��I�U$�l"h���/e���H\̻�/�� �
�ǂH��ѐě{���DB�?j.�=��x4�}�����Q/��T�����\E�H'��%�Q��=����\N&��m2��jnAy��}�d@��$"|�v��Wk��i���QO,轋�MoE�rI��3nIV�_�f�J�v 'Д�]�mt���h��z�B&d_	�ߕo0���d���]�IϢ�&$��GH��Vx��0����'G�p���cn�](M�ɩN6oQ�ډ"͖m����ZHT�r%����!��,�!F���M��.��X�h�1|ݠ��8�SSP�7*SPǸ�̲q��~����pmt���/�.��$ 5#��:W��6�֔L.���.V����Гs/�e:a��en}�qԨ��PL�YNW:UC�^Y���S� IR�Ck�o�k�xoE��JcәE�1�ԫ""��i���CR��1�p:��{�;�K��Xp%�<Phy�M��B)�#oYu�H��p눈��m��Xy�;Z��끈�vLq����"��4�KZ"iSF�;�.�r�^��3�b7�d?�mq׀�p��cYF1�g�8�6d_��;ǌP �h@qH�I`�es�&V�i��{��E��olVn����v�����~ �ֲ�	i�!���ֿ����Q�q�Q�N!]RCֵX�%�#��>���,Bof��N��xI��k�͗�6��i�fo�xPo�R��,=c����"��S�t�|����>{�U�$н��~4�;S���D�5JD����G�!<�����y's0վ�z���D:��I07��[��|��{f�v�G:"h�&�0��װo�E��.�W���Ly�S\8
��Pru|�BϜa������S������j���<���ʇ��'���!k0�=�r�e�,f|��-�e�/���F�����ǖ(w'��.W"-�,i;��U���SW�{��ǜ�z�/s�(��x$�a������-n��Z�f�x9�����*xB���D�JW.�5��P�j=1d�𼤄���~]m���b�67�`�rh���� ڄ�=fL%2��eȫ*���1�}Y$
�
v�J&��u�~u�_(���,A�x7���e���-dtO��7�����??r�2�ܧA�*c7 =�HtR�aU���\F(�B�d�ӯ��f�ok�lY�Y�z#!�UN[hr��l ��
��Y �R����ߺ|ą���vuMY��Hꉻ"��\���� 3��>�� $�Ac�&�������pd�U�����ސ�Ry�*��w���u�b.��oS����]F,����T�6�{{J?+�0�t��a��<�j)�M�dЊ!C��)G��R��H�^�x���z�\���s�#�*Z�W�ݾ:P��[{��d�$G��P�ү�\��|D�A#�Ǝ�z4���As���y��ki�noM_������������ ~F5&�<��ףa? �3krZ�,�w�����ϥV�M/P}���`c��d���:� ���s���<D�kK�����<{sR�ͯ��-��{���d2�bn�IE����n#�C��܅mw"��ک��۔�7�T+Տ�`����2LXb�x�����0õ�^aSr0� ���aM��Waq�3j/t͍>C^>���c��B�g(�K���,jZS�±*��ʪ������z��迷���e_�Q(�4���v�ֆ�}��r���xCd��H�%䱂��X8�:!#�
)�1}����g�������ΞZ6�*D���ϸ�3K�B�>4]J�3+��W!k�*{ʮ`ی;��t�k"�����o3���ք�a|�E~�a��s/�L�4�Gy��V��� ��Ae4�eF�4�N�R�[���l�J=P]�ݑi���g���i�=B޸�6%��{a_�!�Rl����� �=FK�a�Qs�����o��7�I �'�>�_��>�]W�F�a�MMa��cM�6C���*�k�/3��tx�(�Q����2�o��D`�(��&����?ݽ� ��bo�Ƃ7��)І-^dMuA:@� T�<q��T^�MAC���Oz�������@�
��:�����W� ۉ"χR_+e��~3Ԫ�rI�����qc�[�����߫��e��@�W����m��t����z�.s�5�;f8�/@D^�C�����m�x�հ�ϴ×
�l%π_�rl?�����a�LK�SFFo�W�D���|��V��D6�q�i��6�)3o�r�z |aT�T���r��c���J� :I��. �i<'a�@��&|���G4�!�j�B}4#ت���YZ�cAp�����Zq���`g�El2�o�?�$V���C,�Oj�Ȅ�
�(l���M�-H�t�ŝ"b�K�|Q�7�co%}_/��y�2��:�^⹡�VR7�N^,UDM�5���Q
o���JXy�,�1t���i |*⾔[��p����A�����K1v���1����&x=����l����ga�pǪ���=�FP.)������%ry:�F��$���E��vz�|��mxTV!���@�ܷ�Fn�
?2��̧�������Uޟt9��-�ALt���Wi0���R��b�I&�X��ځ��>���ӵ�p �iPm�K����|�����)���?�_��u���=X�d�^�Ld�AQ&-���}�q!ʠJ�iR���c�H����� 7��[H�5�04��乞�����j�7��𗢘J9mM�)>Ӌ)y*�[pYb�s	�����pTX��N��pXM�6���CA�n��1:%�m^�;~�@z2m����a_*5�����ƣ�s|��}p�ر��8�� <��x��}!_Jd�`o��,<Qi�7+��Q(��1����K��+��d;��������;C�^0���
��,�����yb���g��<��>�̞� �n�#��]$�4����)��t��f�K�Ye�$㹷�^nߤ�Q��izkP4FzR�1�@�^'/Sχr����X����n�gS]�S�:��q:{ۘc��f�O�LlJƠ5�]���w��,9��v\�g�A�m���y��s^�v���ҍ�N��L����r/�l$��R�6�r �d�`�95����KŜ��a�EnW �*�'��?�Eu܎�l|�6@��%uυC��5C��[�zeM� �#�!���2A�:5<�B���/�\9D�u��2��~��˴0��� 0��xֿ����Ax()n*�$�h0�iK��3�/���e�QɇR|gs	g㪭E���k7V }���N�ć��)�49K�TOJoi��ǹ���S8a��0̘�"�J���}XY�fuJ�e>���iݐ"[;��Z��o՟������n#֮76��VC#�h�@d�X�;Ư���O-�C��s�>k����?-�d��g�y%W�g�}5"�Ɯ�q��g���g毃�|���C����^���\��7���͌ƙL��g��|�ϸ�K��*.��DM"����ɯE����^p�j�è��*U����r�&\
�	�h�ï�U���{E�+IDT�!���CWş�
张�IN}(�����u6W��+J�='�W*�>�	��,;�+Za|pUY�?��;�a�a�4,��H�z�ր�EUҫD���.E�雑ۆ3�ҙfs}���6s�1J��/
-��0V��P�*!W�>>��~����E�2#|����@	�~P]��w�������.���S���B<7�19�P���.��:F}Q1�����ӫ�,�wB�>����'��3A��^�QV�V�
z�|��8�;⽬�A ��^�������8g�q��A<�0�)�t8�����N��^��La�e��j��d�G9b����$��ga�����WL�+��V&����ilgh�e �Ӫ���5�;�����$³F�I�p繁CÂ�&�y`�<W�	�wƶ�9n�f�{��6��{S�����x�
q�Ь	�
/�L�'����8z�:����sQ�Tx�(㔐P����d��Y�q�,j�E�з	�s��^�S��8.��]j���U�Q��8�<�������`����T����;�`�&l�����O�4�8�cU2�F/ez*�� �u�R�.�C�[�w4[��:׻�-��j-�O�6Go.�*�)��o��94�X�%����u�6b�Z��A)K"^XEB\#k ���\�^���N��%t˪^���x%	2����=����c\-���}O������$V�^���wQ��klH=c����p���g�B���+>���b�x��b�S����{t��3���
z��$�B�5� �mc��ݩ�Ed�w$5W�֪C���6g����s$�`�%���SǢ�i��s��9�G�kP�� ���S�1h�i;3������I�����${	d��p.�o���{2}��'Nd�Z�!Y�\�Q/'ׇ��ˮ���}�Ga�550"�x�4������I�-N$rL2}a�U����ܦ�TQn}�LP䳽�XYE�[g�r����~��柍G�����^�G���K+��8S�� �oP����k^β�q��Ɣ���p# YǥQ�����o4)�����^��Ռ�R5�,RO��iK+��+�7�G��UvQ;#�@���ݛ�XB�(��Vv7$8�sn�X㖣��� 2� �]*�~,`9��*����]E�����`2���o��-��cZ���&.��y�k������5�Hf�1cE�p�o��P�$�f��}���Ŏ��E9��>��ed��x�Q�nk���7y�:�_
xFt�.o�C�Bgc<¹������	x��4Q�
d��c�F�1��"%��9ia�h��(
�NhC�&N$�ਖ�|E��h��G~��W�8&H��nI-ɏ��R�O��~n��X�S�rҩ��fs�s��ji�1i�e�h�&6/C�v��K�U}���x��!�u��	���~�������/�tn�1� �&�x���������slX��?��_ ,��=�.��� ������$60��L�
��EV��"�{M��*��.ᗪI����o72`�o�G0b[APC��S~
��6�*�综]�'��>�v9}�~y�8�zOE���.*A��H�J�Լ�1dK��4�^ �)Qˈ��Y��쒳�Щ���O��q�� ��u�^S/&!ۮvPQ6�bK����<��M���(�Wg�P��5���{}��fp�SP����O���ί5�<$5x��ӡ�b��)Ad�����B��i�W���	��x�c��n>L��P��P��Ƈ�Úg'�3�Yq�p�u���1ɧb��y�@������xRn+���ߌT0���k�c/:�8��]��iL��L��G�bN �J-(Hx͔W����$���<Np6+gck�Nف�9�(�7��O�B��
�f�Jq$��e�/C�������U�g^��)�c��-=%�ݖ�>=���OBz;��hT7�����b���g  �?����e7O,xΡU���r�x�]j��Z�J#�	s�ET�nF��@��ߢy�}Ci���zf���q4��67����z(���n�I�Ok��ZVz6i�P}���x�jL�wS��Bn���A���Ը B������G�ԃ��j
:���4�+�$�s�� �O�m�G}�P���ԡm��'�1�h��F8��DS���h��y�IW՜)zȇ�B�"X����;9�g�Q���!��(�rG�6���# ��Wz`�K��^r��F�[��Ě��̇Me�[(�x2��g���Me�%eD��0q��/�^(C��w�f��L,�тE��o�ץ7�� ���ԍa͂5 �,�z�9,�H�HB�2.1��M%�I�U�ѸRӃ�oIj����M,z��C���@Dչ�ܗB�}��;�œ>���NX�6�',w�}[�*o�<r��C;��S/��?��Zm��7�gs-'�C\9�@���
i0�%��?��@�Ԏ2|�&��;e���� �Q�p��Dg 9L�ˆB�����}A�+���Q�:g������C1j�i�"J.�Qs)��[��𕈜>�z_ҟX�����R��Ф�B������%����R��l?saś����q7��#%�I��x�s.�E��ϥ�+Pt�p��UD'pމ8���A.W�b���_�>�]�|C,�&5�����\�X��OS�36 ���KO,��8PjַێW[�ăs(���x����I=�nZv:{�ye����U���CZۡV���&�Ԕ�7Bm����q���߆��B�-Q�5��X��O4jy�r�Y���}��2�ט��*m^�S�f�K��B{��6�[���{�d��z��p���Q�<E�}=m�!�K�G�������7�u���H~�f�`-2�3�����|�z7)ϕ�ȍS��]�m��f���N��<RUNr�y�E-1������N�a/���OXqX��\��/_�j�]�2��s�udCK#6��9M�w�OQ.����'�˦%♆{k�ar-�d�XP�_�W��G�r��d71��J��x�W���puˇ�>R�;M�_��*��AJ�з�	F�\>~ա�4Ȥݜ���-΁��jr� �'G�>��T��^�\b����ر�����O6CF�����%*L���f>��7��g~�����Yvq�j�t�����OZ��05*Vz��ܭ���}�s^�L`�Q�P��Hᴑza��Xc�j�=/�6�.�,��bc#BV����s+�"B�o4��wcJ�	5�F@����靖ꬹ�U%O�B'��bܵ���-Qt�����I}zJ�/U��b��ߘKP�����s��f�tw��au)�&���p�ϕ�Ie��/t�LM����:���+q��&���0�..p�����;a��n5^��	�������9�B�oLBВvM�L�	3���;�uZo)���5$��O;�/w�.){kY�4���7�,S�@�lkX��E�<!��ދ�����¸��]H�e�v�+��Vt21άgk���'�Z��6�sP9C������Z_j`K������� �Y����hF���9���p��}��L������x�_B,�A:ڸaq���)���4]G��o�x����&幚�~?���}@�}� �<�^�#�)�ү4/�N)�����Gl,mLe�Y�@0CuQ&��@�&y�exU������]��ǀ�K�S��o;e-���?N���jyL�~��s�q��Ó�G����Ï�a���j%��H(���y��{��d���^��;����{�dlf��C-P����3z�9ۢ���8w�m��g#��U�R�l
�QE��GM>G1ȅ���!.���6=�;pI�����B�T	Ĭ %�=�j#��7�T0~,j�����z�Q6�g��ֲx_�AP������y�j�h��-�a��#��Ry��
�4kD��s�$����T�����KE��F�f:}2y�K�:�_(WE�����M���{����D��$�������bQ�HvSpHd��8��l�O��� ��4i˭rbf]lbG`��3��K�@Sʀ<�O�³�9=��J-p�A[���;���>��4FO��O�k�s�fu��,j(�{�<$>ؿ�
��������$�������#Z ��6�	:��`��~��5ҋ�R�`�Ç
S����sx8�S ����l�v���OŶo�}Pe��4o�=Z�˿�(D9�[Vs/uev8�J���>�d�w�n}��K\�奞<��:��d��4)W�zЅ��<��\-W.��ҟ`%9d��XB��8����wt<?2͓j�%�ԈP�1Wa��~��8+��:�T��@�ZlNy�B&���g�{ ���O���[�۾��Q��q���(�Hy���3+i���i`W��H�ǵ'T��5N��;�,L�0�C�� ��@X�����<Afy��H�ԯG�F�vH}�j�U����Ǎ�`���c�a'�G�����2<4��t�뺎�������w$9ӥ���!��Xd4h�3��i�u�b�kaˈ�d�?�<�m�d��7!»-�W���5YoٝtI\|�۪�������V��8�K9�3
�:��o��i�Z*��ވrV}W�=lF��`fJ�K-�}G&�]�ؑ��C�T.�(g|��!��%ܮ�՛
�nZ0�ˑ��w��c]E�;�jw�aQ�ʞ�.���ws�M�L���p���ѥQe���'��p��2SD��9��f���0�t�X��l��a�޲��ƒ[��-߂"2[W������6��rUB��f.�C�����E|pU3μ�)�b"�_�TH��h�߃?\��t��y���Ezp�"�K94:�ԭWS�D#jt3C�ǰTI��4 �6��TV{��G���J�ct�D���V�PeH�rK����rw���p��sY�� �3�Et�`�-�R��9vBR��g�]����C�Fg�db�0g0v�ݤ����\8&j�2��{��<)�X�=�����Kx0�����u��??u�����*���%hI�A׶�Q�o�n�u���)C'/R�S�H����)�yk�x�SF&c"�> !�- N�~_ +Aտ��N�*��k���Ր.�a��?ev��c�1Ϯm)fe�dM�)��d�թЩ���{0�VO�O��[�s�
N�=Yq�ۢ�z�,>��Qi��4{!Dy�A7؇��,JۀQ�C�5�F�Y�q~�����5�
q;Uy"&O�f��\^�&]�O�*=���[dIeHZ�m������T{���|Q��0���.S,���貮�GO.H�Z?N�ٓ�>�O
��'�}���9ʱ��m��p(�_ਧK���<nǸ[�p�ݎ�H���䊒8�P�Kk��Aj�����3�9�S�^}�k[��v����<��;�����S�c"Æ&Z�e�T���V#'f�6&0�[j*��1^ W`��o��N^�1��^��
����گ>ᘠܳU�~0��D8�aYԀ)������׾����)+,zW�<Qk���BM*H��gm(��D�W�{���ı����b.+(gZ���~�\q���ް$���-�*��p�yR�1� ��T��á����n��F�:��I�w��Q�,R� ���i��HB��-�v�v�G�������V�r����=!��I�a����Α�_&B��!%��Wy�Ӭ��O�'%��X6�@�ο�>��8�� �A��Λu�g�L9LsBQS��Q�b�9C]]��m��P��7��."��)�~'�
������7M�Z��-��8a��;߻o�!�L-P\�)��I����Qw���w5�����6M���A�Ծ��/�d�9�
:o�'����?X�Mv�HوP��vU� `a�=�q�n�Z䅶;�t��V�V8�q�Xcu�_hv�S�¦;����=���*T=hq�x{�9j@���h�����P&֎쯍 �i΋3�3���[ud�5�h�QI��F���\l�1�X�\�CLL�^ {�C�z�,4��9��e =1ڕX�)��b���DJY,���r�f�n	$��/A!e��
p9zK|<�%���+���2���5yHj[�\�a���u�)��f�l��VBj�=@���5��}��u��� [�h�bt�ʆ�����7�$�x23������i>4���g�[�&֏�0�*�I�����ʗ�_���cܢ���f3�Z�J�,ho�,ܛ#@¥!�8��2V��P���j)���;%`I���9�� )2;yhg/8~6c������`��]7�%�| �[K��Qe:>F�ɐ�����Td.������j>U=#�D��K�&��*n�I�j�_��[y��j��w�y���3�}/ho��ure�̆{V���?d�N��nq����ɹ�%)��g>�?����~��fp
�n*#���s�K�	����s�}��	V߀ �;� ��D$��D�G�@\�Dq"�n;��~�d7a�J�Sm~�xस����׷���T�=�����
*����PQC��_�h��9�rT_&�D�\�7'^���#���Dib-�s)z:C�W��������-���}c^o"�?�z���"szuO0�����­R�P�
ih�Uĉ��x�sfQ|�5Z�p)���nw"����t��������{@�~S5��X_W��x�T�<Y���Y1���C���������2����-B����:��W&6P�3�$�7�T���p�8�/�ň��&H(�\���i�@?���)��Y��D�H��b��t&����2qJӕ�x1�� �#����qg���[���!�3ֈc���Q.��_9L!|uᮓ�~;e�N�TR',�1{���h$��-RI��� ����Fz�Y<�v{��͗f �B,�Uݢm�t��Ȩ�DAHP��V�Vvf����D)5�XÈ��1%�WJ�S��L	f#h���&O�T��ö�5��o}��a\m�Fh8T�X�T��$@�yL?�$!K/��^��5���;�FV��J����8aL�+?�I��gͦ�
Z3��!� *QEHg���$n���ݖa?P�X�4�fd��1�$�_��F_fw�dy�����jWkM�x�5"��A��c�WF\+���
Zc�'g^c~^���ϓ��9	���p�ԩ/�nu$J7W<)����h+KP���S�S�"&h�p�yk~��z�u{yw�X�aY�bLu$ �g`��O�#��2촗��@ �pIvb����h�y��T�A�\��%H��lf��rY��N�9, b\�߬DB�@�ϹI'בt��7�u�Ё3L��V�NC�#�ݪU�m��5�o�ېi\��h�I} $�c�NSĤ6G��V��#�=�['ȣ'�&=@*�˞����(�I�� ;�QҗC�͂C+�q��^�	#e"�:W*������{AJN����M>ό���^攲�~�-KHh7��T�O��`ӕs{!��Cеn1��#�U�@������}�V�l,���~�o����:�PrC��b�#���3 7����S�43��@���Tc|"]+� E�HwY#��W0*��^�]hz����'�&QS���&u��wQ�,����F�qW���� ���{�b9BԊ�ۑw�;����y���>-�<�gP5�a�qצ��V�{����o��iLu�D!��b�$�k�ׁJ�\oL���5q�e��L�s�FJ�U_���X�}��ΫR�Hd��mǍ}�́d�uC��n����M�����Y��k-1�`<\]��\aƢ��̩r�L}��3r[�>�I&��1��#H�xeY�������bϭWs�u?PV��z�بB���x�0��&m�̕����៊�����k]A����t���'e�r-�xD�x�s���V���O��g����(�
R�c_
�W��+�ȀO��x�����E���U(x������&܈��D�]��pQ��h�{p��j@���:��2�$��\'e���F^RA+t�eo��U�{Zʢ��7hY���X؝��.鄉s��9�n�� ���z]|sǶ��X����V�o���R���0$Ý����?f�!�6��=���7����,"!/��� ��>��7� /`�Oo�N���h�m����t�<
�T�w�8�Z!(��g�Fzޗӿ��vX�q�4~��vgy�`q'� �#l,5K6�t��|��Jl�	��bf\l94�Ҭ>��&�>Caq���:Ջ�\�h� �m�>TZ�k��-���M-��ȷ_�Uh�8��>`ߚ\���y�^t��-{��Ir���|;af�0��U5�1����/DR�y𷓷���}{H����j�����j��Q5�����T@���T�:8i��r"�Х?嬴B��s�	�π���A@f(�2���_��)�ݻt��o���fy�_����y�����s�*�4���P�%ì�!uw�F֫#��Gܙ��l�1D+��e�*���Sk��p��ɾ麙*	�����lвPO�M���{1�؟�چۭ�8��WH��Z��~2RZp�P/�K�� �{+�nH9y�A�����h�$.\�u�?Sxyi`,��Sf}���؇G{'����\��j_�)Sk>y@���$W`ү|Y��5��d^���q��7��A�_�d��P��(��H�G=�mbz|�P����ϹOƭr�n���6����i��d>����us�d0�tm1���~{~� c��h��&�8{ �;g��;�L��_8�t�9�c��n�k=-�ܜG�ع� 4?��ì��,3��o�ډ�V�1�ԉN�%��\�\�1m�iٓ�T\o�J�3�Ptn⢀��h��	�x��g^�q�����\N%x�[	�g�mx�  g�����frh��	�qW��i�����O��M�oa��)��2���2e���j�E��{V��NP�k��B�WK7Lo_W\�.^a�R�$]�J����ؽ����"	��i	t���sS,�9aW{3�t6��0̎���K�1��Rԁ+.�"Ū
H�@dRJR
 ��'	5���gh�Ldg���͸��� �����i������+�ʓƷZ�s�9��pc��9�P�f"���b]��S!�p˟�ۀ��H.f�7Ӗ�78nY�RoQy�(D��U�S����"����-�V1�F���xD&��J4)�	����v�ׇݝ B��Ef�}�~�)�ꝡ��P�(({��hא�ܨ��Ɲ=6���HT���f�e�������m�I;>%�$_�g��
Q�Q�E2�^�o~Q4z�-rt��\Ƴ�4ڕԝ�T�$���3qL4I�~�3$��G��2 ��QZ�-`���P[�:Ϋ�R(6���H�+/�$9�OV�s�f��w��#������ѝ�HE�e��b�Y��QH�Iw�9�1#��)>�*nq|��,�%���%�9:�B)�VX������rl�q�GZ*Et����n�g䜵����H�9���{�<�}�^n ����;�����h3�`S�:�S���=��$@/R:6#w~l_���B�ie�5�?��U�c�7�FaXՙ���E}���^kD�����R��G�nNB]�S�,�+��ielz`��&,i__V����{�����(n
I_oc���mE��@�7�!�m$ᮌ��D��&)6�V�8R&�*s}27�T!+��� �8}