��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0���C	�i��E��$��Ȯ��[c��z�%�Nil�P���b�5���E�`bx�Ȣ�<B���i�f�n���s�b�z�����	���Zq5��AR�P)h58@	���NWm�ՙܿ4+������%pQ&j4C��:O6X�?O�cx9u]�l��
��'�@"$p�:���H�%E���(�a����5�ϭ�Ѷ�4u_���j7t�T}� �I6?@��f��`\�rk_O��]�,��<��5h�W�}��eU�>MDDs4�Y_w��I���G�5K����l���<��U�_�..P��S��ܹ���D|~hp����OI�Y7q\C�!�B;��'Do�%� ����n����`Z�p
���A����n �AFP&	�P��G�\y$�pn��/:�K���ƶb^!6�t��:|�_�m8��W�,R���`�8�N��pɦ��U7��:y����1X��u�A�0[Aq�|v-���i$�ҩE��]���NH�>�?���W� �樱�J��~úZ;ͫ����ڏ��cL��]��Z�������5����W���@�
�_��v,��:�'���-����"��Q*��K�汄�z��LT�S�4�T�ץNt,{�@P���jQ��z|��kZᑐ�����_,g&�J"y��׸XU��G6F�.�5i���,�)V��v���>�xy�|�]��@��'(��L�8��)l^'?r�c�B�K9���v}�#F���&�M�b�9�Y�����1����[3%.￵h0�8�GݫN#��"�����4�`������қ�ȫ�a������}�����;�_a��295�#Kx�Ԋ���)�D'���O���~D1a�j��v;����6��҃�U�)�����4H���#ݔ�Dv��R!�=��^�kV�����u��}�IW0��o�XĻR��%#�;�&��d�,�L��ek�vA�:�3Q�r3-�[��Q���ζJe�(!~H?�	H��eݟR�JG�8��C ^&��YS�t���E��Z�������N~��RY��	�9���^���n���b���4��,H_I�������������\/-���)mM8�(�Ģf�]
_ϣ�n�-�y��i:���*����}���m���*Eۡ��D�k�Qa�,�kGU�}�,���dp�odcÿ#2v�쀶���%��/�8��o��^�F5��{�h���� 	�.DP<�{ٚ��Jf�e��CŵR�̎���k�k��AQ�.�euLn�i��6�gc^뷕u~�`�8E^f�2� jyi��Q�I�L̴l��[�\��g�ݾV�����Do�U��W��$2��3��y^a��"�q�# ��.W(k�V�0���\���/5�֧E}I�5��w^��lK��*�[,aN>�k�d�X���}�c��\���_�����0pf�$_��3�F�����|��&6�q�gv7��4�����E��օ�M8t�d�	K�hJ�x��Q��0~��_=t��$Υ�e�i��hDȿKbܕၖG/�q�l��W�`Kb��ִx��mi\�q��@?3�X��V�ӈ:a�y�`͸��&�U����>�o�ڈ�ZO��q��z��`�*g��6�Eo����-�QQ�5���mg�rq��p.6	)aF�C�q��bSs����Ki�b�m�j{�\
�HVK0s��.��R�E�_+��177_�,� ��Z��P�Q����^����d�m!f�G�[�;�!��V8��m�-S�O�$���J��1�eۻ!����~ȅx��iBj��!�<��W%�ե$Z���A.N���N���A,��D�=�-0��%cl��U�j����[�j���[�a�P�j���橱�t1���4=�yW�&.Nf���b�=�A
v��$��d%Uoq
ս�����I6��J�_'��2�<��B�}�V2s�]��f.�nS��r��Y���H�Y �'73�_���SSA̋� ���喦�1�k�pл"\l���g�x������;~^�P&J����x� �}��.��g�y��Yuָ��h�D[ ��b���N"�?{ �$���j�(>�/ׄ�<�
����񳳖NQt1>vh�`���u6�w��O�L��-�ys5�SR�x7Ǧg�j��;��~�}v��&z��H��a�/��MA�2Ȟں}¼d :ƉQJ��P��<@l��B�J���sCƄ� OV�7}m �&���z�P�^,Y��؂/�/k�����N�ܛ�nE?��NJq�ˁ�.kir���� �9�+��VE���)�N�h����|a{��s��71���-9�X�;�f�ө��1�7剚�F�m��:�UlH�����lh�]dg�
�> ��)�����:r�S��}��kI�H[��6�E��g�eu��L��2%$�߶
�l�{���r�A��J�ͭ��R7�͏3��a=�j�U�6�m�����k�r�N�!�� �M�`b��o��B���5��]v�U��4wJ���_�r)��}���m�6R�4�?Ӟ�D�������B˿�]��%�m8H4���D��a�(w�z]l�pUO��������GD��KAn̬AFkZ}ݛ%8�[���/֘_*�[�S�<B}xA�% �j�Lw���{\-&	�Ͻ)�r{"7���uPZ�ZC�H��`,�����������;�<-���h ��h���V!�!�Jn(���l��k���'��RKBJ�Ld�is���G'���p�el+RG��T}u�h�[[�(y3%L:bvX���N
�t��wY,�FG��@�P�{��ІJ�P���VaW���{,��`�~[�U��{yTew-O��G��j?�b�>E������L���?�d�>��S�{��b4���y|���z?���S�1��.��~^���d^�!i����ۏ=�|խ��iЩJ�hc=QOB.X�� tt͵B+v�j�:��-�14����%�X��Kآ�b?�h3}ܽiN�הW�O"ν�{L #�w�m���'٦��:�@����5$���?<�uA�$Hh	�A�H�T�"�Z��eQ�kQ����r��z��J���j��>R�W��Pf 0�%_*�����.����o_i�X�k���L�k����JR;{���N0����2��J�3����D���ˮ�7?����l/�B����*@�MV�3;;?!¶�H/J��w!\Ty#���9`3�3�G_x�!��� B����������a`R��6U?��D!�V�2��v���F����^�b`!�UnJyjq!�Ѥ���}���O��J����^�����B�N.SΫ�]�D�f.&j�g�F}1<Z]CX]nٌ�[�&"�x�@�,����\h?D�r"uV�=�x�7|�-��k��
�W��'ja���ݛ������O�����jT)r��F�������̱���m�h\w�/㎓�匣2��&�����mSk=����B���6����]U�v���v�k:lAv���8�2̓�����h[���@��v��fRXB�O�%�oE�p�,���z����DMۣy�1�3SbcUp>�;�H�\�*OdݛQ!�(t��Ov�����X�Y��'��]���֕���md-�����#�~�J�A�������z�.N^��������p7<X�V'&��l��\�QY�?�%p�4 I� ڮ*b1ۗ
P)�mFڹ%���Nk���G��|FC)�IH��>� �\����H���hJ�_�a����^oa��j )��s�����G|ش�L�(Mh�y�H ��X]���V+y[��#��)����|BX��W)U��j�4|t0��EgpJg熱�`ˠ-Qo�Ǎ�"�^�}�~�L����;0}f�s�8F�	5]�d�Ѣ�h!���l[|� ��}7�J�X�֎'����/�1� 4���k�\�Θ�whm��5��=��/@�ۄ�aOf�.,��+d/�J��X��o�m�BWrw���6:��0�G_NS��/��_9�J����(�.�ocn�K�
cZ���3�B������4�����$�HL�l�贶
8�k����{��#>ϔ���vq��Nk������*��ZQ����],�d>�GiT,�O#�|ρ���4�����ZD0��l
�FF0��jZe�8�<����)�d�{bo��!d��y�!��Ȫ�n���ϓ`�wc�����=�N���͗�xd%�y�T٢���� �o﷛P~�b)�r���c�!��R��p{��q�s�	s�݊^��@������8-���&5l5h�0w�:���v�Pq�b�W;=�mB���5в��o+��0�j5���*�(3�y�f*�2pt�ӛ���2� Ɯ#���6�6�q�:C�,��Su51���D>�306��=���u�����\�h���؄U�-���R���K�Dѥbw7����aL��R,�B�6s�"W�Us��m-��=���xBt���ە^� ���@-fd�x���(X��F�w��r.#D�֠Nx}8W`�!�n�Ɔ x�Nu����C�8���AVWK4S����l�J���d�~�Mh��J��t�ȷ*���v£��u����+mX=�߻�L>�ƴ���d�I19�Ȉ-��\r>m!]�M :o������R�P�
J��̓P�:"t��D��*j�D+�9>��>^3�ws8��|Z^��c@jC�5�P�ܞ�V������P�����Hs���n���a�����۱��h�S�k1Ob��W�0�V�����3;l���"4��J�{Y�j���o�&,�)3R��<Y;�C0	ou�����C-5'3��@- Έ[t����z�F-v+�a"�R�'���B����R�\�M'�j7�ꗮv���	�t���{�D(�t�
��nX��jU�f8���!Me8}p,do�P���ާ�L���9��lb��� �F�>)�?թ�ާ�\�}�*��֟J:x���$_+��'�g��4�cK��=i^�IG'���Y?�	�Kɰ]�D�t�G��s�g+�;D��gg���"ZJ.�'��`�O�ii�X�w*C$'�ԭò��jK�?��h!�cx`��p���e�Lv�	&��y��tn��-�_�U�h��h��%���)���eT������`�r�C�0ڼcV�=F���E����R��_{ٖ�տ�%����ީ(X��-���`ovt�JTB]��ɗ��dPf�^����a����J��(7�G��5F���ZM���i�oʻ�<�"����9$�� ,�8x[,��=P&"AH���§�4+K6���}2B�K����]���*����q��G���0e��С��=vf����[����4�kQ���u����h�۲-j��c;�i�Kǟ�B�Q5��M�!IW�%����b�CJئ�=>�4��"�I��u��$��b�x
[�'=����9O�}��A�8F~-d�0��M.��2( ����d�pͥs=��]{�g_��{��?�0*�m ���a�Z���(���Q�K�h�K���t�\����!QMIa,)���oq���@W{:2�+u��n$������u��+L7z��*.M���f��ĸ"ƆQ#N��E�9��N���%0S��f#	z/C����Iw��dS�,I��E9�j/π2�~��)��?y�H�} ח'�~���ŬX��������+X�4�}:g��D��,�PO�ɞP��!-�s$���H���[���u.�eʗ �+��U+��bX��H�R�, �v�zX��y�м~;3�n���Km�:��@40��ٴC���5?��Y�D�e&	�|./�Q��_F6����h驛���~ڨd���v�����tYAx���ؓ��0*ܼ:�QmL����f�l��(C�$0Y9ꨴ����r~�����:�Y��ya,��M���s�#lH�O��o��B��+#��:����n#���nZ�>����9DtѲs�T�-�$��\h��n5~_FDٹpe���"�EKW�k-�"�'��3�#֜ ����o�"?�)`�Ր�v:�m�^S�3�;�rv$�eMyen����ʪ��$vo�XU��{J�W�Q.�*�0�#y���AQ����	<�y��$B_�:b�|�༼�����1�����!�Ćr1�����1ƌ���4\�6%c�җ�U�j�V���R��%��0P�`i���E�e߯ﭞֵ�yycHO�a�!R>a�>i�.k��-!F)C�QJ*$�hMjŀy���9'���ZU���#B[!�m�n4����fY��F��4^}k1��:8��;�qB��K�ɭ_Ց�U��j�ox@'�x��f,�V���7��n���{_
SR�J��?������rn��ܮ��4#H�コ�����Z3)83���5��g��2IS�4}	�9-����x��4����q*��3�5���L�!�<�k�⩋���zp:F㝱�پ�7#����9(�v�߱�QrxmP��J�lgg���?�����.����`�k0�Z�3������l�3�n3 ��ଊ1{�暫�����C^���|B�1�� 3��=`�Je�D\bȶ/�._p�oF�����#JGU���$��#r2�xt:"}��4�h*�g���g���G�����L&��~f�Q�@������i�z��JJG���!���t ��i](f9�pP�̔Wd-Ny�̟�J�*݄]1W>�+��4��ݏ��N7҆�4��ծ�ra�x�=>��Ц�C�rκϗ����0@0m�i�9q/�s�h��Yu&/gDgޑv��a��4����Xf��5�i�J}��-���e`��t�_(귥���6S�0O��d���G]77��Z�*��V�K�un�GtN\���R����\�%����7�7;I�O�n�Ɛ0m5�:x���o�R���'�/���O��P��k9�.O6�W�x�ihp$��	��U=�>�gaV�u��
�u�uN�P�L<H[��2R�bd��4�d������nH\���Ȥ�z���`;��ŭ_�=�Ј�����+s$�3˵�n�t��%�R��eи��Q=��bX��^����tP�f��6�M�O�zP|�-q���aN%BR�s�Mщ�Y!X[a���_���&�; Q�.X���)��3gϼ\'f��	�y�q���kP��_�XwZ��:�|������Ҽd�:��2	v���M��L�hղ�&�����_�l ����,Z���%�EM���v���:��UDn������k ��O�>;�x����8��U��]��q��7}�g���MM`��R��^$\#w�t�����<Zz3B�̙��p�_D\(���x���8
Q)d���O�{ؠ~��⯔�i��*n,<�_ыW�nE����<�㍴��D�G�k��sRԣ��\nG�N��,ѷX��s�ՠ7�2͐X��R���x���~����\�s���ɺ-x���t>3_��W���)� ݰAφ��F��@w<B�:G������~b1&�#�ԏ{�y��=C" O���Ti�nL��5�_!��� j��?��d����>~U�M�vQ���{��X�w{���ي��˺���z��Υpr C|����}��n9&:���1��L��f���[�7.�U#c��|e�@�?�+}���6w8�I#��Y��ɭ{���P@�"��}>00V�)[k���Ya�-����ȸ\2A9��}\��R�<���iً����U�x���L�jx�"�b�ӆD���X�߹�mn���δƟ� ����	rK�+������#t�5x�zs�ek[U/6&�TY�4|�6���q�����3��L�?�ր?
�fh�s]�.V#΋�[�I�'��ڢ�7�S�����B��	��̓�m8�?���	�����Ș��A�'g�ӷ~��ʿ�-+�D5��wemD�s�����NdcwآD�Pj�s/�3�l��W�����%�:���4�,@�a�.��nO���oBwu�w<<�]`ʸ��!?��O/K��K��!:��H@�{{Υ��Q�#���B�		&���D�1o��<�*�����f���o�W�~ H�+!Kc�Ib�l%�T`�7�5^�~a��,�w�D��"����V��dI��A�/�L�j�߫ oe�n�����>�c�i��Qʨ�O^�1]�揺;�8��hp�:�c�?㉟�C��/#��r�׶gi�	���M�>槹31?�ű
0�:N������˲���Ղ�s@ڕ�4���Dfj[vq9�8�!~L�=ޠ#�-.�����Ժ^�.�"V���k��a���M)Z����Қ �~r�]P��k��gg>�Y1��A֨��=�F �ʇS_��Ŷa�i��E�s�p?g6�r	=�[IDȽ4��!�05������E�h��hGQ��3_����,y3p?%'���'� �w���3d���K@�@���)�9�=嘔z��]�M�p�>�������q��3/ ��xH�t�t��V����*�U[�qH_Q��e���b�I��-�qæ"�J�	@�׮��?߇o?7���2=)�E��縥�Rc�ts5��G�`���N
��!�9��pE�}(gv9���!�L����t��$�z��JB e�4x�V?��<(�������N��Ɖ��t�;����K�Ӯz�,���G
��ѯ���l�m�B���{a�P�S�e81���/�Ɂ�I�u{�_C��YI��R��%Fh5���r>��H0ͮiϡb��&������#&��wGl2ɝ��M��JAR��z�2�����́e��ڋ9	K�Ұ@pF�q�LX�6�,�0l䘝ߏ؋��&M�һ�^I]A-~<�N5�
��M�A�L���������l�����.ޏs�ɣ����`��/�gd��㹐���c'�Nx�b�)S��z��ԫ�77>��޸2������~�������j �ޢ�s_^�k�}��ÿ'%i�j�d{�z8����
����b4�a�~#b�?�{��,g�����_� \g豽�l���8�X���ܓ��'��^��HX��������-<�ss)�����&� �H��$T���c��Xxvn�����~��<�Ll�6F`8��_�դ��=e˄L̆�Gj�_:��=�*�:vn<�� !��B���)G#';��̘���EQk��A�K�l��y��BLӂ�<O��h˛��2 zG��s.S|��f�18�^��흜$䮁iJ�����j�p�̨`�ϙ[Ƨ�揄?����s�\G�nz����a�&[�;�Ϫ�9]�;��y��!/ZםTw�^�PȁZ��q	r>a]�#1�� ����u6�>�S��0�$$��y�v�^y��ޖ���#\�ʏI���wިxIB���L��N�[M��%;=�k3Ct�}���W��T"8�9�r6v�ӥT6��PU��?�]ˬ�����du�{�XԶƥi%T�b'���V�`�*��3����4�V�S�(��q�-��::q�%�t(7��L�#>����޳���hm8I��|�;t"��>�'L��$Ƿ����������'S�\���ٹ٬�P)��v�$H��`��6�eI�]�q�.h,)�[���f�Պ.�-��̨�2���U]m��x��/��Z`��
t�ޏ�0A�~͕&�7@��ݞaI���� �σ-^�����W�0�5�l�"�^�Oxnl�?�>�����@"d1g�=�+��d �$��d3¢����)��)�"ɏ�5�tJ�{�a��	��9�\���l�Y��
�b��R˶�!ڥ�����X,��lr~6��1���Վ?�Z�������w%S!xD!��M��e'��@,���1-����G��qlW�_�������.xw���L���PQ�ra�C@�;����[��T-��GP�j�[����\�R  I�BK�7��*~Qm#e��Ӝ�> �_~/RK��3�a��S��G�ºTa�p��OՂ�S7'SE	�O�s ��>[B�/����k�Jaq2 �S�q�'}o|�o�pJ�eJ��l��r�O2�p5on*�(g�"��|�(��rG�'o.�B������0��җ�+v���}M��|�!+e 	r\����d�_nE���t�+~�H�L�S�M2
���@��d�zMm�9�S"87y5^Q�4N�~D�.D�uss�s��o�m�M�y���Շ$��h%tG܅`�^h=�`$�g}'�2��d�sY����"��
*���I��3g�ͦ-�V�z��kML!p�f�l�
g�T��5�[�2����?��,�}�	$q\�_��m"ڶ�hQ
U�� \t*:S�1')a�K�F��_��.����vܚL�?� ܥ���� 4<\55a��AY�=�*�ۛu&�XBE��@b������,��u,�&Fʸz�B`�\����������������VJ�!.8ȯm#��%�.{����"�Is�	�aBG(K��Ϩ�p�_��So��7�gd�
b�<C�r��l#��\2����fw��b���s�U]��Y�]�ƹ�2)�[D���.j:�O�[8�u��1
�(�Ks�ok@��1t�Q�P�b0�5��)\9��pD������B���Ѭ�Y]�[��v�d|W0�V/�/��h��<
�Z�Κ�K����\ģSD�k��ʒ@V#>N��N,�Z^���[�pU�����	���(�u�z>$���w�oE}�j�64KR�%ey��J~;�!E�E��'mx�@��x�Tv"g�u*��}�����&�=�lE-�q=%������oS������P; ���veͰ��(�rp��,Oн�=�x�d��,�@�|���|��ë$�q+*���B=�K����&�u��k�$bzћ�  7�������x*��K�"����%�	OŔŀ�r�S�l���*I���v�I�s�>mS-���ڦp��A����Qa�2��B����ܸy��8��@n�dL����Sm˾/S['~kч�14�ͼs�1���樗�+�s���������V�Q���Iv���A�����y�E����O�Z�@�O\�������� ���>����u��LO���ϒ�� �X�&�xR+!�	��{r�bq�8��	]E�5�����n6�Z'#�l-l�$�M+W��pF<$�[�����z���'����~z8-R����=�I�����pŏ�d���vq��=�0�����K]�º������u�yR��/+Y{~{d��q���%{����1p�G����(; sЅ�6&��78��+S `����7w!�\��j�o�CW���nV��|OW��U���O�z�Ϧ��t���l.V[׼e<\��Z��)}v�tP5=M��C���ۻr@�����W�9DI%,ӆ�@�������a�\�OJ�n/�z��֊U`}\S��(O�1h� |�r���T�g��_pOy��79O� .��|A08�u��Máz����a��.�䐀A4�Pm+y�(rL�[)4'�˞�fE5�p�� H�%[��w⻩���q�O����X��Vv����-'�d
{�@�dL���W�4^�)�	P��uq�KEIu)�O��]_m�� '���CicR�պS?�i��ao�%G��F�q������z &,\�~�/_�/���Տ����U�p,ƺ�@�����#/:���B[9CL���)]&�Źy�郴Emh�\M� =���T��F�:�����h.��t�M�ʖ�Q,]����W�)�L��\�Hs��7-�v #��'�N��eJ��	�>(:��&�H'��
�&ҏ�T42W�c�O�)�%����Ϙ��o�`ZȮ�|�K�=و4C�i�T���0"�5[l%v�aز��{7���\J�Yz0����� �d�Dz���/�
���`�r�]YZPm�#��P�ކ|�`�y���&���(�	��h��,z�`�"M:e\��Ѿm���w����CBchִFƺ�l��$�]�;���*�������voT�'B��Mb
@�U�b��]τ�Q	�1��z��A�!�5D�3O1�!�
ݘ�����|{5��_`�D�V�ۇt�S`��Va1̘�F���l�����w��X�A�N��l�	���k%wu�_䈕�r��+÷+���ߕ���K("0k����?�
1�;ܿܤ.�= 9��Q$����~����p}<N�=������R��pE��7 ���K��#Y��>�P��&�@�����ǵI�����o�%nX��uǓ��T���$�<x2�s-���[QD�q�f2=\��������!#;8JP��nU���e�r/ά`�9�9&{��q��F��b �����~t�kR(�%ȫ��],����$�$����/�p�wV�t'H+[a����#�r�6=�\r��<� �Ѧjt���-+�G�I�[hs����M*�~�yWJhS�E~�>.R� ;dm�~�a�5�Z��,��5W㽺 �8bUZ�-g��	��6�ʋ6�T�+OU����*	�撊��2�|�QyN%����&��r�͖��0�cw&k*"�LO"���Ͽ�J��S��3�	@5�I>����0��)(����z�^Pqiq`$}�g�'�h�o��ۨ��c�Q	�\��A�_*�7����!��v܌p%�C�=����'�S�x��� /��r�T�q����mY�fmSazD���n�����$�Y�����:�D�*��p�fK��X�gb|@mҠs�͚��Z㝰]}�����F��Qm��֟]V\|vm5m���Cm�о��JrGC7O�W�|��/9���t��%ߺMӠ��\�gB��&�l��xz��mL4[�@<�,Z	U��ߒ��H�Y��Ņ�eJ��(yvѥ÷G/L��VE��H�'��r���)�L�eؿ����P����6Q��s�`YGa���J�c�~)n�e���F��ٌYx�������� �a�i�Q�����g'znv.��T�5�:��N�~�L�k;㧴��վ�Ť��h*a�}0ͥ迸r�gW�J�!����X
����<����ξ� �:g�e�;��A�;�mkP��H�F�-9D��Js/�v1�h�5���m��]�C����
JK����� ��f:��<Us�2�xl^���`����kѯM��yo�G����6l�yy���=�k�Y�X���V�@|7��l�V�us+�w�D�5�!ź��g͝B^zzAz�h��E�?���7a����uw�fjX�y�o#�G�����ӣI�M76�g���utk#sz|��j�WY(��S
CSϮ��#9�x���x�4�@鼝mlEyj��j���=�jZ܅�5+Q�0��z���l�����x��E[YH�K�)ʗ���#ٞ�� z��.-ߺ[p0PT�_<e��D��l�PYv��O���&�L����Q*!�5D��@2�QU/��*�k<Fj!���J�t�<�b����nۦ����r�2U&k�b�2q��vT��7M0�;A(�{������$tݬxI�1ղ?��M�E�����������x¤���	��x��l0����6��,��?��������'������C�%0�����	2}��n칉zXa���ץ�jr^��Mbq��_qD��@#q��֩'��H�P��,Y"��z�s���m�!赂��-T�a�D��f�ߎ�y���>i�]�=$���`��w��⚷�KwI6z��лo�^�z��c�L��eAm��nY�;����!�ة�(	�O�lIU�w ���
3R�|�	�[C��Մp���������@���%.�͒��V���Ẅ́�Q��w#���4�wY�Un�I��g�9��hsl�G�E�F����
��]=�w�-��!�
�@(Vq9�dOvgl˔�8o#|1	�6���}����!��\p����(� ����N�ѳ����]F�˩�v 3����ڬ���ʩE�*%�=���䉊f_YT�&:A;%���0�:��c�Ņ����h�rǫ\/�Q�S֦�8���%�C�C��6�GG��BX.������JdE�1岡r�^x�s,,<���o���5ЭVZ�у����Ak�_��Q��*FXw͏�f�Ws$a,�Qhۆ�H�c�������\йQF����,w���ŏ2�_k�F���*�X=�D8lF����tw�C|���
f�n�wc�Z�̲�Q":֍�J�r��)�>�W�Hr�[�M�G�#'�$�LʡS2��y��?��x����|q�U����"��lu���3[���K�K@��$]���7|:1�����hP:~��z��/�9��EjJk�%L�IMX����,O�{�2t���s��S�:�=Ԋ6��\�R�ۜ�p��A��9D���Jm36�q������j�sa���p�R0 5�W��U��$���ޓ�x,<�h�Q46���r��p���yB+�߀��f�J����&�B��"Ő��`6B�����Ŧ�%�׾�!\�����_�,��pu�+އ�����!ae>
�����߆z3oz;7�v�����a U���n���S���[s�p�A`vEF[,~Y��),m�sˍ�NA]���}G� �ҳ��ut����Cٱ��gh
-Ԓ�|=2/�j0՞��
0�}oU6j�+`��׎�wK`�n�G
��g�lIOA���?cG5<ݽ�)kxԯN�R__�� �,)!�eu.��hC���Z1�u�	<cڿ�B�޳T��Bh�	��&��'Ap[�����6pF��""}�������y�����M�%<��n�7��1���<<Ѱx4s_�K�_��<r�O[�n��d���3b�𚗋W1�!���Uu{��,�'O&���a:�r�}�*�)�g�̌�=	�\����ƦV��78�{��_���i~�Y�0�9��V&i�ڸ)'�N]>,k� FPci���$�^y�}���':��it��u�։�� �=|I��$O�<�����?���%������=ک>�t�y�P��w�eȢk{��b�Y.�%.M�T�5���J �Bs&�|6��\��a����ElIH�3+�`���V၂�<���C� ���ҍ��ږ�8������� ��.b��N�.�0mF�j蘒jG�fƋ��E�_�6��A;9+�l1C��.Gۀ����*�x!s�>zS� ��@�vΙ���"H�=��"�Y��9y�J!p�d��� Ib<㛕�����+��lA������/��M��z�7�TJ���3o�z!�kb� mC*x�[�7�)��v�c���ڍ�չ�������
���<{��ƐكǍ��v��s�p/�S�>T��m`h��QFHb�IQ��EA	l¬��@$��`��6X+r僮��A��J6�sE:沘}s�S&��kYo^k�L�3
�s�e���1��h��Dn�U�MC��P�]� ��}�O큰�L%d�K,t���╣0GL:��[�=���q����<]����j�/�����Es��jƦ�Y��T�����X��rh�+c�������$5C���]>������D[1�M���Z�����-�c�pO$��ޯ�^��IK��٣R�^�V��<(�ĥ#Riu�bGxm9_?���X0�Z��)Z�Ϳ���&b�,V�Ϟ��9�9���S�0�i>BuZjcuVw��i��̕�b�E�
~��ϛ�a���#�,�5���sk�4l�@�|�Y�R�y�Bj�+�~��Є�Ui���>�b�Ĭ��[��Z���k���G�5����K�{�ȝ���W��3��w�|u6�vJ�����@�|�]�o:fǊQ�M#Y�It_�z]+�O�ܧ�6��4����#��I�
5%)ف���zM��!���`��� r�WdFr<<�1P�0�Ӧ��a��J�Ǖ^��M�!������d�9J���ĽH��?��M�J�5�쯰y������u����5��_�E蝾�@��x鄊j�䷑�1�U	���I�h���<3D���.���.~�sm���-� H��� ֳ�ZΈ�����9�oY_:�B����	���X�˗�I@��m�U}uG��d9-:8�G�����{	P��ൡ����L)v+�s���	��HlM�bG�`��:�RH�(#�hP�b�*��?t���@W@~�s0��Y+ʥ � �l|�ֳٜ���?���y�$g��^�4_����O�[P<J�U��4��Zٴ�NCW5��o�:&K3��}te�y�Q�:�F6խ�'�u��x{ X��^hj%Z���q�҄w�K�q>w�5r[XW!�eh��g�3��^]s;��]&������gW��^�����ަJ�8�#�����AJ䖖O2h_��% ���)h����l����W
$6�2ww~���P�Gm��N�.�E�r��57�ﳘ�YM�*U�&g$I?+��9�9�S�JR�E%�x����q�4�X��� i�a�����RW�
���J�8�;�*9v�KpA+��0��%U4v�9B����iO|��/G�{���,:��2�ʸf�h��)o���/��>_��:�i>��a<%����������)oM����7�<����5��ԉ���̭��w�X��?���X��(��a*m��>�v>�=d~C ������zD��X��o�����;���~���~	�j�ط�,י%9H�'|�;'��ҿM��LφG9�JiN�M{�WZ�ٜ�gyw\%+`�˳��,��+��.���xXS�l���"�&6ğ�θפl�dt-�7�Q�4��e���5�4��z��_�R�c�?_ci�@��F<�:68��xS1�1;hT�r�J�LŪ2��6,�Ī����z���� �̛;ȩ�]��(�&�����>��	b7!�(2t�-Te��R�5����(��8G��ŻV�Pn[W��� �����2�I7 ?è�k�C�&6� ��YN9���6"�����z�f������0d�a���Ԗ�YE����
�sf\_8eص��uސU��� ��0!�_�2Q��K�`���i2����~��K�6�D�\*��T8�soU���A�1v~�-��/��\g�qUCT�6���\sN-��G0�ڞB4��2�s��(4��|��Q�ہo���&n2B&��<"Lsaٯ�����#ta�"���!ֶ�Q�e]\�Xl���
�>��_�3�j�K#�&In�Jz!l03�+�<B��y���)=XdJj5��b�z�Ab�øy
��[9��^�k䵏Y6ڄ�Y�C����"�ifIq�@6ҩ̩����	��Ї�@����?������]������n�s��T��XY����`H��0�/�pZX��I;��w>U���y��6�u���l��Y�� ��E�rtt���QT�gQ�&	q�5L�y�]����@���,l��@��t#��ѾfY�y8%��*1�X���b�C;�@!���!����ݥ�_�NL�v���Zŧ~�%]�@�_ڧ�)ĕ3��ĕVMx��P�W��-���%���/�ZK|l�9����]l�� �7��L �������0&��e���Wz�}ɲye*��m��M��U4{�A+�ug����B�E���ܦ��L>"��42�64�a+�cl���,�ljf�mB\+�����wI�(6���3
���R�%�cŤ�=�K��aCb���l�z�Dv����h
�̆�W�K�~Hh��e2� ����� 3|R�s�f����Q4��g?�g[�ˆ��;�s��g*�S6}���WW�?|��+y�JH��Տ���J�dT<�-УZӚ�ѐp��?&YH���At���+(iD�%���8v���4"u4�V<*�j�ݥ��g�-�B,��M�n6�{���� �0���8㑁����if/N����^��A��(��V�8R[G��<����J��g�&']A�.���K@����
�۵X�o��#�%q���܉dM���]O�R�����4/�Ң8��X߻�-ڠ+?4����#�1ᱶ�M��:NC�U2�룹M���͜��p@��
��{e~����oF������cR��d��Ч~#Qlv^�!��1���JZݾZ�ꎮ�䅎B���o�[hl@�hZ
��+F��1�+X��[;���M�����kz�}�n5�VrH�ǀ܄!]��� ���v�f�dƅ(/���Ú�ܤ%���N�V[��=����\��ҳ��ZI�A�5H4����w���H�@L-�:���{f�~jN8�)^�WK����B�v�Z�M �scĎ��c�eI�N|jtA��S��k��!~��yyn�Jl�ɣy\c���zd��k5����?��!������k۬|���}.���;�)8`���!���WN���7t�ďO��a���F�^z����h;G��ÀS1_1-7��G��z��o����� ��l�x'����;���45�: ��u�
 F�	��s��}j��.�w:ʢv�O�j���n��%����ӿ i0�O����}�5J��sa�1�Ry��1D���������O	����q�t�����'�� 7V/�����B�.<�V6�r��ln�������]����E��@fa�"7�;� {��2(Lg���"��e��oz.J�0��Y��4������r1�4m2�E-� �K�q<jg�I������A@��*�+1gi��A�yP�L�����_���m��X[_
�������=�4�h#�uǦ�B��,��ػV�rr,z%�di����nN���
�L���Г^C�n3ʿ���w�,�b�RKW���*:Äw&�	�x�H,��-w��#��4ÆEyZ �.s��6�� �P�[�>hۥf�'W� ��ɫ�]M�
��x;P��a�f1����Cŋ���AzJ8u/�!'}Pl�=��&��}UDJ�!_*�j}a���PtM�z�]\�T�]S����{����`2�g�RO��(?&�`��ek�gْWJ�M��cE?���.�����$H�K�ȸ��C��j�/�������#������������ݒ)�;[ct�}�v�O5B�}A��������o�ؙ>���{��P�d�Ģ�ѿnE|���� �7�D2��h���-*�1%- }��`>�-o	�5aw�q#�s���@O��3���b��"�x��O���}ln�~y��Su&��2�XD��N�ڭ�ć_sr��"�8T�A���:�oăQ�k�JR����[�N	5�p,ULH8F#O��Y�j<
������~Z�z��]�F��GHW��W�{o(�u5XU"����>g��K�� ��.)
5�q)��������D�l��Y3��e(BWO#�'��(�V��B�F�����	}�,]����j�q��oe���|;�����8L�i7�+���S��;��t��0���3b�cX'ד��b����]��6���U���G�t\�0��A���<
�G2����!EJ���I��<'�� :���8�eư�r���pU�5�!�PV_e����λ����{%��+?�r88��Wq�^�GD�xz~��xCu���-.xx�.�Y\�묉�"�@�q��A5L����j��$�
���S�>`�ъ����j+-���32����Bڼ0DF��� j����d�7R"n$
7�=��[���q��i�]��5r���1#-t���=��0:Rv�ט�jT���vRE�{�K=6
&��*�`�l����aZ0�����z����Y=�@ť*����4� �F[h����1�� x���s:2�Ȱ{��E(ڧ�~/�W�<|T~�����!��/��Զ\g���9���ܢ�¥�:����t�L|�L���:e�l�+�`{L4��V,A�.z�� �#s��%�F*�J��U]\�����`T[�3����qv�ɨ���D遍���xB����q�^j����Ϲ
�5	����|]��u���'�z�8�N�~����C���\��#?�[t�r �q�`b!R�h��Z�%�����8�3ٻ���c$]�I��x,yc���;��ޞ����8���7���j�1N:��7�=�uU�lqarC�`�+�{�m�nC��ӥ�eMW�������G/��ũ�}M��:Ax��=�mt�:�=�C��gq�-���j>��+ߓ�Rsh����i��H���L�7�_q�hXSj�l�Ԧ	#��O��(o����t�5�7b���y]�eF�D�8�I<�q�y3������%r�n�K�n�^��
��&�B��2�d̞y���w�V���X���Q����<7O&t��F�BqqU�'ǵ��=<����	��$���f0���	e2p�X��ҡr�����☶V�w�R�>���|�������0�1*��+�k���]�	kymZ1M$ߛ^#c�������w%Gї���t���(���!K����y�$��
I~�G0�{�q�b�vz�v�ф�xTJ��PGf�� ��	;{�q7������#�O�~q��L�<Q{�d�'��̥g{Z�-��s��wN7�H�P����_Ax��������Y�@)�:N Bt�L�[i�є��WnT��(N<�<�$OX�B0-/��0,�'�����᪫�@��F�J|Wp�p�?�h���n�L�>^ni�V��Ϯq���ac�H�5���(��,�0�
y����qWmy]Au� HOz	[k�yQr͙&�Ñ�r8��Wʚ gd�p0D�WV��.�e@QL�ڍ3]/��|��Ԃl{��g(� �����~����ꩍ�B�ju���u�&�I��ȩ��w�̓�Bw�n���Q1�����<��K�i�:�M�Ģ���#jgX��H�g{a��K,���/�Ho�W�g����ﺵr0�e䫵h�����M�����GT0N��X�߾�h�wTzHgC2��M�iup��p�p�v+;�Ԝ��(M0�YTGi�;����f�a�f;Z\C�����83c=��N�n`9{�LT��m�� "�ȸ��V2���s�gꇙ�n�\�7��=aQ�U�x�+}���Őņ�Tə�X�@�k�3R�e�Ǯ�,:���wg>���,��� t�5�r������=.��7X�-�x�!���E��(i#�7�v#���Ę �/h���X�oZ?�)/��nT�����Pp�&&����J0ݰ4#V��u������P�T"W�Q0'my-�qG�����ǵe�[�s��,��d�2�$��YO�yy���-���}��H�8&�`��V�*����RTs-���qi>���w�$��3e~�{����1�$Z�n���_Ɗ�G	�!Y?38��;�6�:�1��~'Q�]G���v�t�:hG|y�
��~��F�]���&��8	��#�x�M���+丞�"��b"��J�|������?jnNT�,�>;qUDKZ:1�C*�J�1��g���N�R�_��K���,���&5�o5JB����W�Ws��1��`ĩX��R�x����[pD&)��ZM�2�ra��Z�w0Pw�Az{B������º��ۈ7��є�%\@@�BU�_pn�|M
�٧���I7�eݹi4�#}��kyF�\	��	�Z�]կe;�jvg_��Y
��J�0��Ec���:v}.�)'�:�g�g�W L5�k����L����Z��٤�?��Lr���nGO*B�==�tn�y�b�$���j7�ɪ���'EVy�FDRW�I����2���d�,�<9�ԑ6�'a̷���.�7f]>�:�)}�XS<x}k	;������%cA��z���!�s_��-�Z^!t%:Ӽ�H*O��0JM"��?��|�d]ʁ{��:��Ug�h�6a �,�/�%)y�x���o�Z&�h�4��_}�B�!X��鮪"%��od��iy]ڊ&L*�K��sԑ,ʡrPG�z���� �d����vC����6L�0.{U��)y�_1�ڈ��C�-kٍ��N�{�Z��	�AX�֤k�xG��`�X$%ީ��P����9r��|e��疾�\ͣ���O��c��� �1�;N~	��G��F�j��L���g
;˙�}�6s<�~�6 �uP�)�a_�̊�)���'o�|V=_o��#�]M�;q������]�X�L��L9����
�H���	��F�L��Tg���������1�V*S�n��^�.ʥ��z�q�����&��K$y�5��b�^����"������i�b�ŝ�Ǯ;ۧW�]H�nF&:	�9�����[?ܖ��Fq
���NY3X��N�BQ��;��j�*5?�F�`��=t�{X�=�i����.�q����+g��g^�
�^��o_�
Agۏ���CIhk�ϵcL%�4����	��l��#�s`�zK��S�W��ۛDU�(��>kh���Vř�$��H�?�R�7]h�v� �Hqu�A~���TJG� ����J��S0-���{�u<�ض�g����D�CA��s3
/�(c;��c� [��T�"J@]'��Cʜ��Aǰ�>�Y��bo���gs���xA���Z�P��n=�����y�{��Nĵf�*�j|����e8[�iN�=��z��O&���xʽ��n��(�rpD�����QE2�p�O��'��Z&�Re49�,$#ܻ����F��`0 8qf=\��\YL��1�}C�������_+:u(����n��R�Cä�����7Գ`���W=�k}�Y�S��P)v:�(���n2�ҜϘ���'r_��N��ò�>��/@XB���ҽ���P�8
q��P]�I��C03'��ȕf��bo��CL2����Q$�j����8��8�H�Y�,��|�c�y���k;;�%�\ڳ��(�Y�士݃�'Ar��HD�|�i?��V���{�f?V*}tA�6T�������v.����1Pަ���`�l<ȳ|���di�^X-��[N�$ ��?�*�'�"��Lء{��;��9�qJ �͵�?G5&��Z�Z}RZ���0h�$��b�a�P��D��&��όܜH�Cj��N8΁-�������t�����#�B��k��n�� �j��b�Y$2���s��2�O�҅�۹ɣ�)y4�