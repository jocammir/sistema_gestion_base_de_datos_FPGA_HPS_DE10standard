��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��ܼ��e߈SU���AR�>+�y$kgG����)!"���S-�e�%]�gf5Դ���s<G&�,H��gX�
܎­SH��76���kEb���Z,��O�\��X��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�s^W���0A}�����L e����EF^��ຬ�bՃ�-�O�,Ю��s���[ţu�;����!6��ROk:���P�y�?�6���Oj,:O��q;3�bkHR�C@�H}A�:��Ւ	�����ux���y��Au��%�X�c�N��0~�'.d�H���V��TM1����܁�f�=�1�����B��*�Am�ȁ<��N��^�Lh%G��26�k�$��*K*e��|��z���L�O� �9�/�,�7�|z�>L��W�v9�HX�k�t�Hmg�bH��K���i]��A�*�&V��+����?j�ӲN�Lo�P��P�&��>����bo+���7��s�%����bz*QV͜�����Y�9� ��Z�(�&YHJF��`uo�`�ڴ��<��Ot�� y.잏R�<lZ�	�LH�GP%P"#�}�$�@h��y�^B��.i%3�a�%>��΍�I���f.���X�OR1 B���T�H7��2�Y�mf�?���lHŜ�a�cŦ�����tB�Pb	�25@LL�ݞ}&:;a�z.N9�~<�c4�>�hC�y?>��`Ȕ��e�R8�-�z<	�
P��:�,P)�]�7�N��(}u�aLs�|�e>�����˼F�G2��pf6e���^@�̱��{��̄���ɲ� Τ�Kc�ܡ�)��O�P�2��19�.�d�ƕi�TEl~Mhwi�yâ���� ��d��XP�z���uь�W8:�9c����������H�q�_�������D�_���Ǔ�E�H���e�$U���tUIUgB�u�&���߅�Zk��� c*���k�B��将���j"�(}�9��5�p<��D��?��4ȅ=f��r���f¼'���yI��Y"fB���O+"f2�S+V���MēX���<C�i����j��f��L~�)�/�Y�8�����������0�eC�D�G>��>����L	3�@�uA�2!�˦�^���q��O��XŻ���;��t���<t��#U�r�Fj
�?�A��W�@�t����q�t�^[�qcl�Z�;R�b�^b��#�_���{0Er�}At�-Ƹ���n��e:�������\N$Fq�E���G-pl)Q���v�܎�B��ڻ"@'�N♂�R�}[�� B�V;B����Y���"�;���#c�}qZ���1U�̴�1�T�����ҲH���WQ�p��2~VS|�"���'��p�/#������9���t,a{++P���M\�҄F&U.a�1&Ip���d�_Ņ�"�DwL}�hU�YQ�-�A�h��R���e�_�N���,��B�����L	W LȢ���7��(�.��� .D�����rn�v�K���c��x���:Uڢ/��j��{]���9I>�]����N�c�Dm+;`D'#�i�5I��.�B潤��������^Z>�����@�={�ݘ�����I6���N���l�w?H�./a2��D��N��.��m�dnó��C8$oT�8U�[�����x�������2��N��F�x������lri�������� 㯢N��0��ml|�jd55w���1],M
a�,����T��#���x�Ӏ��n�.3XE��a��E���	=��t�a4 4p�|�G� T�z��l7�W��J�����%B;5	�	��� %1����r&kx�#9�@Տ6�!��d�\M\t|&�<3s����Gx ��G<�
T��37�rh,�$t��9_@�>�5'%$$�z�l�e`���Z��o �W`B��u����fN�tA�H���lN<#�T������*
���!%��{�R�Ѕ)<�`V&�ж~��II���t��^�>�	��.�~�ZD���ƕ���E���i��;�i$p��>��d�%	Y����Z��^�:���4������x���W���?}�G����3�gb8T�9���V��0p���V�,���$r��2���8�����m�0�oӤ��t���f�����tz��
�6�[eG�\e^�b#]s���<4o���Vt�U�J��;5�q��p�::.	���Ԅ���P�uŞ�BCeJ7I%[K�Q�I�������3T՝�xH[03��@P�GX�U� �Z�޹B�	�	D	��G����S���Ո�C��ɲ TK���Em��>$zQW��`Ӑ�����8�  ��Z�7`��PTJ��A�t���<��j$B�>M��@TP��-y����(]t��_jkTvK�Icٮ�Np"YvU��*�+��ĖfQ�S������%��V���h���l<:`p�
�)��n��-�8�Ha�����ëb_��`�,��Il!�]�:����pb���VXg�=n��` �V������߭}�l_cSja=��a�h+\���AØ�V��Q<uv螙���*�CL�W�+�Ÿ�0�[�������n�d�p ⯰eզ;b��:>�{�҅��=^ē�`(�Y�{�/�D$�V�G\�^aC��m��ٴ6dxD?ЏK�k��\`�6�I#>R6.�X^ E+l��Gڠ��2���OF�)�:�c�Խ�ؼ]N��� �����,4Zr���6���
 v�o6�1�	FmЇ��^ G���a��|&�%5�g�����y^QX��F�D�
����+ɯm����9:���ꑂ�����ڡ闎>�ĺLǻ�lE�{���D�wζd;^���mbh��^������;�H"CԞ�����#���&,���4��������z��}he����d!�Pk��;.U	�����^6��?��ՍZXbx�~K���� V��9;d����_qx�����g�GF�z�����u�U�;-Q�v�5��h�(�OT������y���J�+�z�m���wO%:\*NCs���V̽�B�5�����I��,�.S��Ә�y������fI�k*�{����xz�]g[�x|�~�y/��T޴_��zy\3�4:tI���JHp��Q�ʝ�y.ᰓ����G��`k��}�d��E7�xN8Zd�R���}��(�'���h��4ahG|�!g�P(�mo
J�gɓhaZ�pK�^V\2�je�}`��<N�{Mb#��%'ic�:��\c�>b�R�$= ��xӥ�P"���׀j��Jе�j���HZ�޵L��"���FՓ��Q��"V�����c�ù}����Q�2H2���q�7�M�^=ލ�V�[����[a��1�o��p7ŉ��ȈYPsv�>��O�Lz�cP�C�@��i��Z&�,r|�`�ܵϤ�CUp1OS�4���kC� t�)�p�5_��)��(ppQ�ӡy�[�M���5�{������K��pO���A�s�Տ�5%��e|������}�4 ?q@���z�3�����۽~B P�uw��H���jZ��ʮl5���m�&{���$�Y�?ij�5̜�e`X�#8K.^�p�_Xd�J�H�5t��hD�&��Ĉ�@g��[����ܮ�7"�Mą�p��ytᮥ��Q�.KR��$��m$L��,�9J|��i2"m;���=�
� @��|A��4�1�]�f' �_L��0�J�}�$m;Iu�-��{q�-&-.Сc��X�g��F��f����3 뽂)J�P���q��&
�����C:ӜDڗ��E7�S7h����U���~]�X�;�{S���#�װ}*�9�	��˒��7Z&,��Q�3�U���l0)��S�l��q]�����1�ۥ62��Tn���%���?��o�g���|���"��3>�;Mߢ�]rm��PsWm`�	�y�F0=V��Wd�	�u��n�<J�bU*Σ���K�����(�6-�L7�$h��Z�����h`�y:����L	�����=9=l
>���W�D��n/��:)���I:/��"��){��7C�#T�;+Z��6�M�oE�QeE��1�E5��?=�?2�dWԘ�y��TB�ԯ��|�l���i2^W��ԩKW��ز�+o7��e��r1�aҖ�/[�����C���z�Z�D��`��X���:&���)1���>�]��j��Ɂ3JJ���#�P���n���,G*�b8N��m���&�V��fh'�x��@mސ��w	���`�5�$�L��.�L��}�����AY��Ѳ����/�F����@,�$�/9��X�h�N�%�7�m�_	O�i�eGށ���x& V���1-�'$������zz����X�kn5���I�)>�ʛ5Y�Ö�>RE�pn��4�[�5@!l��,|�ڏ���Q��8tY���U�_+�CRRz���)���]��pRb�s�m����v�?�,���T��n#��7�g��](��fF���i��`.�� X�](�M�*�a`�.�+k��F�խi��q�
�.f�S��%��X�)�\8��Ɉ���-���d9�C#:G�xo��@�PwS�Ѽ���r�ߤ"�68Q���]=wa���B�$���68짨���Z�a8U���O�t�[���B�P��GJAe�72O9ȟ!twt���?oje'[Vp�t��>մ
���ԳJ{:��j�p����K�����k��'��Bv.P��0Y�W9��L7sQϷ3N��bѠ|��c������&͙�m�%5�U�������|Tf=~��2^�J轁<�9����@�^�9C�N�d�+�g�SZ&�;�}V|b�z����zbF�Fx�UaJ�L�^*���~QT�k�������bh'��c���HʭG��k�Zxr[��T�"	��4����Vs���}y0�N0�٥�1��w~��G6җ�n}}f�e=W{6���U	J'�������?����3g?�Mڎ_`�_8��ʙE�&13c��B��muM��''vG�|��m�KK�;�Z����b��e@�d�p�.�Q��f�.��,+�fbc�F�̻���~e!l\8�4�!�X��C@%f�Dx�EE�$��Kh�/�����M��>A�U����ߊԌT�9@~v+�۝Z�*�P�}���R|dO�}��[�L��\VɁ�X�w?�mUe���d84\�$��E=�<+���Pb��.ы��k�q%%䌂$�b�x������~E�cIw�).�#N����\uؓS���\=�9�5��ކ�*$�@MNb�RT;�2�}���d��M=�o��[ t�C`k�ְŲ����@��v���ࣿZ�%!d����;�(��e��r�Ee%��)�2�����qfi��
4	�c�x�\���T��V�ٱ�>�:��_�������d7l�SB�֪���q����15כL��<������أD�����*�ސ���L��G�z�eN@u
��k߰j���]-���Ӝ����Wje+�;����a��G�q�W�X*�ݦ��B�hT*�W6����[�ְ�(��q��^����lJʿ\�V��ҩ��ߌ���a��C�k�?������F��y��¦��U����\=�Ʃ����fMz g�,/D� 7T�t2�t��ɕ����Ux��0�V����H�ֱs��z��/5����'��$�ߚg�|ڙv��?dcߞ�B���ɲ�\�i��<V�)���?���P�����R�/����N�L`��q�U�	�>zj`�\�&�������Bm��Ş[}�����B
�yȐpО_�>��NH��B2d���z>��ͤy�_�A�E��yX��Z����i�پK,Π�F
�ŭ��@SS��D@A�:V��ކ�c0�#��GmҊ��6��FC� cO��z��p���|HE)�*����KD�tn��x�F����� ܹH���>���ɶ;�"���n�(x~��q��yp�5��1�7���T��-6c�2H��8�#�|�Oʣ���(��*_�fN%�WiF�|�v��]Òf��(N�k`�9�yn:Kk�E��7�{���1t5KW������h��:�ub�+���[A���\�������M��� Z��ki���,�%^"x
s��z�����'�s��#@��"���ix���(��m�!ד��g�dŪ�Wy/NdK�鳺�?�g�*X�,~Gi�^H��y�K��d:<8lQ5yé#��]��S.�Ss�-ݻg�3�kc!�{��o!c�ǀD/�25���3c��0ԣ�q�����*��䋜]~}���1,�'� �4D�!Š�+51b��$�(�L����jzJ�9`�N����VH��+�p���	C�y:]��D���Փ}��Fޠ�y&�M�	Hq(���8��a��ޓ��*�h�)}_�ڮ�Rg����r����~��-��D0�8_�'Xjvd��F���M�l5։�q�o�뫻�����Յ$笉�lB�;�eA4\Pi���'�]�(�����o��>a;�wgD��3y&�LU�DE�e�����<�_�*��5��T��.�7	�t(!U�Ѷ��V'�\���Cb�& ���\�����[B�ࠡ tmR��"h�(��z!o�1y�:qٍ4��D��I�v҂�܁����@FE-�9�(�$tJ���W��������;͐\���v%�_���
�Y���.��`���*X�̤�� ���5^J�S{ks�s[~Z��2cx��jd�x �Ls�B��s�� �̀*)�����p�[�6w���;��9dg��چ�*q��
�Ak�яk������GMg[�CۺD�Wn�P/1Zo�>�%T�Ī����7���8md]��8g})�׎���6z�>`�e#Y���/�0ܗ���t#?k�lϺ�q�����=��f��wk�Y����.�G��s�H�����ު��b��ܮ���yP$���SHZ1ɶ
�xW�3#.D�&O��1,�F�j{�^�a�a�D����é���d��+�~���pkO_�TC���Q��B~+��W�G�����\u0�Z`ooQ+���w���:>;ub��q`cq��L+AZ����g��y��Qu�V�0A�0�Ò�Ҫ֨��0�v�y�/j A�-�<�xP_W���/,�f#�!��~q�D��C���U�&�<^�>�#���
��2��ƽOb��d�qY�'B��gRĻ�����GQӎ�!�?�����`����~�
��	Ω��p��G��A���z}��5HY�������zȖ6�uSk(܏��mxjva�~+$�<W�-�J��PE:^��<]��y2��n��2{z0:���q�t�P�O&�#��٬w��2<\#�F0�>�^p�Ȃ��Op�z�g\RRy�7?S�f='��Y6��V��Z�Ru�ɨF74�;њ[k,��Q������K�A�� �?��sm�`��s�f Y���kn�!n��N�p�	��"�*ˀHP�ݰ�pb8�`$���f]�<���=��<�= �����D#�v*Hj���X��r�y3'��c���A�p���u��-;`�_�<a{DR�L�%Y��:p�������B�F�~�~^����<}�*.���Zcn-h�!���܋Wt� L���R�*��N�]�S=�R-	��|B�oŰ[cW@��j�bt�A�Q��¨�	C}]j�bA�d��)��iZA��$3޴ϵ:����I�oo�ס�}Ja++J�'�i��y�Po�	��Ҥ�,�\�< ��O�:�������J�'��wCG�!~\��ֳ<��Иkw�q/,��{6Źmv0���o�Xۭ;��5��jm�"�Y�%�*���&E�ooAT�./lu��Arc=Q�f��f@a��C*K�SF@�����<�y�����B����Fyk(0��S���lv���n��G-Y�4�3k���뿠��T_��	�����T�Z3�<2�:�mQ�bG��f��3ߔ�f���u�G���lv����'C���6��P|���蠇;�&}�졲�1������G�+�m9�흈?�Gs_���Iܑ���Ɨ����/
�~���LKlG�a�|>������:@8�/N(�e��zi�ΐм7Q_D����[B�ʣ���)d*~�,����
J��Y: !إQ'����ס�n�~���w��otP*��t��2;ؙyE_�t�pGPI�U�k��& 81��?ܼ22�Ki�n'�Zb���/��Q#���`��E���z��g��d�j;
����">N�Q�LDE��S��X��%���<RYڡ���) �X �>}`=��̧*kѺ�d��-jc�GS���<:��J '�@,�nO�gܸ^x�%�=�B��^ؖD�� �Ot�M��U�gA��/';2���|�g��X�R�q�$�pA���8�����Î��d�E�|��O����ښ.��g/\��礋v���xٮ��!D]��KU%Lj�µ���.�@8v�"�����՛�^�����6ni��$��S��$@� �!s_��"�q�e$��ߺ;�>���CˎHV��7�cΘlQ�K�8YV����E�"��9�O�f��6 �\���v���N�T��D�Y�{�Wyx�t ��c� �袄n�����I\6~A4Ӆ��Μ���oH.��9��0��rg�??�$�}RA�E&U<xW3y��<n�ϧs������~6olg�:�����)���Dq�f;y>~s(��c�l���K��A�{���'������� !#7y���V^�������(c$qkײ�Yw��?9C�g���
���Ή찚�s��S��oAg��u�Yv[a �y2���0�S� ���X�� \�*�%dm�P?=������2E�&�=z��7��V�����=jf�CS��kX�C����F�z��x�w�~K0p����d��}1��[���"�[� [�`_I��T�,q�1�qӘ8�-z�3��¤�Y
�K*��9��6�t�,�
���	G>2��G:k����?��~\��v"�yG�Lc[Iq�2�����!��p�*c��DuS�v�y}<�(.��Z~|��>�	0'��!m<'B?@gb��}K�҈�z1b�b��_��y���
D��w��tm+������ ��C%�]zB���Ϥ)N���������,�G��K/o�j�p������a�����	�� O����J�p0�h��4�0/z��U����n�~6bz��=ƽC��=�;�c)B�zG/Z��;\��	N[��������y#��.�R��vo䞝��VYq�>�������sA�u�5�C�d�*e���dUMLY �F���KH���- 1Ff2 ���0XkQg�=��k?I�Uh�CZ`wB����Tm�U�#1���罝��xtC�6l�s�u?W�T�t�,7 ��FSD�t.�J��P�a�i��=;?3���-���
�a��ppF�%� ���@��a���ˢ�p�t��(�G�����Ğ�c�O�����L�>�C{�wӤ�VTY2��?m/
%�.��($�C��tO���C����m�x *��֨�;�H����?��?������FA����eR�D��쫬���
�`l?o��v���ɕ�A��&	��~�yƉ[(� \�-�7�ث�Q��F[�lǪ�e����c˨�.��˽�Ev�d]/g�FU�뻌=`���w��/Xy� n�s��5��g)�V#C�n�j��6T����v�k)�7/��Y*й�8� vt�J�G���֣��'�q�!���a��{V�0���f�%Vu��&߻�hn��n��2�l��$�=J�-�fsΎ��,�lؐ�r�t�MS���͂�)B�u����H�����3L��}�����ȝ�-CO���[�wO�V�Wj�u��l��wi����v�jb�t�([���š8.�\<3��Y���jKaD�oc2IȀ���⼠��SVk_z�����i']���E�N�$t蕍Da��'�ړZ2�{��N��f(��N&��f�G��]�Ws�����^��$�ڊ����&8ٔ��}��ߌ�v��L�T��F
��21���{���}��Ք���/L�&%̥�d��\hI�����}��K�?iF��������DC�u�lV#��!��x�Z�sP5���My�<��v��O[�W�EF}9m�Ȗ�S}?�f ϗ��J�Ԇ���ZvxėZ��6i%���uق�,��5l��%񱊍WT��S��T�g}��on��Ot�ḯ� ̢m�k��.��Z�.�,�k��w��,K��݅(3�#�Dȱ"O辺$�;(y5#B��;^eo�W�+�e�ُ�q�Ԫ�TrC���N
f�ʶ�G�Z#�M�>
��X]T��,��Fw6ѡ�f^�*�/��H�k�C~����� P'&�H�i���Vg�.n }��iUÓ�zuIcmA��88�
.�fX�Qn皞l#߱ju<+��ICP"jI��4�'���Q�����J��g�8Hnhvwlf2p���utAX�@f�0��
��/�푖i�Ѣr�W#Bd�q��\)�����͍J�1͵נrh9�F|�}��~��JsP1Lj#����L���x�$� E;V ,��T��U�������Z�a���\Ɠ⌼^���7�U���p�;�s���W��x�1U���	LNJ��kel�9֪[������2O9[}$�bIi�Di�.�:��l�����d52QW�z4������cry�)�4��k�7C֓�e���c'/]�Z%� �<�v�
��eb�I$��]�Qb-1�F�}��i���F]���26)L�)RO����2�Hha�m��|y�Η��y����%��|޴��;K��Q<����h��!?6n��u���׏��P��H<�-	���2�����؅.����sa94'�!�Hj�@A���6����K,���^�]>̬���*��x5���k]��5��7��"�Х~-��UNz���N�ON��wUY�8�;o��L� ��0��'�j�.B��:t�%;���B��~l�m�UlEL)�I4R �CzV��X'�i��'�D��^�0).L�)������7'^����C�0�#�;gB�:��xzb �Οs�Bt[i�y�T/qzR�� ���U�ͤw��8�a3��rkHb�L�r:��s��;��$�D��Hj����V�;�t�����/#�Cn�Y���J$e��/�%C�c���;�p��j&���+���@�R�5������ I�Jnx� �jvfj��A�No.�x�!5�l��i�&W����[(4NV��0�� Q��A�Z�`��6N�G	����"+�����ݵ�z�R�dC(�龐�u�޲����t�I�lk�[ur��c|��{���던��x�S�7�Z+�Zupl��?=�Y�M;�1N큹�(vb�rNo�_i����6���d�_B�
���e��J���l����+l �*������M��sbR��9�k}�o�ӲCF<_�?��.x[������.��}�["b�;�.���c�EXƜ��
��o�\﹜� �u9˞�Z"�i�Nx[h�3#�����?�+M`�0X���z�c���>���gn*�R�?Y8
�z�!1M�c Ao�*�����ϡ����X]�j�1�-4?�`m~�:C/p7���ծ��nϬ*��Ǥv�{�y8,9�?$-$����aO�O�U$paj}��R�$�c�����Uc��'�Qw�M�JW�V�l Q���7��7Mo읎lY}��
A� tvh�ii��&��D|����r��=ő�֘4�j\�Sy�~��o��D��>���M�Y	�
�.�Z`�\��ro��8h��]ڳ���'L���)��~��N׃�p�����*�6Vkwބ�]E&#0��Gf!|[3��0z�r�B���_J�%�a���v��ۨ$�e/��7oJT� �|�Џ�Orǆ���T.m�}V�x���>S���i��yr�D5m�Q����C�rԼ%[\Q�v����F�K�t�'n<��`�r�mA��!`礭�eY;\.*��p�Wx��v���2o��4vk��<H~��BS#D�l�=���ݵ������p���~�!}�+�Tx7�B�� *]����[��$����*f�"�{�Ǽ;ϵ��i��� #������y�Dx;rru�� ��1�;�z5`���F��α����P$�P��fH.o�Zf���P^�K��Z���YJg삀S�����Y��u����S�(�\59bý�C]5��U�� ����>��8��F�,��.�����׎��/6 i��|-@x���ܡ�� %rL�ז�T�DAU����|��w<���	���(�]�RSk�c�8Ga��Q����o�S+���ĊH�͍�����	G�g~݉*�ؽcb*><H�p�����ʨ��s���V�Kl��b�`�@��DyN�TJ�D555��iIA�:��eYԮ	�� ����CԺ�)I�#��Q��a �����j��)��6Y[�n������dŇ���j��Q�8C�BE�SdB�W����w(s��?�h�m��>b�l�B�Vn�^0�iX��������)MM�lv?�Q�(�bT�v�ԯ)q��]t�3���Zp0O��X"AWXXg�POn�oRx*��=�B/��Rp�����根D��א��mvL��]��fNl;r�c�H:�b�$X�!t�뫃�:��^��F�;b�ZV�EyL^�*P	�[����a�ن���{����ҿ��&�ʩf�%�EɿH�a���Q�r{n&y���eC�j�߾�m�d6� %[=��q�G[h�������ח㖦)�;�_��DρTHǟڪD�j��H�z���t8�,���t(V�t2���җ��J}��q(e p��F�Ø�NA���g���1VISgk���4�z7w��?Lf]IH2����ܳ���"=`�"��s�[�B>;-�w�_H-ڜ���_el�&QOa]�^��A�%P�X��An5��6�b�����䔥pҦ|Ʊ��N;Є�2x_f�YЀ-Rm�p!}���2UK'@�	G8��PXO0/�R`l�ŉ]GZ��[�d]�3A���⥺^4Vy =�|�>�N���p���q��~\C�/�+$�F��a�NG2�?h51d!��.��	�#ً�����`ɜqA�ҽ0+�Qq���$�c�����c� /Z������� �����$y=��o�Z,�Ix��e��������C��(�"���Dt���Rd��r����] A������ �xV�=��!�A��3�'��(1��ɀR?j�����&ё���_��D��&q�~�3T엯����ƀד�[�<v5��,�瞳���{HJ}�SfR��V�����K��2A���EtBu|�\`'"R���|w�*D�*l3��D{8�5:���R�Kmp���6����;�zP%_�EB�3n�	��W4E,������F� �UEع �Lk�J�{Xe�$"��]spkF%����]��=�bO��m4,}j��#�~@H�E�X黎(W��^��2���]�ݢY@�RNW�A�'�ZM�0��>&Gx�K==�28D�J��3�9 =�@zh�9������8�i�`��aܒF�_�C�,.`Ts������m��}�`ݞ��އ�	+��[H�}�	{x�'��0���W4�8<�FYydm�0��GZ�g���!@L��%͸�R�p�BS���qj;!��?{�	(\s��/BDo�h�K�S�ܺヱ��]��.�Hq���[�	��/i�Z�ϰ��-y�����\7�XWE���N7w ���y��t�RL�@��rT*�b`�b8�2��zhA�焿�)�^�nW%cN�I�H��`� ����шtV"$&��c���th���ov|�:�?��޷��\>˺��f�g�(�F�\(�����c7�8^��==�Oؿ��� '��)�\N偸��_o��)7�p���5���_-��kG�^�6_q�K6#��Z+�Q�D!�h&��L!)���c�7Z��O�:��z�$��0�V5~4pD��!�z:m,��W���y�S8L&�d��_���3�Y_��U�o�0�ړS��ܨ0��/`�	���8V�������@A'���/o2�z���Vrn�B���'W�����]������Q��B��&h���� ��$EhZh�Ni,⥟o�N�N��^��OV��d�5�Z�0���T�V��G"������yޏ���cpb�]��	Q��͵&�����%% s�(���E���s"���{������v��� �Q�B����}X���L1@w����	�A$C6�@I��-�>Н5�⫊��H~m�pv��y�rF|���x#�ܒT�l|���Mi�?���j�bp�7�F'C$E��V��e�����/qq\<M�q�K2�\PL�H�n�����:0��	.|����%ܰ&e�-%_����Z0a�c��`��R�
���^Bo~]�>
�;*Ŝ�����zgXM`��G��S{�0F-7{*3�J����[��?ܟ����-Ҏ�d���(�(��>��7��L�z)�.J�/��U!�wU�8rU��T_l(�=4(���TKL�EPhȼ�BW��BoxK�g�(xLͪjo�;�p��˚���j-���kĦIk"z(�8��-c�������=�f��d�� V��$�|Ij�M�	:�5�6r��a��`&���+����oF$]�^��N	>4hw��]V����Al���Ar���lv��AU{�Y&T��`7|���Õr�S�T��ZeЂ���~}�b<��� �x���d4=���YRk�'V)�SuEEM�=���������i�D�8��F%����P��ԡ%vv-��C����Xj����z+v��i��ơ�7w�N^�h_�xܐ.'���2ҭ�t2�sXz�t��U��C	gL�S��=�[ڢ��\��J���k���e��@�Bg_�+(�#��o���4��e���|o��0[�Ȼ+�J�}
����Q��_��D������^X��r��!T�w��.�W�0��QG3��E���k����͠�ZX�3�6�ڴ���R�G�X��Pς��,�ͱ�	�d���V�ˎ�������/7���g�b�b[��J�Y�Y�Y����|s�{0$���>'kL��!���_�$�M�^&�1�FAo~�ڹ@QQ�D�&����?G�B�:�����$��dF�c؂m�!i����ҷrk�h����u����������M��<Ӽ�F(��ATa3���b؊�7�d\͚��g��LwqFG�?�����>��{.�N(�ç
�oЉ/����{{b�s�*fj�rh�GDX���s�\R�3mr� �*\��zqI�n_�����01S�q��u=13&>^� je�T�v8��K��k#����g���G]5���W؀��䂏����[=ZYGթ�K��%�%���͘�_B� �#��M��������C�����	�)f���xb3��[�ѕ�9t׉�Tv��ڊӒCy���p]e���HWh�=�w-���$�-�%�;�vd)�ݖ��T[l�
|!6�BY+�:��r�m3T��o`6�fBa�E�`l�W��]w?S�J��e/�G�x�.u<�IK��������Yo]�������PWF�U� -)m<�K�Ԅ�*^�_���|�OZ�eh{p�8���w�-ٹ�)�Z%�Zd�]�9����'W�.��R��zX+ s_ҝKf^����6a6!爱�돧O�,�������?�@~T?�{�<�\Su�7�ٳeu�ba㼶�4�w炥�G�>U��������`4�������Ę�+n��F1�}g�T��<�YD[�i&��LVa�3�ȅ�I��h�g<R���F�I�m�XL�%:0؊�v��u�(�f^�G�K��|�~��{Cr�7Qt�w4��er�T�l���3b�[H�#��*��!X�����W�ZU�[˒]~O'�f3�Anm���z�#�W7���pD;�Zw߄�vk	���&�$��QY䱺�s}�O� Ԧ��B=�(���~���f��������Η*�k����d��x
�ޠkj�X	���N+�>��t,P/��d�#Z��K���պ���w5R�7s|�����]�H�bAt��.��?��\��/C��DK������F옐���65�oպ�z=i��z�g�5�y��ѽM�?�}a2:���3�U�����>�*�ˁ���ݍaI�î�@�2��������	r�p�C!��e���l�2M�0|aeW#�|Q%�E��)\�}�@K,�$�i�]��ˑP� ]�n%1�": RLT�U�����WO UՁ>њ0κ���M�)i�8�v��M��kK�mG�ċHE����îY� �~g�x�w�}b'���(�x�|W�O7�C����P�*W�|�G�5�M;sik�����BJ2����\��R�"�����j�p��m��F�N!ƛ�'7�J�Ct(�1~g�+W�#L��Nn��A?T��$i	j?p��$	���dvb*M%�|�3R�0�G1��!"�b���(t��������:��j�\����T&9�����4P��A4�yxHne^aV.��B�h*�=�"�2Q�d�Z�X���������JG���k�����T3p���IfJ�8� �2���"-.oC �F.� x�!��< ��XI�l7��9�&�vo���Aw��V���ꦺ��;���C���KH�FFFj��d 0{��<j��y�`��֦x��_�l�w~�R�;(��sQ���f�靂�GYUZ�z��>~o �W�����\�Cd��Q,0v�W_����x1C(}�N'ov�r[���Q7C�ٷ+e��6�P�Z������K���5�i�u��i�7q��m����y
�}gu�j`��H�=��3�{q�%
M�)�Cb��%����k�6	-��P����v�'��|×��c��β�)jI�An���Cˏy��=�+U������u�7@�*�~�,�$����	��#V�n��>Z�K�F'��:ӌT`_I7���B�֗�Y�،����0��ONQjΖ}�0G�rY']��N�=�8�c&�~���;�?��:K�L�����Ph!��g�c�q�s@��y�qi�9��QV��.$wk,�*���d�`
1q�5�B�uK8�B�`�7� 8$Bo��m��͎��
eά���:�|�ЗMo�)n��"�"&]�^� ��z#��3�Q���>ρ���v>W�;�}J��v���TU�����\���_�`>� ��Ujh��/�d##�������Bp��6%�Ծ�����j*N(na��}���������k��"�@88QP�:��VtxD��/�����x�����/a��j�U���	�T��&���+s$]�rhfQE�� ̟�yc��9���s�"&j�ͷ8�hRN0_{���wp����d% ��֪�K*|G>�Q��i��+- �f���u�q��x�KO(EE6��Q��F��RC���s��M�#��j�Ƣ�0]��(C��!VÜ�ecZ�HB�����b"1Q:,O�Wu�w�n�5�1�}��U�p��$��~l�B�/O��^D΋{(�󿯰�S�E:���_�n���n)�|��>h���F��q�O��ă��^�e�GГ6gu��J�?x����^"} �s�NM�Y��Y��;k=肹�5�Z��F��6FV� ղ��V0b��%�������LHF��0�������A����a7,9̵�V����l�T�)V��By꒱R,��.1��45q��&}ϖ`��h�Q�$W.����>DL����r�p�ɚ�J��7<y����}BZ��3��ƽߴ�P����"ת~jk��@��\�������� 02X��}��L�e����I�ɬSذ۵GF{��,�8hܸ��"����l���^5/�4�CmM>�6>��'8������ܜ5h�l�2Ò��U
�F�S=/Η�h��=���oy�7Aq�KJ�z��Ь�ͦ�k���@�
5$�:f�3�&3������Zz��,3F���f��F�ĩ[��d,p`5��Ӌ�˽*������mS��}E���q��X��5i������˿�V$�1�V��eN�����!�	�F�(��	��S���fea�$%��ZȰ�bV�f/jq-�W�G�-�C����P_��y��SK��Jq���<�L�mI�|)��e"��&G����o�vD��Ȍj��jT���z/�:z��]���æj��{���%�=]l��h;�kh=����xq1��)�+놫�bS�~h�FD�����\���-��m5�#�������EV����<Q~��az^ ��M[��=� F����Z�.���@��u{I8�fp%z��ҳ>��p��;�E}�S����J$|'mӶ4�@7��A�.��8W�ƚ��Us�1RJ{����U����O	�G'�2�;��腙��r&N�B*�e�n�P�L�Nh-�D���U%��d��nCxC���].��V�o,-I���y�Ξy2Z��UP�;�G����f)�۪��K`�X��y�zߐv�~J`,x*�_W�N=c��pl� �=1�� F�(0�d�uo���vwV���~m9�b�bGr˷F�5��p�'�u0�m`�<����;�#����@j��u��cR�H���k�@/���U��K&�#8��)�m4�S�tLS�Wt$3����x)Q�'	����z+��C6^|��j����=ƭE	m7���$��	�f�J�e� 
��  �)�~����-��ɐooH����S-m�Y�u!��JzQR��� 0r��������`�Nh�������t ��z^�h������J}�!�M/�sNQ�^bʅ�9T�܌)M�Q�5��>D&7�Zd!�6�rr��5�d��n�%��K{HO�|R�d?Mo����)>��L�M,��Y�Q�)��ג�n�<`�ᵕ�*�
ә�@��H�$�إ}^�H�$������d�� "��ˋ��D/�����[�ρv`�k�	�a^�������a�ķ��vi�6�)�`�oD�O.�~N���'uLGC��=%�Kb�6�B���BfZ]*���º��jɏ�ՠ������ǟ��
�}�a��tɚ�D�.qi3���q��[
�ߺ�h+Ohù]��<(#'y���EC�xa$���甌���c�"���R?�s��kۧ��m dP�ŦYa<T߯}�2=8�GO�SZ��&�.D��͠ZU\v$�5�-�r���gT���c�ɩ�d}� ��R����>���	�g?@ȵ�qG#���N���z�^��K>�y���¾o�8u���^.�[�m>{�5��� ġP�Hp�.��4�rr]�����u/8w�%�^
�^v���~Ru@�5_�Q�o`*�BI���ݤ��L�Ϣ��<���)xVS���M0�	n�[`��
����7�&(h�!��̻�����$Yt`��X2���׋��7�K3��N��@�H�,z�X��TQC�$���wE֣^����-���7���0��{�m����S 2�:�1�����$c;5�� ����lp���A��'|R�e�l��`�o�����pd��}!NjO���ڑ�J�+�^��5��@�=iL�X�B�B�s!��U��P�B��X@pOʿ[���A>�������~!��,�0+��M:;�J�+�����[�q	�9ᮚ�'Q���b�=t�^���v��QZ.�[����}�o~JS)�'�]��K� F�8�c���6y�Q2Ŗ괐J�ss=/�Uyw��
���io�*n4���i<@�K�v_��*��45�s�ㅵo��$�;���ٸ#tΜ���1���fu)6���~�&ɜ�!�qcY�,(���M��\I#�7s�-�զ�����Y=��pA�"���o�:�����چV�Hc�y�?�.���K������djn?�@��w������*,�ފvo~�13͌�S��"ש|�"�X��&�목��P`>���G�Z��޻�� ���dJ�lc�K��D'�l���ۖ�����{D�1)��;0��6�~��|LF����,'���|{�����O��R���ߔ�7�i0oOW.�~�C�',f#�A�����aY7�µP>�sy��ILf�O#{��v�K0�N8X������Y%Qu���C1n]�x�f�iw/jp=�ih�c�,5ۛXYa(��ȷC�9������`�P��Sz��Zk26"H7���`V���͔������
��jfB�ԈV�Dz.J��r&EΤm0༎�I��]��J͢S@߼t�Z⾏kBvb.��0s��i�V��N_� %����^*;nE�|x���	a���Zp$$�B�[O=jECʛ�߹�ߤB�@�6a(�n�xh����N�+���"�~�M���m��w¯���A j�r�,�NL�Wh��^��	>uo��֐n���Ձ��[��5;_+�n��Kn��$�~����n���U!������r.��Ő����Lj��{���4^��Ec���}�ܖ�g��=��gz ���K�-�#p\��J{.�@�L�B�1R�,=O�5gi$&�iRΚ�]%�$�[���#�՚���nO��_�B��ț=+D�A�n潼�#��!"$PJ�9���g��Ia
X���P�T�<
R\7f�����_�d'ۛ!N�5$p� ��9��A#�E���6��er��ӻ���[kd `4�����E����hH�\6�~��h��=��c�7�n؎]>�qu�ӻL�Nt|b_ޅ�VSw����c�V$&o`4g�?I2�QO }��ݬ���:���FX����*������,�]�÷+f_o+ �x3v
�������E��N}�p���hC+=DD�1|'�ÄΧ{���ˡ%[�ٝ:νV(��f�&t(d#%��jm}V
����/F:�5�0v�c�T��e#��`��8�T���d��f�#ƞD� 8&�^0�6d��w��L�͎t.G\���*�J���kbf?�=+�Kԏ���Tǩ�(��r$� c��C��4�%����7��w�]�љ�1�(&0!�6C�'<q~ e����8��O>~/~���t��u��h�{�}��@"Uy�hC��t�\w���pZ��R�y*�bu��~���7� � @c�G��������9$�9�Q�u���`���;���1�N����
�o�.f��q�ZlTȆ.�>5�v?m�$�����d�s�_�`uO��0�8�9���X� ���П�T�ҡ�Y/�2���O���G�M�ڝ>p�Ԁ�IJΊ�� �/�-*�s.�F�:*��v���
YZ��M��*E>�U{�}4.�s<$\,�v�XΖ��HAp%)s0�.�t7���k�8�,�בH����¨իEM2\�^����zQ��s�SA��:�c���K<G7�Uu�o��+����8?�I��zJWs_�ʩo,�fbA婃�U�4���i�Ϭ[��)
5����xA��9?�,)QEP�h�Sp.������I��L�NE�	C���}G����J����=]��ux-�G�2���"��t��d��-������r�#���{�>�OfU\K�/�Ts�Шm�-j��y�_͆*��q�[���-��H2y/� =HՐ$D���ʅ�_! �ڕ}�g�R4?.�> �8�����^fY_#����2���̇6MU+�+��P�G�����04�a+���D�,�|�Y�.y���Р.O�F���y�V+�����+7i���ߢĆ�/D��S;��>�Ϛ�Q��X���$��0}�o�ˇ7"*���Ɠ�g�^�͏����J\~��
��~�t�և~�ی���nm�6Z� ��|�CY��}�����LR��;�N�Tė৐0�!}iY�&��4�^(�9����!iH�>�Y�#�Yx(��f>$7n�G�Kl�CFx�T.��mtWS������:u�l{؂�Z��.-�p�n��Jl��q�)
!b��f��w��䜤B5a��TdT�Ե����ctıt��r cW���t�"�!�34I���!dQV��>2G���=(��p�=<����^����眒��ϓ��r�K��]����)-�z��_��yV-�b�珗�4xwD*NN�8]��ܞCIN��1�VyL	ɲ����g/�Jp�Ct0�h��_�x�|t�g��L4{�����ܧ����K���/r9y��R_�M�7:����y)ͽ�F{(ô}���LM�n4҈3P�&5R��8#}Vgʾ�g�]f��OڬC�~s+<�ZǕ1�7h���H,�W 7��Xn���9���W^5W��G�0�s2��#�E����bc �ݶ홞2 *��E��S��-
;%�CZ0u`}�7��	�3lm� ]v�d��b�%^A:�5�V��ȼ7k��3x� �,��"U���Ga�>�u�'x���wIC�ݳbn{�]r��yg�0'h��ZK�_'"�%2~/�4�k7]7�� A�:��<�p�9Wf����w!��S
�j8��. 8�����\����Y� +k���0q.䬽��s��r �-��'�55�Z/[��$�l�-Fg�-8���H���p�-�!�-�1����A�5�.�F�g3�����e�s�x�R"⪭�U��?�XlB��?\�,U����[ue�*��d��J� �EB�&ڢ��?��Toc��V>�=��
�
�<������)gI$��0��H�}o�g\�e�����Y��� �|\����
���Sގ	��
�p��l�F�J�&c�ʃ�Ix��l@
��S��.��9-�Y�쁧 e�w`�u����7L�P�jcN�����"�񖩍�>m,�6,�0m]��X�fo�X��D?k���_�-t�C[���Ҵ+�{�|���ne�GxMVIp9v�F�W���C%W����z��<� �7������(-���P�)�:�
UN�WxJ���/T�;J��;S2`����9#��sb�Mt�8J�%T�!�U�&��M?�>�5�XT�� Z�̀HAӑ�;8�:I�p�Fս��奱ߺ7�aj��gu�n��5i�ߥ6w_��:NZb�1��h�Z�g�.�!(�_ޙ�x�٩��<aj��?��P<3S�f�[�d-NJB��a�N8�J�F�AF481�.�,�Q��ew���3O"u�?�Y:���D��N��)�3��q��wy�q�|<"r��=L�y��ۼ�(�4L{ kE��Q��-�fcz��U����Ov�
y9�X�� |�W��p=&�ø<�����pܓ����S|7��B�
(����@�����Q'H�!T���c�Џ[�iGX0���F�ͺb@	c�!ǥ^^R�c�e�h�f�]��>~�U��8�{��u��p9ǻ���l��M�vK��p����.[�8�1��N!j��4���;�:�IhB-�结,�����V@��k��i�{�rH�]��*qV~�6�*3�H��T$k�'��b?����x�f�#�pP0e:[�y'<��'&��l]ZS�/��>�Y�D�YM%^��D�E%�x�*ˤ��"&0|τ�q�ݦ4-ӕ�t�wi tڎk=L|eQ�)����c�ښ'!ZknH�XG���ϫ�t��4P߿�q��d�ck2�<�Vr���F�kG�A`�Yک�36u�@���ѕU§�zd*�qBa>���b���HPeR�B���~�c_=���K!q����6�\�\�n��"+'D$�@���q�Q|�|�^�Z{�jeu��L�#�({�އX<Z�0��t��|a����.)C�'vkjʎ�0��];�r+�A���6�MG�W�LI�{�Dف�72���ItCo�W���v3��@�E�:��7)^��˱�2F0p9�F9W&R��BxY�Ks(����;\�Y�^�?&BL��T$K���)4�g�q~�ɘ���M�����f��L�M��t��jo`!���vZ�4|=�	"�Ȼ=f.��<�v�R�bT�0��g���몵�zP�vQ	� �Qf�*���$���cA�?ڠ!�=��b���⭂`G,���:]���ʒ��}�ޠ_���e��b�:fP��*����L�W��"tʥ�8l9~#'�q������˄���,!1r�����?m�k�f��<���b9���F��,��!Df���]�x��ڽ��m��y���L�ٴ�U�����ꇣYѴ@@6D�˺8�]��� ��}z�������Ⱥد�^�x��w���"9e�5�ψ����o@��"t�K�xtJT��H�/�%Ⱥc�_>V�_ǽ�N����8�G��;ǥ���p!��r�$ܦ[��P���^)�i6�.2@�Tc�����r ̢�93��$��12��89��E�� �jw��gH������Z�J�s��֩��K&�p�?�<�l-��}���I�;w�@�ჳ���G���
�q���w3\ʖ�
eK�	E���K�M�B1���a�?���~J  �+��P���brt�u��b`Ŕ�o��Ϟ�mHS'�&w�q�yZ=�g��N�	�:nC����c�&�?������@�@m��R����%���iK�ۯ����O��	�U0�:�F��8� �IDi���1SRua|t����Dgoj���'�ׇ^����B����.��`�������8�ĕ�}D`z�� m�C�*L��̷��ʹg��X�j�!�����v�T�+�01��(ъm�~5[�q�U�l��T�
:�f���L$�����D�$#�ݽi����f���G4t�?�؃��Vc�n����Һ�<�_�[Ұ��s-��UF�Q�Py� �ȁSη@��4��h%��D���CX3���萦?ϓ� ����;I��g�d�k�.gUl����(���(�VXl����v�I��Œq�]1�|yO�ǔ����4Ai�ӟ7��-([�lׂd'ʖ�jb���Ԧ2���W��a��v�	�	�H�G�Y�l����Le�����mP7a'�6 ��V�{.,�FϷx=�'��z�܅rԀ��S��C:��іTKZ�لo��h�KU�jhq=n���պ�0Q&�J���e̡\��r2�o�?Kz�jlb�kʖ�Ϣ?ׇ�͹��L��0�+�Մ�)�e@<�T�>�4�vC����B EYNI��ԡ�Np�T#��[���V��j9�kK�,��Č�����Gx�:�%j%�+@�ɓG�s���ao~5��w��0c�P��O�Z�٪�z�4����*G�xn"r�.ڙF��-�� \�4>uN��=��=��"_�	=�A$W.iM�G ��]F+<:й 0�!��\ǲ�uć�]��T�q�3`+!X3���{��Eq�1:��U�q�~0��)El�`�/��Ð���Ӗ,x�Jx^��u��9�bA6#o�����d�"�8���_�%�ʀ�zڠՖ=�IykUsC���y�&Ӛ�Y�Qf�â2-��	(�qW�xa�lD�o��A�`�u|m��C�9�͝�6%$��_��Y�*��T |��?���h��̸���+m�˺�s�61z�3u�w��{�)��ѿ��[D�w=�T��t�M�< -�ِDJ[��Oi�V��\RP��)y֬��PP?w�::�6����n.��f�\5�W�8a��n�*�M��C�>��V�'"<��YpCT����lz��9���u�S
m@���`��y�-�o����{W�;b��f�E����Y���8G"���'Y ���������/)�4d�P�O�4�g��Z�\m�*N2d��\l�N#�CڥU���q�,`�ٜ�q����g����J����~�˗M�Q�k�)���ϲ�	!�A0͌�:6=W���1��1s�"K��B���ݮ8��alS���ia�<�\$�3m�i��Pc��(��ګGC����d�-�� ��2���-d��i�H�#pبj -H���)^0E�`�]�E���HI��JNz�kt��k!�و����wK��Tmݰ~S漯u�����(�Т�T��&�pGXj�~��WM\��m�6a6 6��z჊��)n�+6hW�A�̌�aD7��}�ˇ!ׅ�?�da �XfSc���x�!^���`�����n�yS'?k����/ ��[��(��AՑX�C%d�B�6ɴ������Gv܃����y��o�wqB��痵�:H3{1l�)p[�o5�j�����zd�E�牒4Ά��äL����2��:d7YҌ~�Og�3�0TA�����Z���;����q�8����/E��=��KjI0j��LL�{��ْ�eJ
�G�Ke��I���Pc@aB�4._��@��\1�G������� p����8���*9�U�n���^�<�o������_��yH�P �@����%�A��A8@̿q9�/��+�m�t�<���j|E�S gA�$
�jr�8�~39��$����6p(C�.5eg�Lkl��K��M'���믏�u�n1��T>Ct��Xl�������P�~FKά�ھ���<��+|��f���hj &��G2��zk�)������uk�A�Z4>MV*7Or���ʂ��е���w��.�3v�4 ܛ?E���������M.�A�K��D�:nW�Z����k	M�<�U�K3�N�
ј�>���G�4��T���몎��}3����C4���f#(nb���B��:_���/��;ess`�q_o�o��L������L��Ղ0�Y<fm�>�қ �:��@���tv��$Aɽlp�i�ʯc��]S"�ވ���qR�0ն����t�Y�K��Jƈ����e�M��3ޓ��i]�pĳ~Y�*4RB�+�gTI*S1
���_��O1gK���oD�jv����3?Q�?�	�|�O^����.�{���f��T��2�P�h��m+�f�-֮{S��L�_�$�d��q��Vo~St,P>�=A��ύ�_Cd� ����>�͍�#�ߟ��gE����2�Ɔ���El/cN����8Ǣ,���!�WO�'	ʉؕ�"[I�����9��}�Uo1zt�5�f�����k�>���ޱ�͒y����t�b���ư�'��0�Z�jhx�v�hD�&��T���]�O7�%M�����6D���'���{��Ӆ9�K��C���5j���̮�i�u>7��D��Ѯ[��1�NL6��/]��l�Ei�Q�Ko���-v����O��L<TԖ.�T$N�#������;<�M��s�2�6ʆ �D�KcSwxW��!˵���8=�\��6��C�ܥi`v8uߠ4��Hr;�@iy�,����8^F5����L��@I�*�FQ.pT�Ğ^�H���a��_������Z ������\9W�����.�*s�z����%�U���4N�x;w�a~������:�E�fl�}�\��0�z�4k�e��S�c*ۖ��X�L�G�1�/��6�j��$5��i"��@����,�?XW���ޮy>�~^I�<kă `�f�f����ʯ�}{O��쳊p�vk48���r� �|<���yq>-�bH��\��R�6�f3qX�pS�+���,M9!�	:B��Y�&AI�YȄW�E��l��X�,�|'6�k���R8�t�N��� �z	:�EDw�k�o�.FA�T�w"xlO ʉ6�,;�����R�F� �{�y�ez�uK"c�	�iTV�{:DA]�2n�X��b�{��.i����}~6�*g�jV`F�i��o�wG�^p�"�?�f�����M�R+��|�
�GZz�hBLk:{0
?ĉ�<L!l��e�*4l��`�:��v�	��k��D��X��L������g��ͩT�P���5�2 ?t��ݓ�"ӭ���6��L��]PM�?\�~����3��f�^H�)ɟљӻ�_cpp��֝%� I�U����2��8�xtP�]�B<_c�1�9��!���o�E���*L�C���&�1��"�@�,A'�Y!����{�wq���L��c�n���7ƍӫ��j*�!'�X�Y񝦓R�ّ�t}�c��,����gy����O�Os�4��a��W�4i����0d*���.X�Ro$2����ʫ"|�ü��`�-��HLq<	#�{q�Ir��:��G�G���H�w��5����P��oM��G�q�@�	y�j�"NŮrML<�'�A����E��5V�{'m�-Q6�7�˄^��F,5�c����~2�>��;���j���w��W���z�A��p,x�UE;�pa���W�╲��<=Z�7U��	P S�Uh��$��L�f5����쵹Rѧ��Jb_�9��I��a�m�@��R�ޅc-�J��<��$�~/rf��p��^���;3(A2�����,��bj��֦@ö'6�'��6YK��s�*?5DD�p����b��*K*�A��zU��[��KF:9(�#�n��3d��M��z�1�7����YC�=�����T���bE]l#���hw��u�ɷ����MLʘ�_b�=��1�Cń���XM�!���2�ų�a�J�6*�m���<�b��j#ը�S��|͖�ࠈm�g<�`YHaA���_�9��V��Pí,l��x:�eb\E�Ԗx%�F�z�w1N�>�,C�6{˂�1Ap2�|�'q��)��}��UR�p�l�amѝ�ؾ�NŹ	�_��ƬW�7^~� ��u�3	-%KJ��&�/}�=lS"\�1amr���l��ڌs�ЈJ?rO��])J��G�&��~�aE>(���e�{���Mlqt\F;o�~�Dٌ�ʑ���!Bb���0[o�wS%sÉR�K�_�p����+ӑ���}Ğ�t@j��y_c�T^1/���z8����qt���T٭)�+j��F�G��X���Ѓ{����=X�W�]���v*^�	�z�7�8����=���}0��ϥ� �}�H&�8���߿�Kd|!�ʹkF��O0d����b�bԳL��~ErߍᢒH�b3 ���F�%���֦Z�f��<��g���g0X���� I�� O=ƪ$��Y�̗��Xӿ$T(ԇי�L��Γ��%�m�'Ww�)�bD�E�7�&vZ}J�mئUW���GP"5#w�h��%a��/ZX�������t>L��iTcI�&?8�P��4�{;avVX��J{%䷌��e��H�;�`=�̜Vb����,�K|���#^�h�U��d6^���\Ղ`��
�>���5�'�Ğ�H1��
��&G�>��p�;3	E��~��N�"����@��5����^!��|W����sP�YB�*2�-g���Ų3�[G}V\n�j�n���+�w%�X��)�Dl���R:��r~�C�d���1Q���ľM�a���5�n4���%ɋ�J5�(���x��x����o�C5l�c[��n���2��_������ ].nB\]0����lI��0�Eɢ�Ζ��S�읂5���K��\aֶ����l���nY�qs����X�a2=NFatc~T�Tz��*��I*�-8jh.d��h1�?i�{����N�]�&�<�L��$b�g|���M�J!��-P�>�x�B'sH�sG� ��{�Yp���q���W���!ʍ�η���n��~ ۲�Cg�a�qA��h����y���V�݌mo�����_�t��w?�u0ӟ�h��.Ԏ_@�O�З;bء�� ���x�����G��>�u�wM����@6\SJ�-�/ȍ*�{����i�\��S�,��zbM�ײv��x�������:d��X;i��!��eVԜcLXP�>ES��n�O�G�أ������y�Ј̽l`��~��<2��@��+Ԑ��"��5!�;B��17�'Ymp�G!��SZ������8 ׃x�,��������-Dvfj�5�ɵ�� ��N>y�I?`Ʉ!����7��ж<z?^�����xL"H�C�[�Կ�	G �`;yvY�����N�3�y��5&BZ���Y΄6I�dk�����+�T%x]?���M�Z0��X��`��W�#3]�\M@��Q��跪$r��;�,�Ή˟�`��GV}8�����S�N9�Ќ�y�f c@PÍ]gM�8�!�1�ɻ��i�^Sz�w�A3���>��(�������D�Hr�]Miu2����1�J���#�y�j�GH�xM���68{��Z�m�P�W� &]���j$E�8��&|_f���*H��z޸�g�~ �&����Ơ��E6�D\>�K�Sp9��a,H$K<ԣ<1�_�`�-��.�'�?2>N0�N-�X��P�_f;������+VT�����V� NP���\n�o�V�mB�q@�i�����{�7��.�mc2�jv�H�Wľ��C���������te˭�YU�:��E�mkBݺm��l��{A���"2V��g�o��W��M,�i���Ӄ�	�R:F�0�@A���C���s>�ҋ��{7F��3$t�^X�A�˦u\�$s��ءk�@D��.md�${�Ú^��G���fH�"���|����8�_xD��׍�;�C���|�[�@�Vb�%{Pq�6~&
��A���)���u�X�Ng��nz@/Y`H�<np^����x���i#��Vh<r��"]�D�y����O��mنT�O���A������[]�/��xF�H�W�8c�v��se��K�&��0�L��.��6�.��H�"�m��m�����J'b����܇kX5'8Yc'T�/�O�=nU˘�s�
�5�$���l��ӆH��V���Pe��"�?"��w��s2R��[k�/Kރ}���k�y��7�>j�+�\��H>�F¯)��^p���:b��?-��)��=�=���F~`y��;��8G~&�g�n�AN��F#��2{��+?�k�,�ќ�[V���:�Ҥ0���Yt��n���d��B��ړ"\<���xAP��.��Y7�2�τ{o�*	��KЮ��Oq}OR�i��ɦ�;��"���� f���<���SjjIKm��4HM��
�uwт���0���W��v#�?� ��$R�͠�V?����;`Tl񆆃�JH���]����G2��M�ᥨQ���Z�Qf�'�`t�c���P���Ok+�u-�$�--�"Y�#����Pi��<��\��,E��7�opE�(�X1�F'_nv�������Q��()�tP�`�l<\eG��TÚ���6ʓ�K�[�*B?������,܍�1�5�pIOE���9���<YK��vj�p:���z�k���[%�GՍc��D����fo�t���cp�ȊO/���Y�ם�'\`��{HQY�&�y*�F�<-n�\��+G�F;G�
)hw,�k�8+Z&��>��V��~T�_��>���3��B�!�ec��m~U��Q�'�#.�X%^��pP2՚{T����P�ێ�����0�i_IC;s����ƒ?*�+s2�Rϼ��p���Ȕ|���ov�j����L_P-,�Y� R͎��E�U�����_�wD�R�'��	x����ٵ��_��'	#`�TQ�i��\ʍ1q�?闇��v柱�a�ʋz\���C@���
�����(���#f�\<.Լ3�Ġ�3|j�A���6 h	���v��z�Z�M�J��ʶ����i��d#��"� W"
j�z{='L�~v��,�V,ڲ3��ӗ}�:h�ɴb�d�!AcS��T+�U��4��R�F���N}���pJ`��;���.>���)��n��\oϸ5�4��B��B�����\Ȼj���=�pl�EXZj��4ʗ�> \�k�7TL�S�^$ֺˉ�ʡp�o?�{"��Q������T�GL��YCaR8O�Ҧtv�M�+[����q���Q��:[�1�`�HZ��q)]�LV7��#����qҞJ3N�v���p,17q�ܘ�X^��qRa9�^��Y���8��OT�$ӟQRv�g�<X�>��hӯ+0�G5jR�2�];X��pL�t**eM��	l¯�` VA@ՆAA|����o��w����Ь�@�9ex�A��oqI��5��Xz��v�B*c� I)I��c6��_��w��IĉQjf�\�8�;p�f�lÆ�ং$ɉ���6��Irm�/06��;��ւcCM�xz2&/\��<���,IGaF#�p� m��g��l���Ȯ����I�l�AH�W�`M��>j)6�f@ē�ڲ��y��3Q+���%�}ҷ�F�O Rx y�p��
�<'1�Yf7}$؞K��u��J����L��̴�/0�tm�Z��񴤚k}Fg�z��>�נ]mi����4%���V���;>��]���v.a^HVƩQ����}�*ɚ����g-D�m�iOme�4 .N�ս�}r��Uo�`GƟ7����p.'g8���� s _4(�(V]��<>'C�68��8�*��ظi������fM�>��D~�	�p�fws���z'���&�&h����H^���m����P��5E۹!�k*O��7`�}@��<���'��_#�*�)�_}�K��l#�W�ÇWc�0�eQc?�|��Hn�D(HU���P��'ʌv�ʫ^5{kjP&������Km���O�I*����.��VrdǣWg�h����a�D�xҔ�@p��X�_�B|�E�f�S*�d� �<F1m?*v�n��s���!BI�)~{M�,�v��c�	�L��%c	7��?҅}s�(�3W��F�,��~��"5�q{�T|듄�@fș�ua��mud��u^�D����ğw�ur���p�2�w�Q1�J���{D�8v�TN"�ܠBr�\��MIx��uM�~"�O�b5\�#mHL�k[p���R��f�g[\vZ�7����1�P�-'���!��Q��[��h�mW���>'f�����.]�e�
��ɣ�p񃋭��/ϹDiNy�1W숫�7]���ɼ��!�+�$~��$W�����yn9`���v=�E ���sM���R�+�\�+S����!����~�Mw�	� L,ɨ��[����y���ܭ�q�N-��P�d5�g��Bq�i��}�<4IWR ��W�)V������ѣ�2$:%��>��&����-W���Ջ�柨a3js�#����I�^�f����1�!��ɹ7Z�h����b"#Q���{�pb�A� p��Z��V�S!᳤���p@�����U����ˀ>��/n�̙�X�����L7^��9S ;�u] t��7:�c?�7�ry�����n|��4�zc��Y�*�XA-���s9�&[۵�4D��n��pѼ1v|XGKq(��,	�㾔���Dp<����^χf�@�#$�-3�yI�%&�.�?A�K�;���R�1�2�	f������k���a���^;Rvι?��
����v�a��'�˫|���/��9�E�I1}9|˴��N΃hS�!�6=V߾*�r���y�G!kj��ꬰx�;0*�h~P�S�-i92W���Rf����|��Q�ip�-%l���琝-����l��k ��1 xTZ9����vPq�aǏI�1*uuN"/�`t�f����O�8:�Cu�/L�+e\�Z��ÏWRjG���]�²����X��������n��l�7�1�xax~�c�5�X1"�!?%�l�zP
\��̄*���+�� G�r� �|bx�����z!+-x0��+���Æ��b˝Is�����'��U�tRos]�ՅH�-&������\܅)M���Y�ALg��+����~��s��� ۆ � eG���O�`�v{Ș�`�N�H��,���ߌv�e��c�psdJ߄�5�l���]�������oŴ`<���,��ݶ���oz~�8$kG#��#��t�> �y� �h���p9f!��$�`��qNd)v���{d����b}7�S�n� 1\.���8�^"��?�\�Ѧ�sM�ћ[�@.����;��I�K��;Q���@	ۖ��!�R��z����A����T��s��M����ynyRM�p���N�oyhds��;�$ �묺~$��S�50E���#��	\񵩉2��	ӹ=�.�	�����挑��L�r�d`��`�׍�b#pt�Y�&o�;������U��OVl���ص�v*,��:C~��2�(6Xj@˽.�F�'n�@�va���~����= 5��%�Ǽ�\2����b� �.Y�٠���g#�T���V^�82�����F�Ϙܸ���<��|�����7�(0�P���Wm1��
�SĽ:���R�V���O�q�Ud)&��-�C���j\F���ꇹ�F����y�f�κ{�N�x����q��|��Mc:��-�����e��r����(�2�P�ѢX��"��j4p �e�B3'b���	�4<��(�<��х�!/�Jg����IT������R(�
>�W�G�[��Es�J�2H�xRIdUa��8����*�@7�͉t`���n����K]r��
��[���\:��[)�.�J):���������qUGފ� ʅ��;@x��T����.$^�4꫻�_+��M�}N~ "40{���Ճz� � `-]ϵT0���n�0\3�j��c���vF�.�F%\s��r����l�vcp}���#�����g����8jJ�5��}��~������J������j�!�p���s����aN�Y7��-Q
.�	�����f�E�j|���՟�Z�O�')tt��A ���[�7��1�lb5+��~�x����s��z0 [h��
��	tVW��a��Ag�Ľ�9# ��غ6��b�ҳP�]')�����K��I?��	�5M���Y��v�P�����[Uߐ�����+c fU�OJ٣ �(tOV��oE�FU,�Y�k�Đ.zO>.iR�9� �I�����%/����yg�_�V!�[;tAvUp7���s��lb�Y�l�������y����w�vzy�/Z�E}A)Y���3��E�=TQ�z��<�.gFC9�(���w��"BV�%��NF�[y��Cڟ�L�X_)PD����r�w�!�q��8>���g]�ʾ�C8��M��8eě���*�$�ND.w�k%����+�����M�&�VT�����hNS(m������-g��`�2��M$�Z�ըΤ�Wy�.p���68��R���/����ZQ
$s��1 �P.{���B+r��̊.<�h0�7�px��o�3!c|�Q���D���(�&�|]��(Xj��E��8��2���ke]��@�$�0��ߠc��5T&=���$������>�^�Z/)+V��1�}�d���v֨�[l����{�k?RT�toB�����c�2B���_�6s�A.�P[&P.�S`�B	K+�+̈o)���p!��fo��Zv:Lm�_�&͟��_u�뛪��ƚ�p�m�N'@�u%[�,�|�p�x�
^��u-��ʌ��n���b�}6�1^ p�ǃ�'f�b毴�>�L������sQ6,�Kb�BʉE�E+!��I�g~ʐ�܅48���Yo?�w�/��&��I|�?�b� �2mw3�����[�mB�t�B�-w~�:� X�f� ��a���#�����c���6�cg��~�����r�l�H�e�Ul��RW �7�l)~"�v�Yug��~�o�����øE@��'��TH��Y���f���8�Ж-l�ڱ��[�ќ���&��7�%U�6����ǓuL���վF��\�U% ���ױ(���<���K�2�kT���F$�s;��*z����hf7�H5
�0
�Q��cW���\��B��a�^���Y���p��X1ω ��K���oC�V��j(�紒e�V���H�EJN�u�˻쯽��e���\j�@�<�[�G�ϡG��R�}�w���g*~�*qc3��#HL�}e�Ii��<��E�I�A����6�G�~�D���S)�����`?[���+	h.j�e���4{��T������פ��s���n��8�qǆ�-Ԕ��!�M��� ����Ҙ������d��i#��H�tz���Lז�f)�f�	��~ f�&��z>aX4S1<Y{o����R�e�ʎ}|;̟9C[B��{tΚ@�z2(̏�,_B<�S���qw��]�8q2���!���"�.��9�������,L�"�9�����^��Щ8�X� ��P�=":���"�'�����Ά�͔�������w;8."Op�.C�ռ	��it��a��T�E?�96#�5��bj�<��.$Dd���;���\}��A�;xS+V!��P\x�f�$_�p��G@��a�������PG�>�o�%�H͚��b��:���!#J�c@-���|E�a��#��$춵�U�̬�gÆ���n>>��m1�Z�YiA�0m�'Ƞ}�����Z� "e;�ǈN����D��ƅ��h��p����-4���O�L��6~�������*��S����`��7�_���ᖋL�!	��2P]\����sdzL��<OY��7v��z:�Ƨ���s/�7*���"�Q����5JN�h:A�^�ai2���G�ч����-�M�,�L��/��Ձ��B\:L�%�.#�5����oRo�����U�k_�����E��L��b��Ǳ�����c�$G%��J��Z'Y�7��G�Nj%��T��:n��6�=��46�g>�[�*�2/sm�n�,�}CA1�Vn����`t���j�&Ü�0uuF.�R��ّG7���o�U+�CrMo�E�Ǉﾍ1��vҳ�1�;t\}e��yd(�)(����գ|����5�t=xs�퐱z�z�d�bs}�J�S��Q����ql� �@a��f��Q�����0�-�����TY��1�fU�q���B�U9n).q�0�C�;�2K;3��i�^��bXA��S����O����<�K�Jm�,����-�ֳ�$\#D&#Wh�5'$�#�����V����I8�x8s�I��'��)�`�Ĭ(+���G�i�8�B���y�����a�*��1�'��ymoT"a9���EnƑ���$��F��=��?q���������Pt��D���C؃J��gG���^PG�u~�ïK���)Da�K�ł�.�]:���>�7޾�K&Uv�wSu�z�����&�Z����L��u��m���4d{��ڣ�g���DܘCż�-�2��X��?�,�,@o�A�]�'a�0��	�v�+�rC&�f6����;����,)6��sK���b(C
 J�F��W���-/~�ei�ˆ����z<n����۱
\~�;'�qE���k�YI�oY54���-�y$�<<���hd��k��C�o������N�џ��E����F��j]4�������D�
��~���Q��$���������2\��w����ly� ��D	��Gv��5H���
ڽ�.X߯Z���Wr����B�x5�L _�%�]�j�m��T����?�$�Yx~����;�I������gd�/L��]:�C��R�YM�^"F���BΊQ"�Ŗ��g�:/Ufc����?��TK��80����7W���T�U� |CKH=�5�7~ЬHX3
>��p����u��ꔧ��ic?N�o��*�`2����a��^�N�n n1�Dټd�z�M�[�$\�A���d&�2B��;�=�Gǎ�Z�eSs�zHe=|���HJ��9��Jg�Xw��.[�7;��L6Z�\�@�{eY~��S_���!�=Ѯ��sA�#�ߜ9��L���j�ϫ�	Rea��>�/:o`~�mS�+oU�Byh�ʵ��mi������|�5O�&P�����13T�����}6�t�93�5����q�1W5c�/����֥��%&oV�}�@� �m�i�^�ҦyYحB�C.̎��6��ۆz-_�c��0fJ͕���j^%���6�U���R{�uR3�fr���&��C3\"P�P�͟�[;���|_��3��cĥ8ҩ/̐ac����GY���l�-�b�)8�+P�c���� n��ĵ�.�ǉ��|t��0�g��;E�u5�B���=dv��g|���M�X�������o��.E�1�{6cÛ:W:*d��Sm�j7#<��>����_E=M�Yr�qQD{�CP�1��k��6�b}z,��l17��G0�,Ѥ���J]�4Yı�.�b���=XR��� #"�l��Q�"S|F0)bC�rtY@���<1�rsGR�wY����0<"�T����pK���l��87	n��N���z}Uf?Ps���bA$ {h��¾z�V���
�!�a��M!@y��dg\&����6��~�|;��m,�-P0h?
�M�<~�L��+�[�D�&��0�i=����s���j�{3葏��GT�����1��BKh��፭hU��0�G��V�~�}ÐuX�D��[���ge��r
�u������څ�8�ׄ�6��]�ڳf�ޚ&ҏ)&�ꀆ�,G��uJM���|��ی�JY1�Z+Ä�L2����gҋ���25
L��t���\e�c/��{"2X(jʷ�ϼ.�Llgw�;l7w
] Iq�Ywe������I�����}�z�kȳ�y��|��q��ܶ��ɤ}L~`p���b.��&9�.�g[h���f�< _5��cX��D� T(�,�����H`Q-7�Up0�	���˚�Ym� �V��}��i����#�ed��r���N�3�g�Z�N���sX?u�ܩ�p=<l��Ek��B�ε��҂�Ln:P#�G��n�]���|��|�ld��6)�X�c��Tf��r~_�b����j��~��j����	�}YE��v9��f�_=Q�#�y(�e�Ou>x2E��PzG��QA80���
����qY�8����N��D�9����������h�rQ�E��������c�҈@)��8)ۦ��Ͼ�S����@�LQ�E��[|gMvȵ��VS}�M}ǳFKhN/��=�4.�b��F%��� �3��d�G+u�꧗�^�U@/:`/�D�Q
���N�purVC1;�Z�Q״.0f���� U���	Q� E�[�/s��-��;Ľ������(�f�!�ޣ8��]�������dQĵ�7�	U9{�BD�(�d`l��B\�e���:伃x,^�]���#�H�X��;��]����s�+ߏ��9�j�G��Q�B}^8�䢟����B3�:9�X�-�z��g�����U%y=��ɐ��9P���N�حk�|i[���3�-���{ �ꡍ/�R���GW�w��(0�U��o�ٽ�4"���\���f�������C�ֿ>��K��:ؓ*찶m�u�MU.�
�TT��P��q[z\������vX����f���.98\Q�|�v��K|9���mF�"4�,�+MB"�*|�o�v��S�/?n�j>�]s�o|��G��f�G����c�oл�2;6F�y@3���a��L̢��w��Pstp2ڠ��>�l�� �<�^���0/(�ᝌ�_�|G�z`P�F�\vu�u�?�A�oZi�w���mR`9���a�5�q�-�ֺU��^qa<c'��Be'��x�IQ�g=V�	�h���M&gǰ�HcTڅ�^�e"OYҘ���D�wY���'�o8�R-UJFn��%ᄳx�����`�<�_�8� R��]���J�-�P�lK��2&l�̢}����2u���+ 3a��'��t�Ϯc-���H?��XR�$�}��?���M	�i�{g��x����x:Xg��5~�h8���9��W��+�w�k��ѧ|�9�	�(����\��Č��Ҹ|�e��\A��MU*�3�F���>�b�s
��T\�Fƭ��P��Ut^��Í���P0�8H��� Bt'%����E�QR��A�΁����.�J�7fL���W�`q���t��J? ����m�1i9�?�W(�����j�Mv��Gs��-��u#��;�����[gB9��m%��ޜ}�A�3Փ��X��������$���bY|9
�!�	"�ލ�������{8^.^����̢���zg�����p�ى
U$�S�ᶵ߅q�o���<>1��l7�7�:��\�1�{$b��,��kD��@ؚb}�/��&���D$����b��IX�P�+>D�Ҹw_l*'w�[������J��@�4����-�+2���V��b��O�y�2S���Zɷxo���_4��>����FO�/Zjf���ϝ��]�W���{�,=��DĦ��v�;+JC�t�І2�V�������F _�9?�M��R�
��-�p�r�C�y�_2�����Uq���ٔ��ew�qm�o�{�G4�e�R�&�A�A�� �/�U��d-ͥa�C���@Oq�G��g�D#!�xU���~��Ϝ�He����^��9.�1�p���OU���1�Z- �:�B]=�� �n8���E#���虻>�y2�vE�����i�J�l��bַA��V�%��rQo���V�sXu��Nڛm.|�dtD�4wl�ܩ�seq!��9��w����iУ�/1�����Z���n��?x+&-�d�!$�ʺNr)��L'���bZ�0d�0�x�V1����
����5�p��]��Ȥ�@�k!��3�y%��9 ;����������	�r���T��g�釡�%<Rʂx(oX�����F0�g�̫{���(!��@���LA*`r"[5��%~�F��[���f����qeZ( U-�֯uYǽ�Q���%��-dH�2m��:���-�6�+RC�M����%�����[�:�Ӏ����?놻8� ����ψ@������#mۗ._3OC����[�F݉�ȶ��t]������W�A���o���/�ԒK��A阜r7`eT�K��b%_ef�,_�+���V&��>F.�p��^w3UN���8��{�@�]��Q��v�(�Ä̀Gr��+�ũ,��2>�Vw1���D�{�J; �Tt#�g/�@�Lx\����_�@s0�4s��ӧl����[��?[Ԕ!Z�~6��(�t�_���E|�U�O�#~P�~O�m���3
�P��zޙ[�RC���YF��x�)2�tF����2�nt$�M�R E@Z�g� �UÓdtm6,|{Iگ��/,�a��~4%�UNJ�X���7V�r��%n���B�h��}V5j��Z���g"��O����Ƙ�	����Yi�K���J�EŞ��U�fܠ�B�����o-b��R�o��ٞ���XTg� ݐV���ʱ;�S,0��*��t�N��D�p�~�2��IV�Ѯ�
���Y=i R���` ����3;�˽N����'7��]�X��L��ރo�s�;��ٶ�m�i�q��SnƆ'+���t��:�T��3NC�+t���0PvV���"!��U0s�s���l�I���Q�^æ��`��)v����
}�**�Q������i4��*�ѵ��VUax#1�����r�.w��5��sH�XC�MP3�;�t$��u��t	q��H'��'�r.�����}Uۤ���D��Y��?�9��bf<��iq���D�$i&���q��;޹����5���&;���)��2���6�bb���fо$L��\��F��&�\�:P��J� ��Kcv3a��Z~��`��ėpS�ĺ�����Ȁ�������XK�`����ڥn͕v���e�Dl�8��C^�S�l�A�Nx�+�,���Wԡl�Z?Z�'d���/��6)�G��z(k&��-^��,nV�^�ES���5��N���(�$�u.C8�����5��Pw�������ޤ�|�iW�/t�p��pQ��5�P��`y��\�&�C�r����JL���9ꄇ4��I�j�^7�>:�����ᅿ{U�VH��A��+pA�:�Jf�A��6 豽�#�)`��6����`� ���K���Lp��Y�=�����"�
VN'�ٜ�����Q�pѮyjj�{3B���=�BkQp���,���%8��'; ~x���`#�� �������K��۪�1i�4�Z�촣4�^����gp���T]9�k��h�2 S�6��IZ�>xڴ�ⵠ_���Ώ��M0���άT��ʱ��6!��9�q��g\���%��;k.p'%>Ō���ѓ��� ԃ��NJ'DP��=|x�Ee�5ҫ�����|�>���� gKa$��,0����.Ɲ0~&8z!�ٱ�~�V�H��v� � ���~�i���ҩx��Բ���e�W:,�7�>$��u3������3�K�S�X��B�:��8���<�Y@�()���8E�����D>Hc������g��N���&���Ѳ��LGF?ʀY�a݇��f|��#'�R���)^�ܵ|I��m=���eDW�@�@)�ӮP=�o��%�@����EKq,7�ڋ<i=��H�[$�]���.N�8}���}�Fh#�?l�~qD��t2G�(�Uo�ɮ0̲M͎����>������ر�?�j��F����0㚥�u����'�j*�|�Vϲ�݁�Ϋb��@;yϒdgt����F9�����U��2�ke�a�>�h���0��&�SL�%,�A*F�����~�IGJ2:Q"f:�L�ƥL`�Mb�RE�r`m�N^���	,\�,��gd��oq!����'hs��^N���H�B���{�%P�Jb^ԭ��E���+��@�����fJ�IJ'p��-�Q�[��KLP	���
�^����WSʐ�t��'ـ^���S �˄���[z{p�	�S�H�FP�`�:�F]7K� PK�ЉqB�<��Q#ǚ�����&��o��)鮄
lJ����}#؊*�Q1�PD�}���M�%�!����/Dǌ�f���B��L��r�m��
��B~<�`����l��j������"�b�&3O�j��U����g@�WW:K��5R[b�Y1�a����Qx�����tL���f����*�>o�v=5qU`�5_-�ݲ����zj�T�6�`\֘����MGX<�X����X���b�"�5��Nx1/ �Z2(~=�V];,��F��Zʁ��z/�;*�5j���&��i0�)j�6���\ �W�O�n8�\�R��a��Ϭ���Ʈy+o�$h��g��2�[�#���/xD!maM�\T�����{������^!���4'RPT���q�b�F%D�b�4�N~A"��������$}Ƿ���B�X�8;�\�@?O�@��!+�`6�#�r�:�<��J�כU�z�d� X��3�н̇�Oo����R
���\�Is����F�LB�����&�n��b��T���T91q�;���x���ׂ�.h��M�m������*�'��YS���&6xl�!Ζ�n��ȕ>�1�{q�BM?1����L��o�ك&��1M?��@X���ҷ�n�Rd�c�|��6�
I�ń��N�x�<�����Er<�ҽ����I�Y��F
W����>͓�����4]�C�TU��ws5(��+�w���K���U��jH\�z7u(�� W\o1¡��g}"�`e�jO).���y��^Ŷ�H��������%�����>/s���bD�=��D����v�,�-�>�g�+'�r�h�Գk�.t^���*e��N��O,d�1��ߐ��9��Yɴ'k���O��d��{Rl�c ��?�]W���*��vJ^�P[Q�gư��G���Z�n���B����H!6H8Ks�{޻4�W��$����a�����L�>�s����N��1�.��$E��2q����ϊxt�Qĺ��AQ	]� Zr��X�;r����a���5�8���d�i��UF9W�fPC|�CS{�#{=-xP�J�Xr6�ª�b��z�ư�~dP��Ct�4[������x�Z��>	���;e�i�[Ĳ�(;Ln��?���4��,�A���m&֠��N����v��G��,X�)�U*Vՠhw�r�ù� |�^���t,��IV�3�wF�!���
<�*��şe�7�M9	�'��Ob|*&NS1� �M^���� ��j��F�*��Q�i�`u���4�)'���g[��F}EklCԦtz�C)�h�>���� ���n(��頛�}��A�n��%'JY�+��$ At�qZe�{���cy��:I�N�s�S�U
�0�4�w�ν2{;8���-�1��������+t�2W�$X��z8!�����ݵ X@-��]`��v������i:ںX��q��+Z���I�e�Q����!�r1[��H���^�g!^?��߭Z�",u�O6&���ȇ�K���L�_*����,6��<��6(���q����u����n������GZ��q���3�8ah&�\��r]@`1� �
���a���p�e�+J��	J~G�,Ƶ����a��W6X]�u:]H凕��)�/!�Ο�F������S`"��QF��qN3Lx�	�)���#O�"\rw��1��5'��b5�v�0^M)���B���r�5�&�{�6��)5@j��M�)0J1����W�{�TԽ{巍f��4�V�ͬ%��W��Μ�]§m��'q0^�v�@����%��h%��iP*lo��m��(	9����g�|e�(g��L��e�X4�WI���=�ԓ߉C4mdGąI����H�mǕg��Ǧa�=qK�~aj�2Tҟ���[�#?��`X�٫�=��&���+~�7;zg�_"K宗��iL}&8�.E�mp�坧+�G3�zDl���AMH�TĴ���Ǆ@6]u�#[!���0uQ�[��:�	�SI�	�;+�H8�5��xD�(�ASu�좢�?y�O@��NM�K��ny�� ��L��.OYw�(�諢���yK�Kg�#B��Q��N�&I�W����
d
�p��,X��	�_���u��?��\,�q3�ZȆ��r�)��n�)�~��鉅7aF�H�;-vT�3!� � *+�(�_ʹ(�h�����)"�!�,��OI��7kn��Y��Ǿ	�1#�?�©�A�-p8���(�#H��ȭ/T����(��L#K��j0¶]d�*!���� lV�/�6+
����:5�
�!Ŗ�i�1�k� ��#����ąV���gm']�����}}~����.E_n��`��4K�9����)0�,��=��01���T���M�_,�a?��i	�c5+˩sL�?>�c���p�Wu_�m��0�'r���Cr��Dr��,k��B�iW��t!�� +�>0�R&�92QhgtdDc�_�ll�l�6`���D�˧�x8�ȆV��:W"vc2�D�@�EϠ2)��C0�J��w��O-�P�ԑ������wv|z�{��J��Ө��~�}u�z@� ��9' -0g$�=H�<g��	5ғ�B�8ae/N(��J/��)��\��E�0�#�-���J'�Ӻ�B�C���Ch?v�ϴB��,?m�|����oz���k�_� NkO]}ܴӿA��V߳��ܐĕ>X��AgLɦ�h�+���G8E�����0*p��J��]���=Ckn�k��y݃�	�\0Tr�,��J$וT�|�����9m�t�wa�߁NC8��v*r9�ʮ?N�9Cn8t ���Jy_z�nS?�Р����H3>VE5K��E6�w�{���@�qP��n2���p�x��ޓ��tEpLy1�M�������fé�
ˇ����j�'F��A|����F�Y�|5wy���z�&lSs�@F��������=��V)hZ%Pd�	��]fO'�<'y�4g ���:�G��� �Y��^�U�'���e�:iʥFN�k�D�%�2��b�� ��G�AP��q����u&s��g����+��ڜ�e��?�+�	_OJI��߫���J�-[J��u��[��j�sM�`ļDX?����!#t	7˾d�F3����1|�k��"}|�X>r<&8+����
���
�K��C:�O����rѮe������-j�����ݬv��:#�`#|�׹8����WAq*�c؝�(D��CHL�O7�r��U�=o:��b�o?q���ە�򯫮sU0-yM���:U�A�Q:�Į�h-���di���t�A�PX:k8���O�^��3ɖD�L�0��w4L���:v�Z������vЌ%K��_zK�'��!��L�&��;â����@"w' �B��K�s��]�5 ^��Lb��K��ٖ��r�}�5{E�ҽ�r*�T�|�;m%*/�/8`g<��ř%a]ܝ�re4+)}ȇ8Nm�B���������g�\�K+u{1��;�t���D'G~(��s����0C�F������J�iG�8��]B[�݄Z�3�KAϻ؛U�8b�/.4w|��6�_@�J��s��� q☽���O	�1O����̫#ý�9�+�H'�2l�>y��}FӋ�	�P}(x.��O�$��s���ֹ��4�z���g%j��D�_=ַ�U��pe7c����"�L�꺖_4	�$H�B�d8�Q�*�)=')M�{,��*]a�b-9=t�mo.�sx�����!-��4���`7�lz �C��۰��8���n�]�)?�|`��H91͸C�n^S���8^���)Fb_��e/W'��%Y��,ʢ��cT��#� q��֝��Z�	�Є�[�+M��Р���,�����od��5��P�SH�^���bh!{QKؙ��Lv����cG�ư@0Wu�X���VNH��8��U�xk��:�ɂ�t.L�����w���\+���������ڴF\��_�0�j����E��m󏜭�� ����_w�rR�c����"�N{�?!��~��k67%t.�6a2ce�x�����\��vP�l�x��ya��+nR�-ȇ�>܃�[�2�/�4_�ɛ"�BG� �����G5�Ƭ�z����C<��U�a�g�s"��Pa}��x��J@���Z�E��#K�/�L?Z���C
ʸlR�+`aNH{��!c����͇rϑ6�OhP
�(�xN�ǣ��d���Xt�-� !�q׽�Z�n|�D�h �=.GM��6Vi�*@�<��Ժ�����v5�v�on�G�V]d*��Й���Q�&�5�g��2�A�(L��掜Jm(��1�r�1�I�c�kœX�E!���ށ�vq��8ݜ��ς��Ҥ��>C��c���3�����7V{��.��m *�d�y3Ƃ�
�Ԙ?����a||/ʯ�zȯ����/�q��X'S<$�(͖�⢳f�|£uO�d�y��#�2i|�?��O��[}ci�L�9�V��}h1�C�8d���C�r�sf��^�!�`��wgs��C�BμvB�ޤ����j_��~�}0�Ě"}������R/}�Hx��+&�?7�BT�.*y��<+��Y�]pd�{��j���V9[B�^�5�N��89^�w�ZA�䵫�!�\������A�����D��=*�<"k����kޥ�?h�E׳��3�`�����F�O���q�BI��@K��+�ҫEe��K�?9e$ƻ/E��u�c�i)*��6*�ia��m`��?T����H����������l�(���A�9����b����궸ּ*��]{(�
���S� ���'����L�!��Ւ�D�{�`?�6��ǗX���P�~@E�һ����/n���T~'?/ٴ��>[�M�`<*-�A�p]�/��r�+41_�����,���cD��h�.{�'��Bu�t�|�C.k+{�1a�!כ�Yw+7	�>�,t�%#_N�e]���A2"5g�'ƶ����]e#��K"�_=�ڎ��б4��%L'���j�L`�c��
�5gz�@6��A����K%l�9m\m��RƆ�\3���u�P�����o���)��[[-F�;:�~Z�����O�M�/2�b)��i[���P�b��7j�㤀����pz����m�t_��o7�>���g'F�e�o�����#5�HXP�1P�d\s�9�5>��O���u����V4Q�<W�R��6�_Y�PTw�|ϱ����7����)8"y��~�H�=��Ց�ȟ���$V��3O�j7��_��u���P��?�R��[ւ�z�ɭ��9��늼E�[�#jp!�ڏ˖`�^b�w&8Q���SI��������޽ȓ�� =v�,����0�� �|����>0���4�S,�5h��DZb8������qb9u-��$�@Vy������aN�Zf�P�\��{���$�5�@�b��Yb��OP�v�-���ϔSv�1iQJ���"�a�EQ���E� o���D�YpE�W9~V�^'`�[�b�P��,n4����a���������ɕ����РiU��yQW���ɒT]�L]\ @c֚y�0�V�ȕɵ/k�ӌ?a�B&��ܳ-�C�9x�m��A�Q�[Y�O"�Spq�u�R[wF#d���ܟ`��oq$F�v��#�wL=jƔ��.�"a^���yZ&���)ZjzT��K��6Y먚\�1(��_"^˺�9^�JJ;����%鱠>����8Pȩ��L�1�����������[{j%�����N�o�����Y6Xf�����c�W��ՠW�u���"WY1o\���Z���e�!���JF���4��VR�O[k�,��j�ح�����m���h����6�_��Cg=�ܒX[���� �RG��~?�x-桺JȊ��
��?�����l�5ĩ��+�'�n?�?	#yݔ?�"c�]t���;�e�Ӷ�����Ǌ7;G���1�>ej�9v�m�;�a�2��t*��,6��a?)�B9>��:x� �ٙ�\�s\p:v��X���t�y:�E�~��ȏ�x�'IS�߇�C(���y[u]���[��ӑ�9PᙝLp��U6��&�0�X�6��K~1 �p�S�%]0�(���}��|�c!1SXr�%	x�U�g ���X�nL�7u>.^�j��U��d�,Z�p&� `g��77�`;�(58���<ò��i��u�i�6�O������:����#�G,[��ll�3;h�>N����ՙ�,�W됴(pF��S�*O�B�3S����l�(0��V2yEp^��xW�J�ҝ���8J>B֞qѝ���3w��Xmt�@���?T�hY2�[ùN���|��͠*�o'����	eJ`�n5"�sk�]R
�G�{5C��ZA{0�Oܩ����i;�1��x�&�Հ|,D�����ɩ2��\�!���-E��Qk_2_Gv�ˣt10ӌ[�ɕ�N\_&0�R���z7�Z�:�(7���PS��͌�$r��F�Z�{֫�N�F�V�^kyl�y���� �0�Ջ[4��\��̮�Lt����*�:��,��Ib4���FBEӘ�oڶu�x�U��<@Z���PoUuϨ<w��)����;8UM�� �d��*5|�<�.�⹅=wSQ�,��A���=����5١LyJp���}ǚ���V���Щ����|��d��y'���Co,c'8�b8;