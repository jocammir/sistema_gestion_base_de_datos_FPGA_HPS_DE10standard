��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0���?E���!�L`����^
d^��,�䞌�b^���Fa��Rx�C�Ժ􋱘�1D(�zq��=n*�t12.�D�T�u��ǳ����?j�B�25��j�޶��-7T��|3WA�K�%t����T��)`*� /~���f>K2[~EwdBdZ#�#ki�hf+�zd�N�l�^��#�E~����m?�t�5r��g(b��������d_���(ʩj��h&H
�w��}���;�뀿&���@=�\�1y�K�q����%����i�^�`�:8�G%A�T�����9�_1��z�d�,6���n��æ�N���sjp� ��F�c�Q�b���p��LO�O��O׬�qy����w_���]R��N�l@�wH��[����]�aT���1Z��u�ny_��RגBV�4�a���l��q����<ܬ^��z��WC2<�m��h��9��$����"�"6�8�'��*�J��ק&�����L���j��Ki`��:��v_�\Y��-������<��/	��̓�0J׋�����0�&~�oG.IY��֢ޡ�{�i,��xa*�\@��ͪ$��	�ƨp*D<S��D?*���'��}����#ڴ$߭��@��1��S�yAВ\����<�F/��j�10˥�Yf�-N�er�B��ZDz\�h��1���HW���5�]��%q�=��w �E0��S_�摴tG̙��$��qe�����{� ��.�2U rw�§֗�լ�!�[;	�>z��s��j�L&��{qa���Tk�+S*,��H�<N/��3vɜ��(��%z/ 1T���Cc��)`�+H��I�.u�?V3B���`0�9���N�t=�D%�@�Syj>4�id�a�.l��N,�e�4]�o�>z��|������U��@�$�}Z��m��Rf�19���|��ȝ�(c���c��!���S� ��\���G>݁$�C|�e#o0�x�sEf�������ck�Iz�7�4Y��6 �u|&ڢ�|��ZJ�𡴳�h*���J�Faٮ)N�	H��w� <�E�F\(S�����<��q��y�'Rz���?\����~�-u�/�:�qy*�S@��Z���=�R�M��(a���i�T� �rR3z���E�̠�����uӠ�����u_D�A���ǰ��%�$�q�J���s����8|��h�ѹA�ø&�{�4ZIB]xЙ@���Ŋ��e���g����G���+�1��Z��W�j9�`�䧗&��$�-�DP���2�H<�+�C��;�����ӧb�%������u��:n7+]�▹���D�i���F�,�f����� ��t����Wv4��y(q�ۧ�tl;���|����5^a |#=����wJ�K�2+��5�U��@@PwΠ��{���@g�6Ʉ�6���$f3"�^�� �z��)��Y�զ�rx�l���-�V��'����∖��L~�~"���8o�$&hbz_��e�	�78B?ܪ��وѕUf�ToC1d�b�˔_]VEu���$��m��a�-y�ײ,�]ۃ#�@5���J��T!�6�_DEO?k�3<w쬲�o�W>��a�WA3evFm�7�Ɨ���QNm4%��R�J�Mk ��QN�?���� N3�ڭwK��=��%��"Kߒ�J��E��P�Z�+�ո3+R���Je|��z[��3Bծ�@�^Q���a߸��ע9�7Ye:)&0������	)�:�W�҇[ۅ��!�r�Dr�� �CA�������ѽ�F����Ɩ�u�&�:�-^|B5Hh��cD���oM�3L��&0%�Bd
Z����+I���Gݞ���rQ�uE��@\�"���wVy?��1���2I������<� ���7�����3����O5�w���k��f�Q���TӤl���BC���;d��Ɖ��5/�G�/��-%�pl�Ʈ_�����6�EHÌ���H>RB;�[�=�*�0;Ѽ