��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���jl�7�x�֫����_��aoY��?#��#�r�m�"R^F�(hb=��pt$��e[5�v� ��n{L�x����o�x�+@wM�ca冐堏����D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0�������ޅ��.��)�_��W=�j�f��Y�dB5&2���.z~��ҭG��7��TNj]�����
9���%�vs��[�P�Ӡ]DMs��I�/˾�[��տ��J��?����j5�~���ng��2��m�R^f�B�=W^��3OH�ݕ��YR�´��c�'�	��Ȃ�M��&٥$P($�*]f�6�4�"Pz�c@�dW������&��oײ�O��c��������xq��s
�IO���Ǥ�첫w�3B�C���/F}z.��V�,���B~{��lA�<�����8�5�B�c�N1�_rF$�c��4���:C�[/[�L��ܽб0,)-\��T���X-m���&�"
�I���*�����qI��m�I�t\�Ѹk�MՑ�� |f�y���4�h�֯ �8�Ug:���PG�a0��HSg�Z�V��a7ʲ7�X�~��9<m5jqnSUm�%��8Q�j�Y=Al��N�����U�e8�Oy�y�kr��W�ɾ����N1�s2(�(�}��i��M���k���{IN������]�8�+n+�$��/�l*���R����]�pQ��gP`%�^j�^��2��}���L��Y]��I��=� gKy=��7ֈ�������&߈כ�'~C�O���pQJY�8�x��1�m� �`jr��J���4Я¡�פ?3�Y��T�i���ʑ�_K�����2	��x��á`�U�9�ɜ�N>�u�k������װu���+��ע�3]/�.�p�������U�/�A7a�:"�W�c$�:'�K��X��U���������K*�n6������ĵ�A�+Z�#)�W�����g�2�.3��nV��>a��]��\��Xu�����5�q�ER/�}7�[��ś�����@��f{�A��H�F(b�M���ps)�@�w�LV�3��bX�)�����@),t9VYJ����l���X��z~���]+6 �8Q�X��A�T��h�Τn`��;G������(w{��&깪
���ϸ�F�������߂���o�s8���f�PR��e���ܙ��Z�M�y#>L�<���B��	�r�*5�W�Q��3�ب��/���c5G�N5�	��x������h+�Dҥ��|�/�FouT�!��-Bt
x^M4���7
��
���E/y����D<�3v��D3�A���gH���ߤMws��DQѩН��_� p���l��U[�ު6��wx?�B��}�t�Ur����U�X�9��fL�Ɋ��a�yFa���b���ྶ��F���B{�KЦ�g�?��N_F�B��.�`y����b��t;���݋o;��_͹�n�g&�������(:%������f��?��j�M~W����P����j�m�.[ ۘ������)��e�w��ظ��Xc>NP;��@�b�zY�:Ě�9��k�16��}��)��<Zǌ�����y�@iE�
��&�Vh�g��T���*�xsz���;N��p԰�q�RA���iȃ ��Z���$��@����f8/�>��� ���Ч����W0��%���7�U`/\�"G9h�j&���0 %v�M��>�a�a��5�����^Z+�k�R��ȤXr��E����<ȯՉ�G��g����R��\v&�e3��V������TH6Yt }r.�Y���Ӫq�������GRvƫ��d��T�Q���Ǭ�9�������ƭ��-��*���c��B���IO�4�ўP��2�V�~��ѡ���{���ɪ���!A�2�3[�V85"F�Q:���}��|�zP�_�}ϔ��
�tw>���;#���ON�~wǥ��i��� /JX�;E��?�k���5�s�iy����.s���8di����ʈ�6z��*��L��/���®g(	��ubu,J؛�Jkĳ%]t�.��;�
 ��~��}��0����.��?J=x�uJv�0�U� r�}S��wE��Uk��5Q@��1"%yģ��C�D�P�|bE,i~����aW6bǧ�tg8n�����Rf�Ă��\��	XrH�`0%%Y| ��"�i��\�t�b���[��k��x$`��I���c�+"SF4�{����4�Fo�m�5L7k��5��Ueg�R�������.��I�͓F�֒��5��_qE|�ۖ�r�Ԗ`^X֬��Z��˛m��o%�Uw���9ih���83��2�zm�{�|���i�dk+�{�Xi�>��H��q �YF�h�dm|2c��b%X��s��d��g,hM%Nt�f�����ܲ�2��+���T��P�87g�v}4�f������w,�=}o���x��)��m��]QNJDK�}��n���4��Z��-� ������}���"� �Q�K��hR����Y��G\��mU�;��$":��3��r3�0~~>F�O�֟R�1�qq����ijmA��j6�6=��Da�u�X	L	K=
u�*�.�vxN�wA]�&!=���K��W���Z���7��]3^�	̾#a��j�����5�zd䴳��LP3�{/hQE�;�-�P�ɹ��2]�if-4O��{��x(%o�6�b{�M�`ws|�#��̆��D�	%������4�!KK#
Bi"��Q�^ё�E�4������?�<�0�]�"J�4��:��S
���*��T`��
~>��0���3�U�c���EN�RҪ�m%�k�y(4��.ߎ�/�1k�|fF����4��,m�f&,���IL��c�SH�r]�����wi����㼓f���w������#:(&D��_��@t�S��ڄ�����C��e`�'��̀s��ɋ��=�ϝ�m 4o3�.�ۜ�=���h9���{���4�fu��������,��R���EL"͉h\��x���
/ߛ���Zz�[���@u~�n�HϮ�}+�x���{�?��/l}vK������ßW����
�炟n�N�"�A��μ��Kt�,\͖(�Y�L��<J��tD^k�B�@Y��b?5^��-F"'���-��ˣy6\�jsB�Ua�2��7��[�_4.W`��N�g�����G��ޗ,�/��Shq;ʀ�H����í�y���>d�������㏎����3�~�@�R©������)�s��N�vG6�a'CM�Em}��'&2��O;l���B�*�(1;�C3F.�� ��1s�D�Z1<ݹduiȀ��kŠan1��W��Y�pC���W���Dv�G %�|`���M�z�[�_�ޓ�Z�e�BFG��U	�k4M��3r�Ĥ��aN[��r��pS�,�P�_=���4��9 &��OK�U�eE$�В
鷂�N:h:��֝��N���N�b)K���h��P���Ĕt�x�� ����A{�v�� �ܤ�n�����
L>U��O�rw�/Z�i�j{�3�-�1fl��W*�ˣ�3�b���6@#;�>�j"�J���9�O��trcKp^�V��S{ᕰ(TY݇r8e��kBh�/��-l���
[���L-�e�t{��BG�x��.�!�0EdmM�u��3�X]���HP5Ƀ�9���Hwm
k��f����� Ju��
w�ሡq��59:F&�:c+�`nO���`G�z`�B�z+��������L��>�!5cV��7`{W�t]� `����m�5���w댖��ͷ��O�������є��0�sj�����9���Y)��YN����6d��v����;y��" vDڢ;�X ��#M�lK��_����??�VT=��#���ڻ)�uSX}�[g�'�� �0\��U��PU�A����#�EK�7��"���'t8�UB��?��l#�ڠ�5j�u��_WR��:0��c�^B���֚~9�[la�"�P�/��X�Tda�t�I3�R�X��ݴL��:Wc��a��X�������?Z��n��ŵ{k��x7*�&K(�y7ɯ�&N��ͮ��~�x��(0�(&�(��4#B�-�.�������%���r��+�\�C.I�Z��J�� �<�g����m��+ؖ�J�$�o�H��(���4��W7����s�d|��{7i�VNo��lA�v#j�p����#�J�������'C���O�ۛ?"#�bw�����pP�'�j�B;�M��^jQ\-�L���^����*ge���M�&5�+ը�����q� ��?���}��L^5~�6�e�CG<W� M�U�t��u?���8/a�� A��jߗTƩE�%��Db;6��a�}�dt���$B�H��}��hzC��=�	�����]<l�����=g�㊌���F�n�.�}������-13�MO�멮��+��{�Z�� ,\�R�n푽5ȯɧ.MA1&���^��Rϸ�jX�y3�N.M8�+����(�\�.L=��&�~B��Q��� ��Ԫ�}
�����uy0�Oe1��1[���m�.1��(�Ր;.�0�A�5�r��xW��VH�1��;�!@f/t+#��O#9h����	��N'�HX,��N	��E�$C�{���推1�3�28������aJG�)�"��,�ܾ�����a\�©� 
q��U�b�>9��w��#��H���
u��=[	]$Xb���%3
%���7���*r�c��bg1���2�w�A>�7/���Z ���i��[K�7���,�4n��1�W�;%���_?;8�@qK�-rfl���<�Mki �C����pȻ�;PI
a��-�X�<QJ�&���.&s��yqkU5!X�6丕�F�C0��G� 
qKќ�hDr*^7E�$�çp�e��w���9��*: �/d<E�L;����>�N� I�l%F����G�[$��8���E,MG�9D`r���E"��}��w�Е���D*eQu:�1)_;�͛1�A�$`��H��y����t<i��l��.�\JT��f���"�c��+`���z6:�,��ܣ\�f���M1Pt�� ��#DW۟�؋�_=QK�Y��{,��'`r�#�(!�����ʉ ��5��S�٩Sw�;�݂�f;H��(�k����<i�9}�$ɭU�m�+K�n(�ϰ�_�0�d���a���vvl�6ᝰ�&(�K��]����u(��Q��I�O���b����(�|�����<�q�3-��Ly��Dѥ(�ݓN�/�i۾��B�����#�HX�Q8v8��u X6 �eK����S�h=� y�?�h�\�|�E3m�����5<􃰁�jQ����%lA�m�&�fyۺ�F��� : ��������E���H�=�4�u����6��䏋"/��\�^����7)��	�J�`]CCT�G6�r ?��KZ[�%%KۡW,A�'k]����{�h5h�]l`"�p�F+]���k6�{��]F%2�L��s�[���v��-u/FFz�ăKSIҖ<{wP�*�ρ&���،Gd4���f���AU#� �l'���*�0U��ؙ��A����)F����\l.�n59�>���d��
?��Q�ag���Bn@�(��TQ��X���ݭ��z���)8���;��Y}9N��LQ�>'=�f���v�2>~��޻%�i�\�rf;�`:��fCH��'@��7��;^>Չ.:�=�N�F^L���oT���ۤ�rzW������K��V�3Y&���\e���6MM��.��3]�� �C����J	�ӥ��L�{�W� I�X�$pb��q��t�e�a�?biph��N�|��Sc�� �r�w�X��ɀg�%z�q����S�+#�#�:4��NW�Ɨ}k��3����}DbGo�  E����H@�j|{~�q�N�ƀ�!�L
2��2.��E�O��[!�Q�z��9�W�앦��mF�8*=ׄR��}�K�[+�j%L��c�	�qq�g��５:g���ױ�2���ѳ<&������J��o(0[�I�#@��FO]F]�p3��o��i
U$h��|1�MWp�5*�Y}�l����^����ʯ�"�����}�"���	+c��+��|�Da7 ޺�Y���TjɃ�i֚H#�V� ��K�����.g?��d�F��est���Ĭ�l��t���}��m�-����(�ʀ�fJ�9�@�]N�� �VQ��mE��:,r�����}拊m��q�>U�5\�ǌ���z�j���vjڙ�G2��6ۃ�/4�e��Ƌ���k�戹Q�H֬m�,�93wEģ3��R����$� z�u�� �dS0|�K���QY��v}�*Qj'�C׌����W�,��ٙ�9��EF�s��ǚD�U����V]�;4G."�E��}Z�����HLx(�n�0�X��od��.s�'�ۤ��"��s�e"�s�<�<��C��U���a毢��%O��"R����ѩ6H�Z�n��hK s�.��O�� �A,���F@�ʵ/���]Ѱ�o-��h��y_������f��sZhY�{��*�Øs�ݰ��{F襦�ˊ����?>ǩR�����z�D?������?7w�P�e��|�<�c��bnd�´ke*���'���8�/��B����q|~��X�u7�����펑�A��FV���r%��ub�>������o.9s�@#�[EHTj�r�@C��R�Q�Q�O{FLӪQ%+�QZ�D�l���������,��E��⏐>��2��൘�㓐ݡ``F�'��ʽQ!��/tg'o� ��uO�h6�YH5��?b�OU�?L�2�0!9��?��-����g��AVƂ��,
,Ґ&�[�V�\}�ci_|E��C8���^=Y%���ߢq��(�	~6�2���w�a�7Ct��'���x�VІ�tEz�|��vq�?���d�(eŲe��qճ���RS| �z�U�A�>�b��}$�KK��D�W�kHs�C.�ֽ+`�˚>�	�]�M�t��B�UA':���A*�&�?��~VeZs�m˸ƂeV�J�Gg�4q��T�Qջj��v����NN��+���䔐���lL�
� �H �Bp����yrh�ЄBSg_�h�������\�n�o�NkZ{�h�NU��>|a��3%�>N�t����.�b�}6JQ�AF����B�~9v��R%�aI�+��i'���\�Q�7)Dݖ�.�ͻ���)��D�q�I�(^���Kp���盷l��艼�k�T�޻-U'���& ���vZ�x�P\ѡ��80���$����CG����!���&�̪W�f�{�=S9"]X\�Wv��Q�"�`,��q���S���ʜ�q��z�kBg��˯a����ɏ8���1�J�Q�I1�J���/>|��$ٴ%���9����-h,]�05u_\���{��%�M���э����h��+�oSkqj�>|���Z�p_U��1Ϗ����ލF�p�ye��s�3��:������ՈN�Ęr�Ir�J��u�]���=�dG7�lY�����&�̤��cH��@�Ue��R�m�������n0�m ��[[z��������wQ`�x:�G���B�9l���r�py�@�ӄ������L�؍�n����	KU�c��$6=�3���6�C�	i���iiܦ
�#�T��sW,^��ޢ�)��An��u��7�?����(U<5O���٤����bz
�q�#	F��v~�-+����!��g�7""L(*a���<���w�%k�u��t3�l�~o\�)�'���f���Ԫ�[w���f���"5F�p��:M+��<���Q9A�៹s��8׼�m��Bu���P�Xx�¦f؆�!��;H�4چ�c��n��Zt\%;h;�������tV9g��k(��]<H�L[9�Cp�j4E-�(�T.a��)��et�ׯ�Tex�ߎqܹ �R�23��/)`n]fK���8Tp{�\I��V`����膪�3���sD�E�L�=� Ԏ�{?��7��P<��+�-_���}���s[M����o����{���eZsk�}��f��xU+h�ߠ儓4F�W�~E�`�7UF������~З	�w<v�ۿ>XIW�z�r�1}�U�x>h��Q?���P��N�L�FZki�)5\R����Ř�a8G��š ,�[�G�B�kk4��~����
�CRF��x3<b�j�gO$�Э҅��;X_�T�]p�)�� ��P*���K�E�_k�)yb%jZ��N�4���^]�'`�BV����g�'�7p;�'☋����4Ƌ�>3�}:������n�w*m��z3� i�%tj(�ԧ>t�UP�|Y��+͘ |Va�(�S��q�(�'}M��=��)W9�8�~GG��O@��Z��>���j�<��joQb^�rmÃ�fŝc��c��#��C�L^(��1��
.��D�Lq��8x�6"��#��cry��d+e^�NB32�ǭ,���e�ڰ�]Q��d/c$��������#�OҚI{ho������$�R��i�7�ע�v~�:rt��'��8C�7�Og�2gD �ob�=#4�[ "�:�<�4��,�ě?��pނ6��[��;�_M\�M�Zɻ�E�0�w�u�Ʌ�l7h�L�OD�Yܨ����g����n�j�mS�}g+����@�4�Y��f{�7#��/n�~{�L^�( !�m�}%���4���Og�:~��f�&rk���bc0ea#ƎN��zNb\��o��]�t!�Tk��n( ��@��j��lc���o7rO�|U$��<��c:���f�%�H�DM[=�<���
>��r~Hp:�t��T�%��:ٛ�����$���gmq��PF�Zff��F�!�!��6��/��ʠ��ů:ܿd�c�5&IHŰ{4N�ϗ"�P���<�ِ��8/�G��%gs̸���M��uշ�f�W|��g܀�*;e��d��4w���Ev�O���3)�wQ�q�Kj�,Q����2�YU5�J��Eh~�g���XɁ���O���hߕ�{���0�C�Rʀc�{�.�ErpN��hAࠃf$�M�Wk�h��@̮��½%�>�$7�?�������+g޷=ȼ���[(։u<��l���[��K��3�j���e�q|��t�K�;���w�&�8Xr2[+���[��p�5U>������&\���.�Q7[;�9��l���]������-��:���r/\��k!m��ʉ�(sc�A���{V]| ڒ�X�RY?`H���ng�D괞�IL�"����T"�,��j5]�ʁ�V� _�bP8���M�%*oWR�I�%T
:Ӭ�Ѱ���F\��鶿�:DW�fR|mf�Gb���5�y�����I`!V���T��<�Kq)ڜ)�����9%ӳ��䳹&�6R������s��ƹڻG���΅�����<��[߰�[��lD�4��ݜ�T>����_9�h!�+f�!�9?����aa-�}ҿ�N�o�0+�"*�6*꡵�� r����N�8�Lp�	��8@X�rĆ5 �H�Vo�]s�t�����y�N��x�8t^�,~B�+�t �A�y�s?́��6���2r�l�� ���o�.R{�Zv�M���'�Ջ�r��@�jZHȽ�j9d:s~�>��hz,5���9�����ǸP�%�H�JPa��U���ќ����z��@���M�G�֕����J���Po�0��U���pPC5�q3�沦� >{�T�Y��jS�n⻔��/Yƾ=���{��'l�p�s����a�n`��7�v�f=|{e�[Ǿ�+3��L�-��s��1�3N�#��\9kT�v\
��6taP��\a�h�ނwZ��7>#���v��f��`)���w�E�)�rgX�U y�s�3,B���k��
��|�0;%Z��ͪ�Ps��I�Ý���ݒ�Y�:��CU!���q�.BpD9�hW� s͉_'�o���3�ǉ���O������#�4a>iI	4jD����8��z�25�]�(^�-0-���+�u f�&�����Jm9�g�����V+Y7��6�B'u����N	���z,=1���T_�t�E������ ��-�`�U���v��v*��m����O��7F���H	��\$��id6t�\I��0��{�,)8�]}$���z����z�|q���*9mCXQ��7��T��d�*����TEUvY�� ņ�|��<)���'u�u�|k��f٣��4t��VT�k*�ѭ��=��
����z�عV�{W��b6�w�V��p38Ң�.�ڝ�MM�o+';"w���#��Fz;���R�i������H�D>��@���Z[g�'k5����%L�.�av賉�,�?�=��C��r�&-��*�:�����A�]�DvjS�<�fC������מ"!�/��8b�2i6���@p?KP� l�T�|�b}��q*ڠ��r��A���|��+ҫ�v���T�c��'1�+i�`�F�$A��a]m_<�0J"E���$f풂���E�@�
�. ��!���{�(w�rL�Q��Gl�gIN����Vx����V���G��,��?�s���B�2?<���GO	��`�v���ۖ\x�6������i�'qe�7�����?K螀İ$:��=�*�����S*�4{�_�n�P�iK
�嘱���ha��)��*�tKB�gJ	����I��8���S�j �nn�z�*؇)��Ɲٛ�`Q�g�\Uы}�hP��T$~�X\��~^��r�j�fFEr�:}�۳vI�����w��%�����V��b�+�}���f �2$6�'��N�vĊ�(�[��虔�T�˭
��Ps�s�Di$�Gu��b��J�q�R�k�%���[;����6�����%&����^�c5U"$���Xx����S��$�q�^gU�R4s��#���
�M��;k8�!_�ӑ��c�'	�(�o"jXr����z�>�M6���jބ��sfVѰkű@`9�9�X瘝j^0~�֊��'{	��E�'���8�"k:�l�~�&�������B[,_@��A�RԄ����/M�1(p�N��8�	VC��A.�-5z��9���%b"��B�
���~�z���l\�;\s�z�̱��KIq��K�뽑�ȶ��_�����Mt���C�TҁN�ݐ��r��̮�jK��J� >���)�WA��1Rj�9��>�����N�K�`�!')������-}�dJmF�7Wz/�~�֓f���~���8�!L� *�x�����^��ePP\7�"v�%	��튘�f4�΋ ��fh,�ce/�T�{�ƨnM�c���eݝچS���ڬ�ߕ'+r\阸�͹�������ߴ~�
��jw��s�jWY+g�Sᔀ�߹�σf����l��]�t����Q~�*�t�`D��Wp����D�f.?��OL�^ �,Y�cIfk�RTM�p}4�O>�л�lS���z�!1��mv� �mt�t����5	Vl��,Av�ѭ0��a4ݭ��R�� ����ĳ�,������1�?c��>����O��+ed9����~��f��L"��� ��҃����0�+0����"ΔMD]���ʕ2�s�A��ľ:����j�ȾƋ����bJ	��y
;N"ҦNGU1�'P���B��nJ8�Gg�Y'��\�^@#43�Ҩz?���&�#.�~]ڋ�W���ޣs8/ņ��$\��Y$��|LDq��Y-��!��P�G�D���[���'�˛��N��u,��N0�o� �Q
��l̗�������S�M�����V����U�P��O4�Mk�!^���8AxP���2'Ex5cn����-���X�6�28H��ZS|K=w�c�6�m��p�*�2��k?�M�BBffN��gG��;���w���m��n��~Ƙ��V����:��j[�vU�BG��Lp�r��%Q�[w-^��������Q�̇��ƒs�*�k�i�<��gJ��>������&P�Z��W{�{�{;x����B;������G�B��0~m�4'�%�ß���}���w07�0����2���RJ$iH�2O�kL[xƮ��&��S`�Jh�DB]<�%9ዒD��>�)�X��|�64aG�ؼVߍc��v�����Yh�]�E�D�A�:jW��B�~)L�6B�����mF0�w�iD�����|�=�d(�"�#�9}F����=�P�^A����j��dU���e�	r'�8M,v����T��B�ܐo�/�مP/�`�L�/6����������d�vN�%�R������BM��vF�\fM�?�򍋒��P�&5�����O�1 ���Ei�g��@���'�1�x�-$�rb��)Zh��M��U�Ɠ�n-/�����%/���ְ)/Q!8��}��E��3g1���7��U����D*>�J���+�E�h9�؉j�u$�f�$âE��)�Q"=٪]�p�
��m�:I�P���$R��Z��E��,Ĝ{M�HOz[ظ���`��r;	��5�������c��\��c�#�}ĀQ-�1ӾIY�Ʌ��YY���44!m�^��� ʥ8� ��D��_��t6�ND�d��I9�D������a�O�UF��?�`�*�/m�*�9�: �� r� ��ym���2�RR<�SZ���f/Wj��%7F�vK;�g���|â�n"��.��Y��+7'oJ�VQ?��.����2��������Q��sξA��^�9.�.��4Щdr���`��x�
V�:{ВIEF��ZF���bu�(T���8�C�����d�x����=0�<)��.l^�!�d�
`�l�T�� yO���=_�e� ��n��}�]�"ˬx��_�!��?O����r���\���r�o%����� e/�殟�2R�CL/?�q���1�n7�a�0�`�G���v�*�K��%	�f~��S��~h�XcK:��	1��oP�qa<�p�P�Q�"L�oddI�'������γ�`i�/>*eRn�^�'��n@��ƺG��L!̅-��S��ow2��_/��1��"C�C#�p�]��ћ9^��(�`�Ui��.t�ǜSL��T�ӯ��)1���`�)30&D9�Ő�)�߬|x8E:cw���4��=��Yc���pa�x�����~
���6aۋ�4z�G(n���?f��9���z��	 �����~1O	6�P�Aof*�'���~��	��@�уV<�"��Q]��N:�E��ÁG���}��f�aq�>^��'��D�]����v=<U������HSf���������b��bʌy FC�ُ�]�S��l����Ȫ��#lއ�l�+�ɖ��>|!���Z$�����8�M��k��f�W2�v��CZo���Cݐ �c\�J[+R��Rnk�����pH��1	����֒�V&X|�\<)߆�?,+�����z���5���F���k����#������U#��%��p_X�S!�sU�]S�"pU��\\Ơ|�H��53�S��p�k��"yrk9b(2�֎
/qpL�h(3�A���W��y�q���C�M�V�F�@J
_��Yr]��0�͗��~��6$�!)�׸Nf�J�2#8
I��4BÑ�pwfS���:�DgX�vǟ���>��,����FsEa>M�C�(���4����\���޷ں���!��c�y!��=O���.
����F�kkj�Yt�%a����>���5�����E�@t�B��$<��4�@kwq�s	���ܯ��6w"�
J�~��� �L����mT���Oҥ��Max�4Kx��̄4���+�:�H��4h4
'	��AF6�Ūc���]�U�KT�
 �x�ij�EH�������vC�f{#����g�H�(��3+W]I���	2�旻'�e�|����¤�9ЍtuJ�p�bV��riڦ�A�?)�|wt��J�l�����_<�U�n�`�PXc�i|Y"z���=��]�:<��#�5Zޅ3,~<&�b2��Z:��"�G�SL�?���=����9�1ۥo}�{�
�6��U]8���C�P��ț��(�d��Ju}�Ε2P���سp����_�B��:���!N�C�Eω�K����~��d�
�E�\F��#�&CF��4:AՓ���N�*ؑ�MEA
:����������P�vp��?����82��[���n���[n;�x%���N�Τ�uO����F�>R�4%=�B$�>��zlk��o��e��eS+�Y>V
�ǔ�#؇��m	�fEpa���?4^�"-�����Wm�'\��ˤG��_����9���멈�qɛ��P�?Uo�$��'w��P�N�{_�oC��jJ^ܵ����ጫ�tgo�U��.�|��J�dci�ys"�~�>���������]�gUA$<5��޹��Yrm���j\<�z�|�R월 �X�Z��W��TK̬!WWlD��Z+!!��g'�K��^���RP�ݞ[��4�l��5�&A'����^7։���{6������M!z��X�E�<$�~���6(�ݑ���@����n�P��16K/5מŭ�'mD2�����šh��(U(�P*��]&�X�q�`��'�E6���	z�φd(��%�8q3Hf�zG����1-�ش)]}���h�$�R'1�TL�oRrD�z�A��@R�\�4�ag��7r��"�"�۽�A�Ww��d:%����XH"�o<���#����#^H��b�%�<m���Y���w�֙��J�9x)U���H�^zk'5�cN)4�u�y_�ӕw��Ph���tes.\�["!�	ߔ6����Mr��װ`�}2n���R�S�/�B/i�@�x�=֯ļJK$���'33�,�Z��}�іtӞ�;{�ͭ$��3.�!�Y陠-�TȨ$�t>������F��fکO�3�`U.�����x��%�Q.|p5��	��Jl��5rF�[�S+�o;����a.e&,�4�A1�8��g-�U2�T�}��Vk�������I�l|�u��w�,x�_�'�Зp�9�3���*Q���ĪY��+�֦��CT1���|��=����o�z�?����%cHqK�	b�_��^d+�,�YX���O�u��~�Q�E��#ͽ6(
3����٘ު�ե;l!k� z��	'#�-��?��1EL$H��m��-���C�G���]W�v7�!��>#����q`�B�?n��σq��I��!�9Ȓ�ba"�Erx~x����C���Cs
�8|*�w6�c@�9*�Ne�d�v�N�$�E�b;?�}5��?���Q���b5\��֋�U����.Z מ!�@�������v_����������2bfF���a�Y�1��T�G���#�2OY<�p���1R.�y�~�>����+��N�:P�Ҳ� Y�h�g�y���gmpL<���r���|? �ΐ�,� �j�g�.̞Ȭ2��穮<�<��ע}XڅC���}P.���
�_��=�P���
�l��c|x���@�MG{Y��ț%�H|�<��h�	��g���':�TI����m;G�V��.��i�QXi��y�����cj�A`	l�����f��G��Ź�+�Rt��*:
0�q���#�<P��%����r �D$����y(�v��J����O���������6'��1��X\(�#��E���h�/��Éǌ�}�<}���U+]�Ly _k%a�m����Tåu�Gv7M�;w�̨�k�����L��S�/�ǤG��Ш��=h�c�$��[�d}�_�M�������¿�����7m���r�C'�Y�����^�l��N�)�%��؍�S����B�1/�l�:�6�|	��Ӝ�99'��?��%��v<�17��r�.�UG�ӣ���4��	m�3L�8��		��?��˪���K��ȡ�6I�I�'�q���[��P"�����sR��@����~2�1ں"Hhk�6 �=�����g����Lb��~��,2ت������Y�$e~2�;R� פ3����K�k �f�xgH�
�]1k��Vt�hI�����3�����#����<�Q��|�t;�p��~Hyu�􌼫c����� ;Jw�|�^S�u�5���B^ ���5����LsJ��4�9���70���~"���
OǤ��%[̡cM8r����겆m��(a�Ȃn45'���w7�&�;-���5_�}��50:9�;����2�x<����w�_�'r��N*g�J�VXC��LY���4�`���c�,�C�k���{�H�l�:��/e�
��7����X&�}���OZc|4q�s�zV��W�\F��@_\�oj~���<;�izՎ,�#����յ�Qэ!)y���T� �K�:��E
�m����o�̕(���]��e���LQ��s���������['�7�#�P�r|�W���O3�}���G���,������O�Q�H�oAej��E>��E�{y/xC��f8������T��ű���n�E�5a����)LR���B/b��S)}�O�:)�L����̫��rn������I�O���
�U�����-�"�t�Z�dhbf�<�8�!����3�T	��0�J|�K;�}�G�f9��g��s���L��t_B۠f�OJ���a�;z���=�&�e������B����{�0��DSF˪-�k��~E�PoԌ�Ni;*��
2�¶�

����b�'�m��
a���5T�ì`3i��tO�b�b�q�l·O�>�N0��]"�N�ٚ�/x��np�fՈ��3W9�^���	��'l�V��G��r�K�l^�ѽ0H��C����
��:��2���/�п��hE��N s�WO7��-,6�P����<��l�����q���u��;�LuI��(��+�t�ECv;��a-F�̏���6Iԡ`D�[f�S�����sEr�D2�l�n$����Cd����47خ�[_a�r��O�=e�N���{��Y��བྷ��w֊��s�]�@�k3~ TNZ#���o��A�o���VS��(J{��V�m��ɨP�z�ѡK�^���1g&�ǜx����_�H�����{���wE_XV&K��.��Η���ʮʛ"�w��M�x,�xgy�����j�w�vm��`��{q6I 
cCO���/�W�u\J�'"n����Y	L������n�����QB��7cswc���ABH����ZTxǜ�f0�f��jF1ç��oS���$1�.��7'��'�Wڣ��U�n):gτ�QW��㊁ E��rT�"������]z�_���>�s틺7��u�A�t<�?R	�N�B1���Ũ���5B�{���r��M'vK�@��)��N7qfp͘�J~�,-啎�(X�FgH�������i�a%W��N���za}I����p�Ԉ`��M��1J	 uv�B\F��.�Y�(&�E���b��d�ɯp@�	���_d��.X�N7�niy��nV�ڋ�+3s5!KlA�!_��h����F�w�{x��Z``��U*Y�������r�!�;ɡ��"�4�1��Z�2��jͥ��Xx.c!G��r����<m�B'F0���氎�B��S�2���<����_��j��Ӹ��2��C�R���J۝-i�m��΋k�).�J�5Ś����'�6��T8�-��+�X�������@���I��mBMd���^(;-��r4'�x��ry����=�����L��g����̿C�k� �:��N�D.]�0��������V#��F��3ʿ,M	H^��D���x�����L���C�4����q������~��Y.�o,��o�P�v�N X-���8���`��<ưJ^h������+i_ �^�\�jnf|z�#���̼�'�������Zp�i��(���U�>"
Q�~`:������(��H��@���k8�����A5g�)Ycv>� ��SThj�gK}c��
��I:����2���\���RA˟�<A;�Co�-G��$����?�[��Sg���Wi>� u��DY$g�
k�!�����[q��i\�ϵ��h{��*�\�k�����6�HվC��'=��7��1`}[N9��h��'L��j�n���}) v����>��o}�gV���v7X�z��Cs)"!T�t*�C�x��(���u��ZY�o���\�Sz�G�Y�^�*>MW�,���@���c�+A��B[����Ԡ�𧉴�[
�}��3�&������yJ��"� l�Y;)%��������i^bI:�C�8t��/�.�|B}Yw+�'�y���s�S�M�ܫ^� ��R3@��-����`��|:�	\��83�A'�
�z�0��	GfJ'�4v\,�❔3��-ܜ�T�	�m�|rJ�<�T�cX�	��8��2���70GU�t����S�/��J�Ѧ�������ڕ�o���>jF�������o6��ѺPc�D�џ���sw�\�S�)���yTRU�E+���U�l�jk�TI�
'��Rv�H�~�Y*^�e�	&�A��G��K�2|�	�/�!�-�.�cX$��9�{�ao�dp�Ob!W�kا�{P�9���/�X����߸JQdƜ��P*6��CS+,� A.��w{*ȶ�梃��'�MC(��ȯ5��k� D�r�IK=�'��3���@��憻�y�).k��ɋEz���oN� = �����e��(��+ͷz�?���2� &Ϥ��u��V��$��'��+7�v�X��O(��v�e9a�x��Q-e��pB�Xdh��`n���%��:�2qc3/�J]�?��"���n���,m2w�(���z�5�>�i�AdK�sk���;��E^=Y��<~'�,�;�yő��[(j7�?�����V���OFm$J2z��>|�o���m{���0�[x+���@C�����ru_ej����E�:4�2e�w���3��k�z���e��>[�D��"�@AUN�v��7|��_�r�Mg2��3e����oi���؋kI�t�Kl��Q����H:��\�%�;��"�ٲ��t��N�.\q�Q�b���w��h�9K�|��H��7d�$xm���}�P~�Se�o���{��蓏�g�9���h2ǂ����}�;��Cv��^o����%Wmz�Y�c������S~������-s��Ӷ;���Ve�y�24.��ʯ�vʅ�/O(ʑҵU�}��@�7}R\����^7@��
?Smg.����{���o�dQ���,�v�>P�.��R�j�4�[��g�|� �D��H�az�����"�St�nQ팹�Y�(nH�����CR+�(�?�]�b�I��W�sa���������0ٿ��S�ʸ��Z�U���u�6�!0�n^9�c�W�U\6 }1ҡ���K��I��Lo.T��
�X�-%X�yc�@G�8�[T�&\�g��C,rY�6q��1y�n9a
<C_OMq.��WyK]�����\Џ�:���09��+���	��Q�-"w��Ͼ�G�*w�n�̮��i�T>��W�l5u!S�A�M���I�P��;Y�jd��|5�q��hT�J#�Pw:�g�~�{"]�Sdp�~�~$W�	��M1�N������VYf��ߩVj��`��$��N�{ۚ0����ö�9\ؘ��_[�8�Gpˮ�
��X�Y��$V>|��u�Yd�R�����5��2,W��!"X��_�
�*n�Q�!�.Ꙥ1t~����<V
�R@q����~�F��&�D�yL.S��-���*����G�I������gvBH!�1؋^�B8~_k�V&�6��wX�������Fp��[�#%\m��n�������`P}�wԡ�ө'(ى�*Ԑ9�.5�"��5�T�9��4	�o(a�N�Zp���<��" �a����W���ڽM��q��+�P*ՠ�wt����4p�'b�')E�u��-���^�33����+�ҝ�A	R����ES,��6c�\��0|Ȋ��,��M�b0.]޿B����'[E���9���j�R��BX�w!0�k)��7��u�z�]~�G���7ӭZ ��X��o�6;k�h�?U_O�Ë7���#,���D��p��%Ye�x("�C!�(cߑX�o����U�� ��u-���J3�	�3'R�x�FcU�@�H<J�E�M�b���&��*�;�o��\t����7�[��oq�ͳ����I4}Q�&����~��Oڲ46N|�r�ԉ�5+�Tw�4@R9l�O��E7O�Lo��3��k*�l��D�Ǚ�%O��@_�3��e�m�_�)]��$e>9jm�Zj9��c�����a̫k�a��ҫO��IZSL�jP��Ғ�ﮓ<k�(N���ev�`d���4��>��Iw~��ꌏ���w��8U�A����� �<�Ν�т��w&b�%讅�|�����L��� $;�PA�윢S��-�� ������td)E��}�$99�E8W�,��)Ԍ���;h�}��b�B����Y�k�sLhE��a!�%�ڏR�p�R��"$(W�z,u��|�^���&���B�X��0&X���[���v�^Q�0Wё�O�U[��v�>"�������.����A|o��閿��)��r9q�O���%I����I�O�N{��
�uz������yﷱo���x�\��D��	�\<�=�4��bc���5��Nw�'"+I����� q����M�93���I;��cﵠ����8��{՚٤U"Ӕ�ѝ��^/&�F,���/�� ����OP4I?8A��`v�^',~�5��^�}
���������2}��m��	��N��.�G��|X�4S;޲h���h�l� Z�n1>��Q��=�s�ϫ�˸��!����.6�	NgI�\̱�U�j��
��� �����!Du]�j[�L0l�!�O�X����������5$=!���):]����P�.'m�$���C�T~�N`k��e�D�PQ�7��o��0��~�����rD�1|�A�C�T��������h}v^��'m�
��8s5��3��n5�&�@ڙ<�>��j�{ԕ��m1<�qW��1<�],�����W��:��Ԝٖ���ũ�ZX�����hb
]�=�	%X	�]g�FA!��G�!���'w�r�O;��>N4M;����">�*nuX#X��둑�|�L�C���rٽ��D��:� �/K �����	�&�Dy�F�,j.��%w~[�g�2|v�4�J��pMn�
�+��o�!,�0���=�"B_b��=C��A��H��&����i�"���̦�G�0d3Ѻ��vi�����a�|8�)�#i'����S*��*�����{v�D�;C��n�rXA S7>p�1��*��F���dD���
�Y����S�v����s�9M�,Y�n��xpdx�L�)�������6#©�F�M�7��k�'��qj
Vd�FA�~c��r[sڠm�^;�C;�ȋ�=o�r)]��OP-�54 ���A�	 ����Y�jCH���Q�ߧ�����\rY��5����pW���Gp�#�iD��_<d�(ይ������M�Y��r�u�z;G\���?��8㵫�"�h��Z]�a�w���j6s�	���8a���J�=ޱ���G�+����aJ��*0<�ǯ'�A��-qy]H�� ��7j8Wq���$7�uB��RNn5�y=��T�����
p@��ۭFŊ����֪�*�x��
�������5�q<5�k���y��> z>ˢ�MG�X0��2+�[�[�^ѻ§9C��3�)S�f�>yP:꼠3�5��%o`�qG���!�ٛK:|	#E��ž}�7�`x7z@h�l����U�bI�l?ď�۪guiy�����K{��{�F��r�"�S��$ֽYH�k]rͳ��R ���f?��4b����U �^��=M��Nd�?E���|�O�!p (R����D,���S��Nx�A����+B��M������	����v��Ț3s��s�?�NQn�V~�0�������C���-/�-�FcщR�4j6/�/'��o�uI���$t�$���9>s���q?BP���dS�"Z�cm��J����,s��~R�-�0�և�풔6�ǁ��v���_�]+
�{����Jmf�
&P�_ bWL��Ȉ�����hD?�BJ��Aj���b�J0p"΁R�q���pp�x�;)o)�$��~]�0�h�iV�D�QCi3m�Ի������bZ+zy�vR.D��1��In��/��]h���o�̽hN.�{�9ɻ�-�x����k�W�ǳ*�?P�o�<������Nĉl`����N�8���f,��J�L���O\L�X��*�@̔�� ��Q�j�'�<��� *�̚ �\�%Z-�`Nr��[AĨ�eE����b�ڋKo�'��Fm�d����S�/(�`�)$U�g�cR<	��2f�/���]?����p�|�1fH5�A�<E@,�g&���g�����*�{�EO�-Ma�������j|	�9IXd)�umŶC��.��DN�_aq���)x��R�4\M�ţ�C7Ɗ�.��b���L�߰�ޏ�`��,4gf�����}��̮��~`�&c�u�p��<���0�����9��2���}u��)Ow��*�7 gͱ���S k���������w�����K��CMMt�.:�,@ҍ�gYv������w��]ꡖݸ�W~��mx�hO�eH���x�@���#������c� � ׂG�Vw%��>s���.u!:����m͂�W8������\3S�}R)�^��ɠHh�C��:�&��I�aR�-�k�XP����{���5�9	'���m�n�4�>�ڍq�;w��y�נ#������]p��^Z�딜L�X��� �.�7�8'�{�(a�Z(wg1�~$�1�D�	rRĝŒ��6�k��5��|���G��ü��+HO�~>%q-��応�U��	#�#&{�F����I�a�� � ڼ��Ψ�w �2���'���	m��D	`*�I�ƀ��Q)F� Dy�@��g�5�ZB�ôr�6�&�Pl \�Z�I��w���Y�������{�����Dmwwh�<{(^���������C�n��K�t?e����K(�R
3߁&7�̀q���:B��ت��)��X�o
��_~�@��'w0�F�%¤�k<�%z��s3��|W8��Vն�ް?�6!�p�w1�d��?8��=�_#F_��̚�Ŋ҄*��%��》E��S���+�'�b&�x�#��<=���%��I(�3�&�����F�	)�F��n!eSa�}�"2Gbm6����|g���9�Y��Z0�/�$ÿ�,�D�&�&�c�Bk�Z-#��d\�He��_�fB��*��(O�5* U	i#ܬ���ShQ>hŲ��H6�����;#@{�rΑ!H�[`4$M��Wx��i��ʉ�@�M�4Ҏ�LFcY��|:�c}'^��'vQjQ�o�����`Qzv�� 5�d<�[�?�\'�ѵ�Z��Rb�N�| U�t��i�p����z`���������u�9|'��`���x�v=w�@\(�i�ʯ2e��Ḥ ��y���O�d҃3nS���!���s8�ICpJ�cGș�=��)���kv�:$�{�\--9�c��M�(P�ų.m��)��W����nt�!@��T���#�bߒ��!C�A;�_M(���><�7�Z�<���.�8��Ӽ����+��v]���-�6��O:4W]���=��.<�~���2T{��G3h�'�A�5�C%�)�����И��x�� ����=X���r֮i�nz�_0�U�!Qus��R1.��J���w��һl�o��8�gY�[<]�d��� ����1К=�Ⱦ�BV��g$\Ȱ��R���H`�%����o#l�;�&4��݀�hi�����doG�n��*#�^��&'���D��_p����~0/�o�ə�Wn6S�N'	𑈸8��C$xp�5�D�Y���It;���I�1�]���!hN��xa��=^��_-N��g"���^|57"+��13_��y�R���ޗ�d���i�\�����C�.E�L�&��h8��3�A4�� �����I�K��6l@�p�`���J���@/�y|7/]4�-ť� �8�R?��X���J�6��pp
�f-w�C��88�j�,}��~׫x�6"�b��7�ʁoB ���]ޑ�`��rr�/Ic�	z�g�=���|E���c�mD�,/�<�<�Zj��͂__��_����e���˕M�[�b��z���Д�5�^x��`b�#��Ԧ�}�9C[�[2��.�abv��'�#�㦲;�`����Ogw[)�'���R�������R^<C�/�s���k�q��� �@�u�g�(��W�H����SPc�z�?�p����
�rL|n�&L����ґMhP�i*�{�����u	G�w�8*��utm@�t�:$���6�O �lh'!)n�\-�:���I���YB>�PB${�hxvT��O���5�<R�D�I��z��7>����J���$c��O���s`�v�؀r�L�ԣT]n⴪~��N�sS��`�~NxƖ�g$�A{Zh ��CO�mp�v9c�o��!�P��@���ּ��H!�(_GMW���˹R��iO����A����1G������P�6��Œ������]���È�؞�)b��#�,��I�e>�94cuO��m�yq�x��� -5�6�����Х�|F�������67�uD��߬���7NA��m6��FX-��ݨs��a��2��w�/���\V^9B���!N�Y<	�Tͼp���|��������s�z������.�/�8��h�/�'���j���3���5@j �# �@[W^���D��y�����@SB�Iw�^�
i���ܳ���y5�a�q�Y���x� � �r�c�����`u]�	�CY�J�y�8��K�u�	�0���sk����ĿT�Hܩ�{*b�O'غt=䍊fWqb�lY�PN;������2Sp�W"ɞ+��ـ���B*~����8hNo�H3�����K�/�p��j�~�.�V��O1� C�u(��Y�$���[����I��˱$�����$��1�z��9�%D�7�(�tbY�7���f�1`S�{*S|4�]�y�eE�;�(��Ϭ�}'o4U8�Z��q�@�}>�0!�E�(�f��s~���/�a�y��֨xA�����'�_L2������;�o����4j!5��'��Y�Y�K�DG��!q�g Q�jTHg'B>�	��C�^����m?��Q��fB+�D��8R{G荾"����dNހ�B7�?~�*�tMJLtN� dh�s������p���P��b�� W�ď��\Ĭ5�gaC`R{���X��<�b� Vj�k�VwKm�|�!6,4V�"�w��R]s��Gد0��zo��P�C'��1�h4ō4OA�P�~������aK�D��8�*-�<�i��U�N3�O@=�������8cEГ_�ɾ�]�;th�F�L�a�v>�v�FB���8��?Z������3c !�.�M8Z���o��J�
����yߙ�!�0��?#3��i��1�=��u���^E�mTgH�����C^�(7$�:܂:�����sv����PȔ�D����r�#��0�R���'R>�M��0���O;�E[��aG�u���]�����B�?��_�
�w|�����v���$�ю��3���f HܧF�h��yEʊY��_��*��\c+�H͖k9?~���y;���#y����Nz̵�| �;�ʴ*����p�b�ꩆ|5 ���l˻_�+��$��+6S�t��i�V�mN�׵ܖ����iӧ:�.�t�OW��Ŋ���R�m�9�2XB�,u����n��JE�[��B^�J�O�ͯ[ �}8'�I�`+{l�p��~� �p����&�4�����Um1~���ߊ���?��+h�G�� ����=;�1RP}h��[�{��b|�%��alVm�`�),ଉD=�����v��`�r�����X�h��!)_����z�����yI�b��#پ�~]�c�R���ؔ�}�a.�a���áĽ���*q�e�!q�+��q���SLc��FҜ�̸^��18���X]>bA�/�tB�;� ̍��U�DJ�/M�4 �e�A(	aj�v��̟��v�]X�]� ��ŕ�����.�+t��$u��Ǻ9�\oz��r��s� _���ѡ��@R��N���B���ӒFG�����z\�iBX�	lt������,�	q��S~����K�:���E���v���"���@?Ey�G�T���4��M�R����v��7y	��� kΙ�CLs�c)\��ρ��D;�r3������"�"�Ѹ�Z0=�jr㜎|��{�<�hbQO�y���´^�%�i4s���,H>��������o���'���u���{&Φ�p���B�B���U�#�3�d����n`q��{e �=��,��/�Y���.ɯj]5�:ZzbJ��4%�+��ƶ��R���lW~]� 4|�$�`�ŀ�,"�N�	v�3k	���cb�����a��n0���O|����G3��	��o�g�.��<H<[�B��y�P=%J�"n�	��2�[8[�^@&�;���}l+��D &J�ҝ�ڥeyfE
�^���-5ء��$�4F�Pf��l}O"!h��O���@���[�5��w7�������t�S)��jEQ	Aǽ���)X��_K��I����6�!9Ԧ��	�!�5��}��Z@#����F:��^���h���Ҧ����Q��1-ط�|���oP%���<�Jev�,�M�X��}��w�l%$�Q�Ŗ'��Qì�Y�w��W�y��@���}ݐ�;��̡��� ����$T�N)}l�⻍�P'��E�M�Mb7:�@m���2S(��<����`���f����(�
�2�,qІ�"������C�,7Q�ǎ�$��:#���jyK5�z���r��08k�({���#��ׄ[����tQba�-(�%d1�{ƚ-�bP�Vq B����TL�f�9��P풮�-/pO�.��rM����֥G���+N #��%�0�6��W/��eG7�=�ί,���i�y�_�{>��K��p��2wӻ�{1���}U����������v���(X�������{���S{*k(�k]V�	`g�K�W�}�E`��O�崎�c	Ȫ��lJJR�P��:^��U{=��ɾ��7���d�|��
�*�\�k�@�<C���ǥ�s߯��3����z-A>M�2P/h��QXB =��u3a|#��T#�c鵁YNT�W��t0����Q��jD���
[6����0	>m���9KOW#f�	$o��8��oG��c�S�fV��&Kޕ�����NU�����F�Uv+���)|sx�@L�
ppLYk�|xq �U3}MŌP�T"z��R�ֈEͳ��i�ȅ<�� ������R���.�!�s�����m�"�\���^{�[�S���w�W M}(7�;A���XSk����zz��.�uZ�홫�f��{���<T��*c섮ϽT�b�tZ��>u�h�&M��:ͯÐ���=gMN����ɠ^�P��c�=+�ll�x�=)�0�j��c|��E�� �g��� �_%H.�3���?�TR8(ŐS%���U�\y���R֣é����"��`Q��$�'�g�~�k�w�p����^$S1��nT,���������]��b�V�~?B�O���1/�}���y���G]�2ql��V	�˻�B*�c˪�U>.���-,��u���>I�m9��D/�?��y�,8��K���Zo�r�d���n����"�]��Y��]����zOF�|����KU@F��e�Q�c�9�`G�Rk�"s��(]��+j����;gƖ8�]�d�Ӌ�P8/�^�%_݊.�P��(��**�LQ���s�r��e~T�J���&�43�'�>UdY^�m̨��-d��=!����ظ��8�W��	�z�n����7M`�/��ˈ>����c2�@����H����}X��\ޟL0< �u��N���y�b�&bXfQ-�B�[0ތ�B�Xƞ����� xܸ$X 6Y��lD��Hr�I�c�8�ݴ��F{��bh}5�<`�4�0�F��a�`3g��'��ݓ��D�ภ|�1"�'�m��J-r��5>��$f!���}S����4o�Sш���D���l[זu��?�&�����,���.��f�0;�������`x��� ���|2P
��<5��7��=�%.�^�1(Y/˃���N�uT6ߑr	�x̥վ��w���t�-T(o�k/���2�t]�?�2��5r?IT̕?������N��4��B�T>)E�D3�4d���%��z���7��}�"�kZW^SǷ�����%��~��n ��r�8�T�?��8G�G��@�c4��Y���)����U�O='�h7��7!��˱K���;�p�/�Ab~zݿ��`r�jKN�y.�p5	���`����_�~����m�|�<"n�s1��Rx������#�U��A���l��Z�(����l�:��k_焥ϐJ�,�(s���Z��|��S1Q%Uz�3��Ԝ��c�W��ca(�5�Qt�_�Tx�>��o��$%�u�Y+�q�}��vw�U�_(�}d��1�����Q�s����7��u|�N1FS��=�9��A�r��2����W-������k�,�������qZ�A[�Nnҧ���z�V|�J8��+#�.z>�LZu �O�QA-���(iPt��@��ޗ)��S�z��.�J&7J3����0�i��b��XM��[X;P2��c��Io��[~�Mr�Lw��Q����q����S��"�Hl�:�/���{h��Bu �g��Ai�y���R�WB�f�G���(��Y�(Cq���	���3�~/��3�`��!4��D �ڗ�ڔ��}8�o	o6y����^�gL����Ad(ݹ�"9ǟO٢��_�����wd�);�n��)Gd}�]����M��7k�6�UԢ���P_�:@�����'����U�	��/Ղo�!��.�"��&��+i0қ��v7�Y�r2���]SV��n|R�ĝ>�h[�	�U(-��ԭ!-X�ŉ���il�����B�	B�Ӆ4k�y�����U��,�$dZ�7�)�[ �+�҈��$M�EP0�H��b����U?���`�!��Md��� �C/1ҋ���r��q?��0
�/����D�p�9�(53qX9F,��N��N�����f��o2^���p�
�/����Yy�6Ҵ����~Ttr����m_����3��h�5	,��)|M	m��'��L�z	m6�O�GT�C�Pc��\��.(y(�Z����A�D~ES��"�O�dd��ݍ�!�U�P�w�B�(�2��(�(-�:���_��aO`09Dق�7��?�Ŷ��[~�ٴ��IEj/�7�2M�̮1��6<��
��eK����=2�{U�)v��d
'i�tU�|�k�Ǐ��ſ�Y76�f���]�S�rʙ�t���k�q&[�D�� ��DT��@]���K4e�z�.:��9�cdfxĬ����+EB�f�����\Z��.�[2t�!���n���G?�f�*zx�ҘD=�u9�����٦�_aj�ȿ�L��^��kRy��&>�:��?Ǣ���W�D���y�pMg̥?Z���Z���<����$VS�e��"�Լ���0�����&�b�#�u/�ww}��CT��KrX	Ϻj�n�`�����YΏ�:zͣu�?JB��\��JS��<���ν����W�!�V����r_��Z
t}� ���Gl�9�R��T�����h{���0��r	�}�O�����2�i����c����`���v�\3Ue#r�������@�h�)cL��g��cim�0�^�u5�1���X(Z�c]��I�;�N6�W:��=��+���FH;�	XW1�=�K=�	�5 ��w���b{/ؠA�����4��՚�����[��a�����ܺ/��#%�. �dP�-Q|��e?ex��N,�H���f_��S�ĉ���^����+kj�E�r�EbND�������ɍ��l=u$�,a{�����dl���u��5M�\���;zQ�5U�"�x����<���n���]��:�� (�.=�f17)4h2��:��AFL�RkA���q�$�ګT����2�6lu��B_��҂���ruh�Ȳ�.�m1�1f����[u����y��\�ѼVʯ9�Z��	���E��vVWpܬd���I<�ne����~3L���֦a��^m�/��ܦ��<dV]z 7���#e�7�=	�\��	�8�d!�=6<��x�WQM͍:2�jy���k��Lq���B)F@��%6���.��V��-�g�^apJ3�P���}�u��� �L���u��� ��n�d^Ad�����B/�u+�����otQ@`?�vt:,� �D��tD�������Q�$�4?�4̥��n%��B��x�9�rj?�G�.�O.H�^i��1(�x�؛8$|˘bW�q@�1���]�ո�cu��1ʥͤ�S���8U��ڙ{W>�怠l�/��/�bsf�ZG?6��C��T��UW�+H!B�Y�U��&��ea?�zq�k�*_��S��D& �bsV�.�%����fD��\�}0��1CA�8k9�~c(s���e@��a���!;H} ���ƢER��D}6"§�}���
K��@�/���"���CrTݫ	�	�)�3.*���F�Y�X�5B��--��+��o�GS�E���+�)&�l��~�-�W��(�2��檭iGz��0,ω�Y���3Vm�]C�S�F���%�u��3Nf ��4xj�$��Л~OB2�[�ب�9�޴8^�߮3��'T�] /Z�Q�b�W���ݯ9X�A����������51Б{���=���׫����}�W�|\�IM��9���b/��B,��5������Kpv��q�<(�ɳ�3��Ջ(��O��'@Av�O��k�q�o(�����ԡw˓���Dn�^�/"����6��MU�'b|�3��6�����F.0��g���d�8:���+�y��]��uzrN��CA1!�d1��Q5h O��f&��$x��W��r.Ҧ�,`�K�����6�	���OWjS�b�7œ������.�m���������S�S�t/��� ��ؔ����nMgw�5�Ҷ	�9�>��9ݴ6%�,��-u�F�$�Ac�7������C	�5fض�<�j(�y �~u��͌�#�(Mu��c�~����"d��'�Qu*������5�����sxW�t�@��� ��#M9��B�wEn���Xk��d�������z/�^p�"x��3��D"ui��Yz� ���.�s)`.tAcm��k�5O�Q��*�	�����k�蝽�����Դ��H�t�����:�	�P}6z�Z�N��z�K�:IW�s�1���Eu۾!w�a�g�rM9(?}���4�Q�g}��� ��!��`*+���YYj�^�B���N�o3kl"Ԭr�O*w:��⥜yQ�G�X�ֹ���c�xYfs�-źs�s��g�9�q���Г]o��}�t��I+f����qx�]�G�� ~xՃ��\��G�h�*�"5�����:���6�w�*��_��7� �}3B���P7{W8]��xqcq3?	׀��2�Ӆ��6SRj�0���9OH�!��H�m�L�L�w�n���
�'�3��z[.�O�Þ����ŗ�T�$�z-��n�`�fנzݹ/�{6���:t��b���z��0���jgx��˫���Ʃ���՛
M��;�����J{0��\�Nn�)w��!�i>#0��h��(a$ӏ}s�ڱ��_�.o6��xUu�f)�\��o�չ��fW$d	�������&K��ԩ4�1���Yt��f�G�_���i������y-o�Q�3K��lqRFLg����=���G鏩��bת�R6`�:H��Nox�Y@�p�����̳ [��Փ��d](�m�ς�I�Bn���i:�cjRl�Y-N�I[R�Q�';Ժ��e'û���#��6���\��O�p�g{X1��ι�����m6���r����^d�"Aw�v�g_��6'�����q����R��'y�Td[`�{b�`�ՠ֫0��a�?�ׁ&�-��A��H�Eè��=g���Z�|v��W��CT◤������%��#n�(�ƝQ�>N�ɕ�,_��!�1^�/� +�	%�T2@�L���/��Bk����kj��CQ0��g��_
/��W�>d�2I,��z�9����V8�����W�b�$֑U5���@��R&�'����18"�vtH���k�~�[V�������$v�U��X"K�&�]0��W&�dj�o�Ll�À��/����4iﰑ������@2�<�&v�?�l��	,��Z� ��6~��R�ojY\��'�$͡��Ii�*�)_���t�&*g59P�H t��%��1���&=�T������k��Y̱�1RB�����n<��w��|�F�֎������hs�
C���`���K�(�]�"I�%k���г�\/A'��D���3���q2d�b`�ߴN�Й�D���9�i/�E�7D�+� (>?�,���r to��ɞA�F!{*��
S��˗�ō3����Q�5�gk[��������pj��B��JUC�j�ܩ�YsH�^)uv���	�s7&�	�qZ��t�<&g�!��|]nl�u�}�K�kz�1t���<ϓ���P\]�Y;1��o.1{(��6cA�|�8FL��h����1�qD^[(1��ʉ%A����9 ��'�8�{����$�V������E��m��֚G&`A�e�s�Z>�CG>��ӻ�]SW�j�t� ����
X��'/�b�>w��l�ڴ�_�e��ӄ�O1S�c<[S�(eG�Z�"�s¡a�
:j0�O�ӋS/%����(�)]\��kfX~�m�z+�t��odTJK��xR�ǻM��b9A0{a��A�N�B8�Ʈ�.kg��)�Τ>Hu����"���Ia5$�rԀL����i���]e�Xo��*�9�|��2ے��4��ZE�q+�*!|�cC�d�S�u9�4�mv�;��tDi��ߒO$N�)_�������b�i�F�W!��A� D\���g��+�[��&G:�c������e�+0�k\b7�3��a)��VP=8�n���Eܡ��L$�s9huP*��)�&�c�h>��>�c�����8[|�$�OA�Zw��X|�B��I�x#����4/�,�ā��c�T��y�l@Z%��k�ɱ����0If�t��%��MjY=���`���6���"�8Ёu�oc�#�O* r<�������>ws:X	��+H�Wm�� gx:zrK`k�h�E�׽�BZc�����+�On1�"|�btvó�{���.)�ǂ�"����3��0~���c����wd�(�6������b�&���/��L<@����BJ�^2�V5Yi`~�8��p���2��Fj���]�����`RA�*"�Ѽ�ӷѫ������zj�z�n�29�*���υ��W�g}`i\��!$j�$i!���`�2-�h����$�G� @���L��	�L#{!}/��lT�)�$��k}���7����R�V`�r��x=Ql�*���z�ރY`�YЬ��%`(�	�Ԛ��n�s��F��Փw�攪��'�BanH��#Ԝ��,"w���_�,��- l@�cW:��Wĩt�߀A�c7.����{n�%���QB[�Tv�Ƅ4��y��r�	��O���k(6���0�s��*MI���C7n�=z��|�C1���2���]����tmj��F�H�XQ`�b\��̞lz���?���ҵX����Uޚ�9��W`t}��9��_
m�-�]5��=!e�a`'�R�B�5�&z��֗�=i_��b)}Ĩ��8����� ��q�����\����D��U
�$�?�~�ʶ�Pc/6��� �A_�d^��c��ʉ�=���u]%U}Ӡ�=sl����r�B�b��S˵~j9� �M��q�@x�X�I�4��\��b�u�s&T�k�H�4����b�h4��;�Q.��9f�@<%�M7��S!�O�,����/;i��uhVv�Qi��k�J�	)������@>^,'U��{d���%?�%�M/��Y}4�)��ࣩΤ�;-��v��n"�������^W~\��ɪ]��k�Hܶzn��53�!v����X7,ė; FC�+����!񫩦� ��N��6��ȯ�p��!ׁg�~Ҟ�wT��O�Hk�X��^^<.
i�$<�l ��p���h.7`�U������T"%14'4O��\D?&#}m|�ldʃ�gr)�,`	��0��]�����d'��,�kR� �a9�,�z��WY2�mZ�A'�dhL�0l����f�sù�8�����NƟ )�~���Ј6��ʬ8=�]9Z�����}=S�, ��*�_�h��2]�]�����)-X��W��ҁ������Ճ��BN���r|]�W<�4D���9�2-G���Y� kY�~�^`�8i�G]K��TЃ�D���N����Ɗf�4)�z�`���B�k�eO@!+M��Q�R��+(���M��a�XJi�Ԧa�SmI�	.@?��	��%��n8��_�'��O��j���&�j����%u��S+�^�닜Gz��c,���@�	�vL	��5�'9@�;h�*��h�#��`��
���t/B�k���WИ+��� Ա2h[a �[G�仰���:�����RKa�+��ГH��XkȾM�Q`��v��<�{��!|�@;	`�va�C2�.�k���;~��ڢ�h���~˿�Ю�F.B�3W�B��5!^a#O��MS�6�8��@�9�}���#;A��Ж�a	A��90
��7O�(0b�T����'/K3o���bï[hAm�a�B���Qk6;�%�����1�fJ/���"����9%��)m��
���j�~ƴ��*�}�flc�V�J�)�e�+�݉�u�mF~ʣhp�~�*)�sT 6r���!:g,�YڕEF�[����r)f�[yk����[�}A��Vt��l.H\�*Q���c^�𐝁ld��|�@�pOB�LBB'�>
��Q�D�Еpp#��
�hz(�������y_����ew�;?j �����)«&:v�ih���ql��s7�-�@�+Fdca	�0��d�-�p�F5�}��l�}�F���x��%����3��Nm��Mn��C��%|�����ZǪpm���Y��M���Ϲ�{<x���:f�R�n?�,jXٞ�l�")�g�U�Z�љ��7l�@D�{=5�])�`�&��ǭ�w�#�K5�	:\��S�ۚ(X�M�,���8�[k��ֈ�ڡ��_~�u:����P�)55d��+��w��#�������H~��ey��쮌37�]>��+)<R�W�'�STAVf�kcM?������`[!	۴�e�!� Mb��5R3���~�(��ᬞP�߱Y4�"Û(����5o{�L|��t�a���b�D�X�׫�20����m@�GD6}��d�Is$�4���f�X�6��z>��תּ��x�W� �q�T����i���:̨ɩ�x�#l�Jtz��+:AD.�i�`� �²~�p�]5/��(@3J)��==\B����>�}{�A����,r��N���8Q���@?3��1&.�����V�p0.4�o�󗪸��z�T�����fD�������T!���xRußOK�w�N�!2�[�@Ӥ�M������S�)2�R_!�/��U03�N����R|��o�P*N��	=<�e�A��0�5B58�����/���m�h�OH��3��8���_���N^�c]�縶�R "I��j|"r=F�=.'kY�*��0���~�7�`�oaˉ�3�R�<�`X$һmG�С��U٩5��-3����C������T9�k{ĭ��ͬ2��=��1Xa*�� �Vʜ�#B�� GJUX~�p�%V*BF���2X0<A�Z�L��X\q[���fϭt$����BdrX��K�������C�8����X*�d*s��t�>SR�˦�9�g�F~�2�%i�9������i�	vT
��XI�EP���Nc/7�|�te��+n$�nu�Z�/�Gl���ҕr14� �T=�gs�h#h�I�A
rw2g�&����_<84���+/��)���A��H|s���*͓Y�'�a&ܘ��f�m��ʵM�[�?�n����|�D-���?��22*gNg�5��i��@#p&e�*E�r�3CW��q�?L�O�Ⱥ��h��^�5�lu�u�΋g0��3Q���.0v��@�&n/�*��~�-����s�`Y���?�Xyb�"�3�]���A5���Vi��#�Q�l�8�)�`G<d���K�F��4P��,�z߬[hf�¶C�-��ծq^�.e����������j���$D�f���87�b���)��0�>8����O"?���L
�Ў4ߙؘ���OUq�~��g���jg0�
�@̹��m߷Y�L- �{��y��W"k=�8=,�{�Sn�7_���:�	��zM �.��V�} �%��B�
!^�~�*���m,�SJ�/#��d;3������}l��}UR:����ҥm㶼�V펿̇��7����)�Ec�D>�M߂f�@��*�e�ݐ�ԅ0�s��vRck���r�wp�����4��B ���^�D{��h���t���3A�V�Ԃ�K�¹	Juf�J�D�0���#����9��B�b�!�8A�(2�D�����-	;W+����/H�-s����l���q���\ܛ��C�&GN!���h*`�9�ΞG-�׸��gb�ȹ
�s)7K����hS���RЦ�]�I��0gs掼Q��+�+#�6M_$4��]r�/�#� ���gl�����7)�߽/�P.�}V��|���&GXP��<�*w�4���'.��4�$� �0f��k�FY��+���Rva��Ǭ|�e>t�sU��AV�^-k��J���N�H�S�J�tR��!�	����C���;%c��|Uώ�m��c�bǑ���:|+���EM0��p*�:�G��:���H~�D��<`1IH�߆�wuM���6��PO<����3�����?OF%������?�=�V�+�Fd�ũ�ID]��/iʬ��vN �J��%<�bK �ަ����$���L(�M����;���˳�+J��p�jT��z�tr��l5�)@�� m�$?�,���R�:��P��+V˸�̛���/�T���$KpVT� 6XxF�[�����~L����;�Ju�aMEi�x�;(�-[:4��L�Dr ��#Z����D��"mھ�%����,�d��v�/r�b�V��v;r,k��cw��j� �_���������l��T��͖�q���x�#mfSLӹ�<
'r\��&���0��)�!�Ͼ#,jR�B�rđ�$~�҅J+�^og�r -��a��$vJp*c
xoa/���#��1�yI�7��(I��"ׅ�(j��WZw�v�M�hI�L�e��UN����}�٤��M���dj�v���>v��>])}��Z����9w�Y�.��-����p����y1˶�J�v�U4��iM�;՘AX�t`α�����i�ٙ1k&
��U�N0Sta��=�,z����c����]��a�����L���q%qt�iP쨈!j�f`�e�22�
Ho�@�^O�4V�3�Vy�rΰ�}��U�\�ͬ�FhVdD���s�2��l1�=z�r�p�jd�Gu�Y�u�y��z���Y� �d�s|�P��E��^�!$e�®?�{x,R�t���_��N��Cw�"�x4�
������ׂ`I���?+(���2���ۢi�ػ\�\b����U��N,�O�s�vXl��v�5�]7�Lq��i�3��|�#9Um��PnOH�*z�>+�>� �9X�j�ō�-u�O~nIՃ��uM����$im��婍7��R�S����p�D������&\Ϋ)��)m<��:1�4b�L��`�gʝaF��ǊQ�|3d�98=����H}����˛@��qw��.�v/V�S8s�лd�M��;�
h�d-E�]�.a܆P�G�zO����`4���zbI���|�`
@�,MvƧ�`�"a�VizX~��
h�$�0]t�YD��uuJ.8�&(E�d8~
�!/8�2r�ax�76�2��Z��nI��fY�p�����sl}��<n9�(�Ja�����^��,s��o�2����]�	В4jW'��1��ɚ�	�M�7u���p�'y�Oq�]�-��)�5��9�BZ���W��3��S�7�����V���?�\��p��oJ"0}��))��p+H���9�q�_i;$z.�dk�i dأ��
�Fw�lp�A�I��wz3) 	,m.e��K{pl �� �k��$��h�P�S˰^e�"��Ǎ��J���/���I櫑*����p�i�<vy��-n��KyY�p�k��_1����u��!j�<��,}�y1�a�>�I:�8��a�ɶ�̆�xk�?�WB������I��q`~:q��e^����ȥr��f�b�	\��W��<.�_���X
��!m�"�BQݾ���R�OUH�/����,���~�r���~����;��7ˠ�	52kK�#!�Ai�k|�;�����ځ�j��&�{����T���
�,��BA�X{����*�)��,U��Z�~���f�I`fHl�7u��sV8��EQ�G4Ɉ|F�|�/��/V���y�"IBF���Յ���8��WB5`e^�}�~��h�NDN���tT���H�үv�P��_�!L�6C���Ǆ���.�t �����_پ@�:u ��RR�r���Q;`��pN8㌼�����Q)��jYҙ�weIxB�� y����Fq&ph}0KQ9�G|P����:�st���?.�5���}��Ȼ�:�2�n�u���o��l�)��tPho�@�5����'�Ȑ}�L��*i/���*E�����d�G�%�/Īy��ō��$.t4��ļ�h���if�*�1��+NlasGu�e4���0�H��b��p~aj�?���н��\Yc��j�l+������BG�-W�7K�g^.��������I[S��'�%x�~��nk�8�{���;���fi�cc��w�vŶ�r�	ƈ:(��%Q���=Zڰ^?�\��J�����,�⏊ ,�@V&�5Q/�vBu�4���������q��+����d�XQ�-{6T�S�]�w2������IbϣZ�P*�ToG}߹���+���/�F�˝��m%Ѣx5�����Y���HA��-sd�� أM�}]#W�Hd��VZ�����,f<f���xe�σ9��3X��+�@��zW�](ٙܛ�K_Y*��o�R��eD�/!ֿ��W��vS�D9�%,-�0��%���L��]��A�H�Q���Ұ6@���'qT�ǫ4S�h�k��a;mg㎗�׭@v�W�85���`a/��B��
]M����c(�����^�x9�Y�4��=�9�CӛÙXIe΀ȉ�C��+�0U���m����i8z,�V��Y�@1$s�z�!D`�M�� ���_��e���@;���]�����fE��Y`���9��.��������[DOڰ��9�5q�o���]Q%�T�ggS�	�t�b�Z�9�_��Y%fʊe����@�*7�^�Ӆ��d���dN"e�ˬ�ND���11Z�}
'Zu��ܛׇj�P��wC��꺈ظ� ���!�K�[�;3�S(`���j��i��q�dg�t��ϸEB!�O�#\��8>�[�1�֚_e��Q{��ߢ$%�"R4V4 ��š��h�t8i�%O�'-��EXI{�'	&��n}�v�C/h��'�,� �X���{n�:��b��y���-���X>%*�Ѱ*v��Q�.6Mͣk�]D
�)���D�/'��L�"�0W�=}E�P���/bd��/b�m�� �s�-_�d䖄/��Ǫ��O3���o��Ղ1�^�Ĥ="ls�������κ;䍕���@�}��q[�1z�`'��Ko�h
��8쿾�����k�ٛC�a�.�
 ���Y��`l�#�'�C����~i������ PG@�P���H�6$1Q�̍0e㿬�!�EOp�,�f��CE6��{�M��z�ugۃ4�En+y����P�}Hm�Ž.W
�m��oDxC����	�����5�*?�+׊p|�:�)�Z��ϴ	r�ڛL�^9zU�;[+�aٻ1H(�|�	��X�my��0�0��z��X�@�|Ͼ�Xy��$�,��ǎ�{��X���W�)����4#G1��i?VT�p�Vo����Yy��n���=����y�}�{�>4��¥"����$Ox�а� �ޱV}W$ځVRB%C.Z��NG'o'�/]T`T�곒��jXa���kPΪ�X��q:�T󳦾���
D���A����};}��g��~��e)��zyg`Re����(F�s7i�䢊�TX�'-���S�f��2�H�[7�|D�j1P�quY��G�焌�4O�G��TD����w�T	_���LN�5M�yZ=��(�
G��݀DX�j�+4�(3;Q�t;���놖tng��Q�~�_�W������K�v��	�(h��Ԡ���]�h[��R& WY�u}�S�$$��@�}?V=q�^�����O�k:�Aia��Ge� �7�Q���><,u�Z�����y����7���K߮\��殠,���'��&�6�!��L%���P����$<�=�95"*B���N��4Y4m8�N�0^u���͢U����זLX���������Q�O66��׃��������X��y:����$��15�O"�@x�|E"����`���;�A)=�8��M�����*���F�Y.��=Z�[nv�4���Z�M�U:���ư�C��Y��s�]d�WIovy�4�i�͎~�AuNˣ�Gh�[��V��X�ɒw:X�� j���w/рR�ˀ����v.qV�G��p��ԩ��'Fc\��
/�ާ�Z���4��cwbP5�y��\�)KB	�ъ6��, �����~n����	!����+-���nJ�S>8�m�YwЄ��``�>���q�(���`�.�uLfRs@gS	��� n�Hu4I���:YEρ"ײ�k�8�)����R�2����=Ȳ�+�B�6C<���	G��'��&�L���K.��R"��la�y�7���m�y�-�]l�K���)fҸw^i]�[����^r%I=� �^쪲���^�@*�Y���-ߝ4g�
⋽���	0\��ia��q�W-�4��� U@>��34�紐���	����<ҁ�i�<h6|:d�	#?(�!����Ir#�\�nx�M�i�D=R+��9��L6�/�$=��;���Bz���g�0�^��x�%6��-X�h��ҡ�¥���GF�U1��:=읽��.��W��w��9�AR���XŅkj�_��^�ԧ-ۤ��B�c�p���[�Q��=w���e_ivz �U�����Y�AN��Z�C���1�^�0�Z�Hc��DS$���	5��o@�#z7R�
̖QUh�afD��4jMig��_C<2ibwb��U�ȏ�:F��ʪ9Z2Cȓ�z6�{��+�ݝ� C�����Ox#X����<'
��j��qtt�	�t�o����`/�w���DJ��
���b�Tǟ	��fS�v��L)�Ņǫ��lFY�>�{%·�#�69b�L���}��Ճ$���'n��Fwʷ)nW��k��
�>�C$�j�V�X:{�s�c[���NN"�U��̖�:��3���v�6��L�"��h-���a��2�Ȫ@V����l���gV>{K#D\�5+�����47�)�»�=�8j��;�\Ϙ~4ec���=�f��h�q�ȡ�ǯw��@)9���_�c���[��lqE��J�	:!=Ѹ����H9¼˶O[�_>MC	E��M�,]I�LS�W��yA*���uR7��.�y��+�q��{}�_H�^�¨��!��v՘\'���N�*��ҮAa�e#7[��pT)�_���s�º��f���"�c?>!h�W�se���|��4�xd�k�<�!Gx6i���G,n)6}u�W8�����C�8�*�(��H����i\�q��/ie�b�)�j�r1&MHd�b\���ڛE�exW?��D�F�l?��͖}Mmp�)nE4��$�$}�cf��'�K�,���ρ\�����+�!"N����v��u������&��j8\�kc��Y�a�Y�'���_�8tD��:
��e���m���	��R�uMS᪒A�ݪ��s��pV=���"�J$�M�毸Rb���b�&��cc2�����0C��%w����4�wI�cb3H�m�X�KTݺ����jO���3�#�,���a�b4:�a
��S����e��@�􀶴�"���"�W{�0P+e�X���힯�H{�
?E,EOڱ| �-l�'��$�H��i�� �?�$�р��"wz�'ڣ��J����%�.G�	����d��cD�f�Y���րw{{���MW���*����Pt��*���Y��ՎH/���Kx85�Q��?3�RT��R�{��Ga�|2b��^%�,�(Ha����DYwhS"���)�b��7��r�hh������oQ���{�tW0�I�Y�;��,�r	 U=���@��ߏ��e��Qu`�9�7 .�Z��޻�w|hI�q��@�qM�W)�����Tar����]-W�����	����L��W߮؜[�*������D��N���R�%h�b� �PP1�φ�g �H�^`?sAR:�:��ř5!{-X����;@X�g�N,:5!|���>��4��&�Q�n$�7���� �۸�2�(BF��<g��K7��wĺ�,
j�>E���R��CS�N^�W(y�,F�pw���eLkGC>�fl��]�E�m�J�;Cke���n�Eg�g]T�!�И�G��ʵ�`V���ε.����c���c�͓Γ���J*|_�K�p̓���_�����8]2h4�k��uH(NF�uJ��-1��	7�O<SY��G^���45�)��l�F� T���K�K�Z��!Z@H��@;5)k��-s�@a���`���!�1��o�v�;�`��q���OHO�dQޔ6d)�EO�B�aݐ���-��]�,�E�T���<��!�0cQs>Ӥ䖝���+�bҲ�F�w+���>Da��
���q>eM=���*F�yn�����Gbx�Յt���Z
��[h=-+��~��7�ͷ�s?����kSB�O0nв'��C����g�w'�"��."�Ü�y �bx��
�`��%��$U�rh ��{%/2�M#�°�F��H��3�oB�\
,���t|9l~�.�f��fAVb��]f5�`�@���'�~��O�ZV�б��,eD��$�ʦ������E�R&��bŰ������9Đ�ܙƥ���|B�C���&�lM��E6A|r�s|H%7?Ӓc�?��2�zW�J��,='6��Y�$���b�]�L����P��P��c���4;�Ue;��e��%b)K�L��|%S��e.��pPq����,���b=f?��#+τݙS�W�4����A���/Ԥ��4r e~�t}yɬ��"���Yc�2H%i�_vm�����aj��yG��Ύ^�t�n��V��U��]��]�kS�<]D�6�w�r �5�T~I#�VӦ4h�N����inŶ}/���ׅ0@=��F�ʚ��D�H0��ODì�H�=yh��ώ�H�kIck�����M�+�3�v��סP*�m�k���!��n|��*+��D�1O�!�"BGf]O�F��V��?"mZk�����V�+٠tR������v���@���F�FA����2=V���j���ӓ^4!�X�e8�q� �8atp�	F[A��JX�7M�Gj�r���t��&�%�105��~��&J7G��2���u}Ñm'��e��9��c��Ů�[*?B��K�?=�B���8
n)6P�0B�1���F6>Ѩ���U./��3��6+̷n^:��r�ȳ����R�-�]8�e`��r�s-.�