��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��Nڭ�	�����B�#Z���?�4�j��0�ΐz�A�y�[��I4�fB���_Ɛ���-����B���M'~��k,���'zf���]A�� -̭���ҧ���D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T��P�]��h�� �x��ɻ/�akB�����L%��s�A�ۆ�)�a7�$�HID	���� �ձll�ɱ/�hsp2�|�U��%ʹ�	�݌�Ц�MCC��C����I��1Pf�A$����7�4���)�"�`C6\5�'Y���=��hJ�g�łIK0�.���;N�T��ǟ5��6{3Y��9c9jB�m����m�c��QT2�TU�o��&���i�K�1��d:�%���ܠ�U�춣��q�$�ҏ�l1�ɩ��o{��cv}�Y�d=�j�2��Й��6��v��7�SΌ| ;���7Sf"�v}
|+L��ܣ�;vǏB{��L"Rz��N�G=z���C�ΐ�[��)�#�����$�j��"5�"�K�/J) �1���p��(�Sr\��(	0�|��(u�Z�(�ӳVKW����k�[6`~r��DS�S��4g�S��@*���M	;�&�$_GJ!@���~rb��#�-�-�Q���N}�B��S�x�Z�Ӈ*���������dzs~5��z��(�X�@g�Wxv�l��y-�-���:������ʴ)80Q�T-�3�7����v���M+��Ht��$��i�;��f�?%�����;�O�J��Mb4��U����q�j��i���8".)\��1Q[Z�aҢH� e��e�OM}g#X�dp�n��~4�H��G���^�� W��͗�<kcO��v��j��/��	UK�� ΋����T���P�v���+��]D=�X�'��͍T
�n�P1o]�6�H��������YfӠ�}�%��	�����<O/�uY!���5��F�����+R����;m�o�� ��\���]��/y�S���%��"6�F���>��UΡ>�t���8�;1]b}Q=�5��?�1��>l�����Z�8����_�a+ʹ���^�6G�a�{gR�@���I røp�"m��N ��΍��)�m �W>���T��n. �����n��&^�iQxD�s$~"r�À�8+�.�e���6
F5$2ۯ��H;\}���O����Z<�(/��%�k�����@B��k"�b�{G��$�d�Q�f���1���kq�.쟐'�!O�9��ѓDWD`M�����6�M�9�t��g�~�&~~��p�����]�K�v�N���!ȏ���o�`�a��O�!y�f0���Y� @�4�L�U~s��w�>��}V�������<�T*d3�f�aJ9�O�=?���|�߆Ŗ���)�K&k�S�v;�£;���D���:���`"[��Ǆ���M�|�i()7��tk��і��W.m�%E:/�5�J�5���hw�sS��ۚ�5!���^D�jW0R���TQ�5"3n	>y��MΥT
id�P��4��#&��ѿ�+?\ )W��hg�E(�m���4�Pv�����il'+M�P 6�e,#�}�%��!���B���9�3�D<��ŨƧ�~��F�I��`ub��'��m!P�I���������-���XB6�.'�=���8)����s3���>5=f�m�
����v���J����R@�^��8�z�X����I���V4���؜�H��Oal�+7����cl�0�l�,�&�)d���l �U�ɱ�9܍��FOP���f�|��y^���Pp���C�E��z�}GA^�0��Oi�N���%�+��|����H�j-�v��v�݉�S$�Joꪳ��["l����b&O5S�J��l&�Fg����g6���C �n�z������#p���Xر=�2�V��l�wΉ�J�]�������ؾz�u7��ф3��}.]Y6U��Fz���k��2�;`۫�� �Gǫ��6� cv3Iˆ�\8�+�Px����?�^6iF�1k3%@�@��_��h&š<	����|V_��]�-��Rp�4p�w�0ҕ�(��hY�>h�~M�Y��F*�
Čy�[��:�3�W�.Y�3�.RCl_��!�zs�Au������9�����ܟ����� �eJ��x��������� ����%�GM}�1x�s�B�@�M�I}��>7m�t���s+����sc3�������5\�ĨM׍ݽ��D<C�ھ�>p�<�$ �F(2���<�~Ɂ_L�S��{1��:��Nj��Q�3%PLQ�{�<L�Ah�M��> ��͑��S�յ����G$c���_݁_k
��Z��(9]�N�M�;���y�\6?��?�U�r	Ñ�M����e�%T�D1��������M�d%����L��ⲿ��ڗ�![��P�������+`Lyj���,+6���H�v+h<t�zu���#,8k�����՞˚�\�
}-ll�>Q�m�q�)y�Ct!��h�^�S���ʜ�"����D\w���&ϥ�z�K�w~�6���W����R>�rY�A����[o%*��<{����l�I��8�Wc]�AL'*�tE=K&�m�
�Ն��e&[�G��z�} ��Z��I �	��F��������%��ڧ>�MIa?4�LK#����Q�Y��[�������cF_s��v�������.@�t���"�œI�~�9����7aqK�-;æ[��Y���Ѷ���W�D4 ��6�p�h6h'��[c�30���j����_���9���|��n7k��*eIQ j�Y]�e��w��� ���8:ZFe].��z��Շ�� T���m��9S.a|2��(#��T�� ��x1��2H��	4��G���͘��|�����{bb��a�lxF�OVnrU��>��%!��Y�vM�n=s��&"j�z�!�®�3 Y��%nϨdg`�F�x�=%�����8�X��0��K+]B��H(��\o��nv�y�0��Ź���u�r�:����8u\5���}��P����}�B��T�Zi�!�\LBr[pTY�֗t�tV�6���Q�Z�����}���Az`�AJQүC�vEc��� �d!]�b��sC��ce4Uc�?@�&�Ȏ��&� E[�~��Ů-� �s���MF`,���,�r��H��g� �Ť�)/.�U|#x�Ȼ�]N�BF�.'��L��;�s��D�HBz��8A*سh�l�l�����g��F� ��Z�[�H5tx�T$��@u�Ld�h�a��^�U����;|����) r��q��'������2�+����-���rz\&� ���Sf�d�+��Q��б��+��i�	C.�|U�Ὧf.Xn�B%�jS�W#��s�S��~��]8F�H���Ƹ���z��,�ma��l�Db@��0s/����&}����hĭV�-��_Yt ���nL���x�S~�y�(ِ�;,[x�UY�Y���AV����#\�^^�������I��c�i��2�<E��nb#�V&�%�MM�6�c���9�RR�+���F�Kc�m���Z���d�E-������5��KN+���5�ՋS��7��\���c��\D)�9�z�G���pQm�/a��'GK�ˈ���ڬp��tn(�
�8��rԀRH�F5�'3���Q�uԣ|����Ƀ���h�ޘ}���<�H�Ca�6�F��8S?�^�%"�j\9}���eg%�2���� �E)�vYt�qmN�(T�$�U���� ���|��b���C���	A���5C�,)E�$��G��g!����8B��v���(}��Bvf���M���R^� ��E�ᴮ���M�o,*v��B_'�|��i�e�4�p%�#ޔ�,�Vur���k��E
��J�,SA�=�d�ͮ� }��1�TK�n�U�+�?�/ٖ�r�#��$��c�]7�3> އ�NR�J��T��e UW\�4������T��`��rY�߸O�m��W}�O>p޿����J�{�)~�ǅG��4�*�����{A2#��!O� 58���I4k���G�Նf����03�mD����$$"k�!��@HK����Gw��7BZ���c����$�@��4kˊ�L��ʈ�hE)y����Y���)GV���f���
?8z-ֲ�I}��`�Z��몽BR��U�K���^�!�0 �����\�ՄH�\2�����U����gu"U��=^���y�ܫ(�Q�{/�G�Xn��7;��780c��ݷ7�mc���IV�i�K�Qc��SϷ+�o+��")k�s��j�xl~/�M�e*$�7 �|�|T����M�y�FP�l$5A7�˝;�}Q.'
�Ĝʝ?F�8.e�
률�A��mx΅V�Ι��4�#��+B2rP��e�(�����G����������H�v��A�oW��b�#Ck�ǇL����.�o�܉[���`l'�eh;��6',JbgG�ė��6?��7�]����l���۬�7��{�> {����1�\` ,��k��N�)�2��$�mw&}
lI�1w�/�U���G�J�s�|`t���Jȸ��A�v|�7	�}*�\t�˵S�Ê㨞ٵ���D?_Q�Ar�&�&}9���*�(�T�����K�ƞ=��z<�`rٴC�����H�i�0�Ԙ$�J m]*�%��ڞ�畖�!&�1���1�jJ�����-RmO��0qu~��a�fE��F�~q��kׅ��� kWX���I�Ȱ��zXjD\D>O�S$в��WG]F �o���
�g��s�Y���C8�']��#���.��T��fːA�Sz�X�v)�=�~�i��X5/@d�ǉ�3C��ت������a�+P>�G��h��Y�|��6{��"Z{j�	T�&�R�K� y�G�[��1��E�Q"��$i�?�S�(mt���) ���:��c�}�a�1��f����h�8�p���h�	eY�6#�:G�S�Ў��>8�>P�Q̫�H8\��e�B�"_o�D�+3�$`��'��P3t*�?k3��ꔷj(@{�� ��4m)� �P�U�u��'&7/0Nr��⣋~�u���ظ1f�@�}5V��S#���m�fg6%���qr�J��g	�g�ü�����r���͵i�wW�*��%x2�]�cw�Z|��Ϲ|���ǌ9�c, ��2\"[�{离����)T�S֞�1�bJ�/.��z�y��~�8����c����i�M�u�HҦ֓��8����Uy�LO�"�-�F?�H �����S⡔�}`�� >1ïh�����!�����ԡw�r�]~n
��f�S�=��	�(�M��g��U*����E;���u����+!�_���_�w��~��d�h�����M{�O�8�G�BؼPԠX{��3��=b#��"�5Lh"{�����6nx~�(iQ� ۴��l\Hۗ�c|��o�
�}
�T���{X+h&����f�w`J�ϻ���[��~��bJ��5�#eQ4U�ޝ���7q��m�1���8�q��߼q#ѭB����MC�����n����|$�x#c�Y��_�I&gHdu�ș`�wdF��o���#���r�TL'%s8�k��q�/�v؏T��f��cB�8H�+�5�JL8�BQ�	2'�����̍f��I~�����N���e3��b�;�����mR�J�X������+�
~[,Fq��'5�s^h�Z�룇O�#�Q��`�7�����"�}H+���.�����`Mr{�>�@�c�bS2�;A�[�۞Cb��Z��o�����9���ɏpQ��R���"���h��";��s��o���V�U1�O��e<����Ćc�N�D�Y���?�t�%�L@R7UΟ�5��U�2�����N�&��
U��Q�Pu��<�[���IL9Ԋ�m�qb�Y�c�Y�Jӈ�7Hs�3$�m��#h��\z����)B�2EQYS�נ�?8ܭ��*5=�C���GFzt1V,���J�빤[��[�j���!�ë�)n���l2�(�ܰml2���S�Lz�-�~M�m����w��ԗ���>xŁӬ��R#Y��!1��WCP�������i���`<(7MR����G�6\���TD��~&4P��������p d�('4=Xߐ�X��V��5�R�a�Jn�h���cZY��A��46��z{@�k��@GD�����,�����b�1��0����$!��W���4*����fN$L���*�A���-DB��e�R��	��l���z�u/Oi�7a��7�g~�rWYc_{�Ȩ��*Vq����/{a��k%ݨ-$6��?��'�[-.����D�D;u�>n�~�a�o��$.�h��޻k����p�M�O��/����j���u8�x�i�"�:��H+B$�Z,�HW�ʑ0�r�:Z�1ut���TGВ� }�Cռ��:H+�����6�����/z����JT��@�R׀��3[@� ���<��s�q���ix.޻	AN�%c?��࿲��jp�t�w�fP�[����C�_���D�/��U�]����=��JZ�7����n�� )���l̋��H��*��z�M�M/Q�� ���������-�T��
�,@|�Ofȗ�_l�g�H!�q��Tg�\�5����+����G���u9\R�G�����
Pɰ/v�Æ�"�;�H������0�̛���E�D6��#PS��)q��Is˰���tCS���A.2':ڎ�9�S�do�4p4g,����/�L!V@�[����\+a2���*���S!�N)���?E-�@����x����ep~h��-@~���q+�9���x����@�����CVDo��L�*�R|�3P��/�E|\zv�58HNQ�:�u�E �c�!��W�/��D>�ҹ}�����<6ta�w������f+R��@��%ˋ�9��1��g �l�2�q,�1����RB:R�.a	������%Ӆ��S~��0��"s���bH~��+�BcT+K��W��'>H�%{���Ͷ���]��Ӻՙ��'O�"n3Rikq���L������E�zbn����ٿ
y�tҏ�=�U�[IE�t�m$���K���<ӕ5Eڃ���W������y�]��0�^�V�?nZ0[Ǒ�n�p�ѥ���B���5�8O��Fs�$5{�笝��� f��h�UP/r�
G���_B��K
w[έ���B	�`���R��{KO&�r�"'�r����m�qƍGSo�ԏ���� ����]�e# ,�b"�]�i�Kv�O��`�B�Ye|A��,�ٞ�Ǡ��n~릧�x��Ä��o��䂪i��cn���dc%��˝��s�,�&�zN I��e���5lWy8�˓�1L��e~�Fi)]����R�*
t�7h��Pl�7���Jr����`�ݭ��g
4]�}�0^_�]s�9��i,6�x[n��R��� D���C�KÏ'G)��Q���/f"���*�������h"tw���qK�%B�.~���翣%1����Ή�����ל��{y��Q�*6yЙ\i�A�\�z�������h�>v<�@���鰬-'n�.��M�E��}\�5ata����߬(�+t�� ������y��6��R��9��f'�G�7s�5��xMn���L�� �����{���}����s,��Q~7�?t.&_�.�נUd);"痃���4��EL�ub�#9�v��A�W;����n�Y\z�o����� (�?4��.9ǉ'E���h�yK$��*vz'%�9�+� ��ÝU�7]X^߅����!�\���%
�4�|�~}���!��3v:FB2r�C�'����@}v�l���<�^-�%�����v�7��U'��iP!+�h���(v������ԧ�C�+ٙݓ��Y8K�|���{���Ͱ�7
���uк�
|��#}6���+����A,!O@Bn��*�m�������${���J�ֽ;��]]:}��= &H?�y�	ڄ���ky �5�*X-�W}�3	q_7~������7�\�.\�X*)���� W����{H��f��ȁJ}��%�vYΪ��\���O�u(������қ�8�D#|��}fRo{���l"|V�����זF�{���?�9C?X�10��D�.�Ҁ�����S�Ha�xh���P"��G,5_������H)xf!�y��':�����\�K���qS����p�z�3�퀠���K�&F����G�e��eDμİr��JEڄa��}[����=��@��p��-�@K�z� �W��d����C�������H�P|�ʹQʇ��w&�V�q����@M�1�ce�}�[����2�3��}�@q�f:2S�(�����znwn��	��ꫫ��d��VK�iҝt�(�4�r��~�"�<����J�)Jud(��9�qY!8�C����B_�h� T��F���x"M��aw9UU�v����թ
�����oŮ��9�VLW��*��]+$��*��A����O�FC������s쨽����)���{�����#aG]���t����8���?�A=��+Lt3��`���~�
~�^��Y�5��)I'�8�. �;Ņ�&�ۮG�X�!�Y=�������̇<�f�!F[0�l�|��"<��88�a��{{�j���Hc�c����c;i�?ֻj��k�G�:����(�3��sћO�H�W�s-ր�"�&�2����?�f����r���tqt��� e]�K����3=x=TO"��E���:�ŉ)�r,��Ҙ8�iƸg3��
�l��7/j��+�
&�0�ۑqK�F���4�@��~�"�eج��K�f��7� i��3����d*$\rS��JW�f�4_���A���zAQk:#����@�>b#��F�����:,w��v����Q�|��m��9X��A&��2D���"�Y����f2�-�w�j�ih!
�K��#Z�՛8�ET>O27S�����
�� �wh�����K}y�8���h����^�5����s�-j��� �c#�c�è�&����y>���[ϫ���m�����	R3���&�*+���U�4
��$)�o#R���6(�[&�!�3�Ӧ�Ah�a�������5R�x�A�g�bI5��BѨ�2���hɡ�-�����#bc��/*&�~���XK��V�{5�M.��SU�OL�6W|�yI�G{��Ĥ2��	B�\�Y�^]11�0L6C��#����_�yB�>9�1)�	)�I�H�9��X����#4Aj/Ɲ��)�!Q;��p���*��sD,���v�E�lL{�珽Z4�=N�����j���� �50�Qw}q��Vz��[�;6m<�!5	H��]������|����F�!p�f�ϓ&���B��C���\x��;��S�G�+��7����� `�Q �k��B�;bn�14P����[�k���^�}w�׼��x�a�Xi!L�2�Db,E�O��F�w�p*��v�����
v����hZ�9^䂹�ڗk�	����3�9�����{ٗLNm��p���K%]}�;-��qסΈ����Ḓ��dN7�EQ0�mH��d���!"_h�{ؑ(."�_���x�H�MkQo�"PG�"j"Q�IO�ֶ<�#vd����)r�y��¢ڣj}B.M�6ƪS1SYL��-��.� �ù�.L�22_��n��$"�!gSF��e�b�y�H�eo\�����S[���Gt`�Ʉ�S�0��y��jPo�A&
5C��L��CS*��O�}�3���8��:��IG�յ�X�R�\�!�����C7�������O�=������t�:����S��#��a�t^�n�cWz��f�����)f:�k���������/M�+����@k�a��eÿ\E�o&��c�[�F[�~�Ү5s%El�x���0kw=D�l[�g~Cy�Uͣ�Y ��azg����f0H�h�e�ޅo "��S�W1��a��^�\b�J��\������2\)@��Dt@W�Xˑ��2��Ҕ�z��҃I�z�G����Y����d�Z�E��F!��i=��`� (!O5o�fcǉ�3�!#��-dG�ӎ�6���c��{J�����D�s�i-�mD�k$$;��X��B$e+�[=��������Mu�a�&p>����@�m�� (z��e�u����,.%Q��.���66C�>+�	H��b�H�*!}+q�4u�KS�.�[��1hK�43��U��̬�)0�3،"7���Ms�/H�Q��˖�,��4���D�D�7���O�?�X�E+<T�y�b�XS0(]#���v0͌#��t��q���gi�)O�/hQ��`>N<��ǀ���ͼ!�T��ݵ�+���YJ5��*�=na0�W�QuŻ��1`��Ґ	��)���C��b�y�'[����8�F7�saF��Mc���̑��w�Q����^1}Ln��U���c�[SS�_��R���e|�{ٳ�N�]5H��!H΁�f#�B�<3��n3_S�]�.C 2?�����0���d��@n�:ST�AͥL�|�4�W�l�Z�/G�r��q�
���_`�����iӈ��Id(��y���Ns�%�pY�g�.q�3fm���K�(���R{9{�*ʵ�8�����������(Cqk~z�PZ��M r�l �&�>��N�<�Չ�*c�Gfc�N#p���բ�PZs4w�;�/�(ٚ��сi����*4�Q���K"g�#0e���!��ƶDRǞ�r�Z��m��xU�_�Am�N簻�μT�}{����a��/���͜�l����� �\�[�	�D u��mXNn�H�]�^����B��w̃4y�ףg�yD,9���)��x&�o�\(�������Y��3�m�LG9V/�a��3꾽�\:j�Q/;�q�� gL�0�OB� �Cw\�g�]s+�D����W�R���k|M�o���;��YY]�C�d��ɋ��L��%�-Y3�9�3�%m�����l����9%䗙����uʰ���H�^r��QH�0X��(�v0֣[�(��#����C�� 2Q?�_��ݳ�P����DLe�O9Y�,��4w�UjB�C��҂�b�PY}��[qӕ�����}\@�H�J:BEN�b�>�o�o�8�;�h���.�}]FG}ZO���n	�V���ME9���c��alP�W$K��j�D0b�He�.��ZPK��ڛ�	&��K�TGX�v�2w'%	쮍�����9���r�J�����������Cćo�j;� mt~���R�q�>) v���_$J1��� \����'�r_R�^�Y��T#�Ͽ[��M���yi���$�j=(�{��W��֛:��ID�6��ʙ�3�S�m�ˤ���<.R�0���k��nt��MK�ۑ��3��znQ���N��(7
p���D�����U����ܐZ�"en
�����T�������-:�,n����� �d�UO���:��T4��4}^�+5s��,!B�^�V��!��M���Ҹ��s��t5Q��g�+k?�=�
��e#�7��zr3{��?�O���(q�h�D�+]@�e>�)4�p�HV��~�T#�ʔm���;�M��l��@v������6��!\G^~tFbf��H�V�����ȁ��9��$��]��L��ͳ�ր�5V�����>��Os�9_��Z	5э�Q�g<�y���]���<���C��F52�9@�ꭨ�O��>�Ǩ����VZ=o P�>m�JZvú���A�x��W>�VS�Ⱦ���C��p.gI6�n��v�����H�X���Oޔ��`߳B���W�{L.���ZlN~
jX�s�"��P'�&}�=��OЂ`WQf��NWVo݅��cOѳ�'�xcŊ qL�HbO2'uv���e���c3ok1���Į�|
z��.��Ht����T"y��*�[�� ��g'�?N�9�@�<��F���bJoW���>P0��w���RH+��sZ��E�����|q\`�S^�k�R2u|j����v��.��\z����o�BwO�E9�i��*!���s��ni�RUB��Zc��^i�yy��}���*Fz�\��d?BM�>����R�$Xu(����U�p�S h
�%W�*1Zn������0V�Pa#/�Q
�Uڌ}-P��u��7'�<Q��X@ZQ������6�6?��e�vE�f�g������5���wb{�����{(i""\�^��w9)Tn��Ʋ�&y]���p��k�" z~x�Z��B� �TQ)��k����sLL.@rJ� ����t���S�Z�뺘^1�zO���q����0C��&V��ES�Bn��	�ό�E47��6�<'�P���� lx��q��ޠ,h�ҿ�������ᓑ�2������p�x�Q {����s���!�ou�B����z�-aԗx�pb����W0��|��TgͶ<�تe�oU)جY�.L��+��;��g-��.J�-���?�3���*>���S2!����\t�{��/!��f��&	�Fݕ����NO�[X��eS�:�>��bm}T��G�຋�jDP2�@w����5�E��[�S�W�2vT|4�C�_&^�G����:�'|=�d�Q{��Ig�4p�Ou��ڰv��C|�O��w5�8��^[+ܰ<:�{�km��J�	�ÓC	��������ǜN\��c�#-�v��!*5��Ņ����Z���WG��[�]�L�������Ǥa����%0*�8�T󢠱Tf<�./�+Y�	�B9�c�ev�%�;S����7��iG�%�fyp�#=/`���!�1(%��-�,�?�[�6 �n%���U�J�]4�j����x<Sm���=H�i��F	�#��!U����gU9T[]�7�������<V˗��	q/�ԁ˴�4�Y�$7�,g
E�Ċ86ծ�,��� m��Ne��P�/�2�i�y۾��#�S\.�eY}�`��Fu����������G����_��|
����3ˬ�P�a~�(h��!�/��U�ܲ5�7���2ѷ�oi*�	gѦ�A�Z]�n
Ƚ�D�n��a�9��
���iT6��FuAd�m��#i�/*�>�UT���0g�����DQ^ k@5�X��d�vsպyT�3��7T����k"{"Q=�IjL2gd�$?�`<��� %����F�"'�Â��ţ�S��]H5a��b����~v��6��ܺn�R@�#��
&l|�|mc��� M{L�%�sR%�ޤ��g3Y�8�|I��]~�����fƛD��P$~ceb�X���'f��Na���b�K"�=�=����~`E!t�@*V���7��^�(�Y����0���H�UHJԗ�Lj*F�����>$)�G�����A�\,��.jNw�t߄���"��q1@U���iº0��0m�M�Y��p�.\9m �ܖ���ŵ?WqW��LB�� ��9�3\T�&J����W[k@�WFq_��	�Y1.$���j`KC.��E$��T��4���P�^�]�^ )�W��[ӏ��as�+���:W����N��|���i��q��@pt�z�I���IH�����e#ӶՇ�Uuk�P��'����D@����%�2�������Ҧ��V����N�6�GH����O7
N'IV�$P�MQ��A�A��O�|cm�L��G����+�����g�o^0��KM`W��-W�k��M�nd���~x���#)��:��~#�ܺ���x潆P3%ح+�������K�Z���I�K��π�{�����ƣ��up:ʍ/��B4�j!�&1�>�JLv�~ĘeM�E�e>�j�!Z�h/(�y�H��}�_���y�P�~����#=q��<ݾk�l`C��t�[�(vK���py���l�d��{o�%U��CA��&���!w��JMk���0Kꓮ-�!O,����n	L��Z&�IF��ߞOj�t�C/c��]�[����R��?Z)+��&L�C�{��>�d�Alj8���*'l���ԝ�~���wl���h�;���ǚ�!j߿~o^*�	㴑s��H�Uw��/�b�V�Sя����Pa�����RK:`n�_���`\�#�l�bP�u�+
)g�!$A�]= �hM�Y�:��1���J ��/I��Lp�,ɠ��-(�r��x.dm,',�H-�(�.�O;�
	� ��u��-�WB�m)��įϊ�-[��>��vB�����NI���=it��7�e%Э��TUz���
�"\��	��ۦ�	���v����N,�?���yLԫ�R�6 ��̷�PP��2�zΘ x�
N�W�"�⾂B��&�H�8���2�S{S+5�j%㺲ߐ'���"\~��x2�4Dt��?�$ۙ��,j!)�P]単�⋜�4v���r��p�tr"��9��d�����\�����c$���b�����B��5N[���⮒�R8�rv-J�����sBE�[~���W~�r�,:;/'�5��9�5�\�Ǚ���vjT�����$���x��I�����ͫ����>H5n��h��C����m�r�"l����"1ʳ
�'f�y}�_tMg����vy��B6u����o��B��:��vrG���m]͡��/�oXU�_�G&+�&$S�!nEv�����\J�ȼ�R`�Ǵ�"�ޖ۾7䣭)܃��v�F��y�"[&ΚT�g�4O&�R���_,��=�ra��:D�i!L2ȼ˼"q�D�ඒ�v/\�Ȑ��a:)����;3����r0.����hw�sO�5����F"��"сf�?��mb+�鿪ϟ	�qMc@�q��y��݁Vj���u�PVqy`�2��.�)Q�ǔ1/;z�	�h��"�V`;a^h�6NT�s`���ݵ:uT�P�7��L]z%T�dE�,?4�̝��C�K���JPx���5�%�v�"	�i,U��ir��X�2�^�^��IҢ�"�g�`��2�l�&�皩�v~����� ���?���V�:�}i���ce��8��[����i�iƉ��?;����'�:�۴_�-2��6r��������֊��aⶇ�?�s����b|.�����z���)�bb���@NʧiےJF�" ��o��r?	����2ͩ���[1������ Cܮ�ѯ�����,��~,�g�Q:Z�D��S�BS)�+q�1雷�!M�sn�X6�{D�*�μ����V�:�2���S}a��������# ���8��r�nWk��FiE�xuڟ�#���V���s�`F�U��5X� 
������̚�o��̕�ȋ�M�������Z���$6T����Md�P�(ե�0)r����ΓnJV�=����(��0�N������O��+h��W��SvH"�%��lP�iQ4���s���5�����|lu���a��lQ���ڴj8��}I%���ip	�6]�^�?�yK��ɮ |��rw4���`Sxv8Ԡ�Y#��G�i����zhVj)�8}�,V����TU"$�z|qw\N���P�PD�Ĕ�b��_)�f�dc$>X?Pi{V����{�jȼ����e'"$q�ę� }/Xo�K `u��#$���_�"d�����wˤp�?��
ZM���8�3� R���`�Rz�