��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0���l�=�&�D����F�n6��"�,t1g�Eo��g��mb|�c�	�l{�ȩP[��K~����"i�stɠ��(�F���Q��������b��y�=�y�S����b$�nN`���ӵ����[��U�rkc�>�0�
�i+�Sv��T�`Gޗ"��~�cF�m��arR�@
�%����{~����m�~h��I�a��H���$mx ]��>��lZ@9dx�'�AeV�.W�˼�(�G�2�q%	�~���Q�NJ�1���h͸1���,&�Ɋp�N�P�|;%hH-h�Q٪1��\l"�aM� �]l.�j��l�� N��<�h?p�';%m�1��$�] @	��b�ݗVJ=FV�6L��X�����V�A�w'�T8JG=Y	���H�&�{���a�+�:��/�N�&�7�iFj�;o���቟s��N�����O�sos֔?	]�v���h�漙- ҋ�R������9���w���+7�s��-�rU���{�ֳԯ5��F���c�Y��T��s4��{6IS�~OC�V�m����$Ǿ��}kW�é�*��V˼j`7�T����}:<T�NOY�`��k����N�4���s$���{j�:9f�:�v��G��U3�,(���~��C�"�G�?���5���!�>ɔe�s�R��/Bg��"?��+&)��LK�:1v=��0�8���I�?״7�Q �FeEУ�`[)�/�v�����&��\�\!�)��]�ܘ(�� ���P_w��]���C|�/���%a�wG�����필a�~ί�|5I�Ae��y��"����DB�¦�ie�W��l���s{�;�x��o�;ڦ~����5@=��Jd�P�T�7bA#\-@��G0n��lz�Rz��:�pvGs�ή�N��S�����=!��_��6�ϰҘ{���\��J:�w~�7ߠ��IG��˳j�	Gz(x	Z�0��=CR�"�0�H�t��\��~�S�p�xn�?��1��G���}�[��@���ԥ�}D����V�ǋ�y$ �j��h_'�Z��ѓ��jv9�P�׎w0S��/�ڂ�:�͊��f��V�[�����3����`&�w{
�*k0�|��b;�~��8�u�䀰i��tӷ�S0� �!.��Nh�rq6sdꢻ�n���:x鐷Ѕz��f	�ۤ��\gYpv_����=��Bm(޼��T �.�Drn9D9��7˖�*r�`x�`���t�����($��g�@�:r/i
Y�G���뽃�Ny		��`ӊC���$��2X�z��#���޽#K��o���B�6��i\?���tT��8��='W�ې�zL+� )x�A��������V����erE{�G��ixK��+Ȧq9X��K���N��)�`�M�$hh��V���y,uȧ˲�Ǣ8��G���ϖEo�.�ݕ�c�#�vr:=�{�qܸ���P���L�=W�^I&}��N&m$#���O~�lCQ���՛'D#� a�C��lt�eJ�Qw��N�gh��(��MF.�f��h��5X��S)۱�v��}�D,�]�%y��Y3,��2�,>=���b����j��R�F�t��a5zր��p=ob�����Z��oO�ͻ9שM�u�2�sy/��S2���Bi�&'=��1&F����NN8n���C4��Ƹ���$���N���2c�8B�2?^b�_��0��EoS,�`^G|a_�i��܊)�����b)�zl���:x��2��_�j�aC�m���ؒV@�<�� ���q�5��S?��
OF�yR�$pm�S �A�a��"���I�Ti����N*����.a	�,��觗�&�̤co���X����Vyʤ.v*Y��[�U_��#k�+�%�)��ʥ���s�+���c�{�2�.b���9Rӫр��*IIEi��+��-N}%G�⍣E���zՙϣ|��F�M�7l��"0٩+�1�5:YH~��X�g�����&��4���:P�O���}m�%3��hd`y�^�B������Z����"wY;
[ꀔ�>	3�//^aaq���	�}����R,�垑�o�{�)����Beoq��$C�s�֩5��[Y��yE#+@�3s�H���H�C>\zS�l��H�(yq�2���5$�$�<Kh('�L��n/����ȳ9`a���8���	[Z:�P�b���կft0}^ϫ�ҢEAo�(���"�Ճ���R`6��a�uR���\A�`�����c�i�(�u{D���4%Y�1���M�z\��S���=��
d8~�_��w��?�0_�w:.d '���%�e��c���;�5��JG_��/%k��6�sa�4� �>�RyӸ��+g;7i�<��8�Ѻ#����{��Vh��/gE�vr瘘�b�r�fGsE��=�������y!�/fKׄ�`9��2������qS�L�h��iQ�68���ϱ+��,����m�/:�	Ҧv�)>_�$��~f�pg���s�ِ�o���N���	�|�Qr�ݘ��!���Y(N-zoF���J�������S�H9��M�r%aĝ�Lfƿ3eh��V�<ڛ��0��4��ѺW�)_%��� Iֽ�^#½��O�s�2�����jm9*)6�\}������Bh�/�>�]&�5w� ncpV\��s�S����R��\�E�W����sg1s����(�P��6��ʛ�)_9\E1���>����xR3�nGn�y���C4T�,e�R�ĘT ҭ���x�����l;҄׊��Ɣ���!�q��i] �4���_������r-"$L,8�����+���EigJi ���xŹ,q� kî�#Dz˥]m[��E�l\F��b+q���X��a���І�!A���{ёG"�.֭>~�I]~� ���i���k��̫vbGM���0�X��$�o�$���q�0
�]�΅��m���>Y�+�Š��� @���H~��0y�T� ��AE�z5'�<De�4Ј�+J|��<��~�¡�7\9X��ꣀ���I.��T��P��Dl �����	��I���������=x�+��kϝ��W&��9�����	麸QD~�[��5x�ۿ��fI��po�,��{LT�󜌍�.�_'�6����G�P���7`V�ɇ��=��r�-p*_�<���ڴ�8m	�:ٸ�Qz{:g���C�c8��^4&]P�#��ؙy���@��d޼����e���.BH�B��V��7�ju���`��+�����v�=LƝ$�7 BQ�V;mCV>�`���AxZH\��͂���{�׶2�w����[��D�]��J3X�+	���&XD�9�L=]��n����X��J�r�C���Ͽ�7���u���n���f�O� ����5�S�<F 5�׵��:�5E9����z�|L�S�j�
�;���;�������y�*�M}�
0-���K1TW�f�Y5�����F��gh��
�_��é��%���r��C��J�m�kg��epft��Se~؉�=��`Y�{Z�V�؜H�g�c�|�S"n`����g���Db���t�$c�`i ��q{����*gl%�X���������Ϝ�e*�b�'��7-�2��d�=��V�
���3��^U�R\W|��\ڲ6��L+�WT_�� Cgs=+��ňF�(o�,A���7��C�}����z���#�_cD��KQ׆��"+;�p[��}��բ��n?���;/�_M;�y���	�T$���|l��p��%��T\4����ʑK�}��A4ς6�QO>�]=z@�
Ү�kB���R��O���/l��VVۍ'��(/A��¹=�)X���B1�\����)μ�~*s�(���-N�9��ä`�9Z��Q�R��G�!�@t���b'�G�ʁ�h9'�gD��S*�E���:m�H�^��^��q�ϙ�f�a`K&l�����>{�H��&������"L���0���]M�p��������7�s��O�.[�h���sSq�������[1v�2{���0�;���'���$��U���~�?�2t]>0Cwq���-ы���F���.Ⱥ_
yK��9t�i)����L�z�t�]*�`��?���O�~}r��Y��c9n�*~	
$*�br� �~�2y�˿���3��1�e7��Z=+���7���`$2{�r3-��c���BL2�V,�D*��S�s�CWt�V'���JЮ��K��X��'�+��O!c�V��i�?A����!K�e,�Bt:C��Gԧ���b�!'��x��\�� �Z��P��,�є/9�%6�٨�x�o����Ɵ�EH����|�k��U}��`��3���6�?uUW\ރ8y�5Z��ΰOJ��TU�Chj:N�(�f:C� �!����8��$t�����h뫛\���� Ԫ��\������p']�-?��K�j��1����Ҭ�����x�6������c[@��[7��r�����K���!s�C8[��LD�2(�.v]���پ8u�K �M�l��k����n�*%����h��7�l��� ��k&$Ϩ�c�}a���T�S��iݱ�/q��"1Ě�&x��>�ΰ��2¢:
��/ǁ�Y�>w��up���+
{3��� ��������d<o֖X ����W�d� ͞��^���&H��<uc�9��T^��	_a�n�7�R��>"/�ؕ�m[Cg�K��[�Pzf��B�Q���g%��>Cϟzx�.����g ��W�=kV��O<��X���&�Y�܁�
��:b�/���-7?��������pP�)KҤ�~|IT��
,f��!��7�;��ڗے��Ϯ�o�78�mHW)�#x�sT�)4�%�h�0�\��p��|?&�Y�U��2�nG/�v��r %]�i��$"��ƀ*O�cm�{��k[\=n����ɮ",'A��)��$h� Wgyź2NE��$WG��%-�8��L��IjcB�}~�\A����4���G˟\��lɅ��Y�'6v�)�Y2�%z<�k��Kfot�z�:�ݾBL��J^@���"&���;N����;!�Uqgc&�L8����=Ǝ�kx6H���G��TF5�Hh'�f�+f�~�H}hp��N�i3̯G��Vq����_!h�B!��<1*w�Y!�f�ށ��.�S^K���b��
0s��o)�I��#n��FB���ok	?B��uj:��I�},���@NT�@O�}�2.�ʷ����V���Q�iǰ��hi���9���B+��,��T�g� � �X.�uh���
2gdq?s�?w�9�Kݧ��ց�^H��P��3��H$�G�Nv�r�[�<����9��d��A>/$��F)���=w�w__Հy����$?[z�f�����BOʞ�Ӕ�18�Ȁ{V]C����F�s ��r�Q��s�����w�c�u�O�=��|d�V����Z�"|%r�Y�����*Y���6�������V���P��^�'GE$.���s�!=`~#' �P8��w��噍�@gsJ>�Pw���5 7���*Δ,&];�j�v�ѵ�5��q�U<�'�g{R,�hΘ8'���,z&թH��.5���:r���KG󞞋��`[�#<�D��5��5��s��W3/�B@�}aTsZ=�=[ ½FNk�UZ�6�GE�%f@r/\B�k��˾`�H���gm�X/~��V>�1��h���}��3kl�����
2,�ecG���e,�@=�i�ztq��Ķt��Xb5����	G�P�3ﱊ����ݩ�ҳ,?�"4��5��O`��k��R����Y�1��F�v������r��rh�Ux<!�s��N��#�$^dC�t�g.r0^3Ŭ�{�xD
	�{lȠP�^��0[��qҋ�3%��$"(ڿU�ݣ�`6U�>H�xF��b|�k�{ Т�&BY�Y��7�Ca��qJ8V��Z#��J�2��@G���ݬY��5u�^��#���"���ʑzIZ �G��\ X�����G�+3�&��yS�r�g3�G	���2�P2Z��
�ZW�w/"��Y�|]�)�BW*~���7U�#D1�Y�V���|�\�0��I��@?�+n@m�v�$�׻m�=V&X�rc&up��r�ob�,9��˽~��"Eb@]?\β�2���&��T�g�ϸ��ԩH�o�>Y��Q��R_Jx���o�',w���~a���c�tAWފ�QTq�g�^�Qq�3yKF��o�r�=1Ob��è���/���O�"R�����-���߯W�:W��i�O3��]���h ��ö�f�J�j�m�"������r8p�?z��,��:��H��@�k�:�q� P�i>:�O��H5�yL��m�o<�<�L��Py�RT"jȵ�����s�I��"��2�'�Q�v(|!q�9_����a�m�;��h&5(8����b��d'P�ջo�i)�)/��T�l˲�lQ�'����DGp#�Ө�,�B�� �v������Ztof_�����zP�/��R7��%`�ܴ�ΨL_q�4�
`��e��df��]�� 4I�����6�__��;Z��Ð��5��a�C�ECyH�8�5c��\���������'>4F�mI���V�*�l��� M��Ό� N���Ygk��S��IS+�%���a�Ed�� 74~w�1!�����n�7��`_?��J�b��n�S�C�S��mk�d4	�����I$��w�\i�b���<�ϴ;� �s�����5��9'�J��,(iN����]��"W��Wݜ ��1e(��}RZ��{H���@�6��E=�+�꣙��viW9%�,��N!6����{]Ք^���d��b����
��)&�RS�V���P�J��s���):���(�IN��nF�5��J�T �y�Q�I���:�?���-?�v#��9�G���&&�iI���� tqhn5t�Y*��	Ce�u#R|�m�ڙ�Wn�uJp˪N�.��s�O�qb���!夫~�V�I;h�Sl&��]زm�df�&b��ѝ� �޸X�?�?��,<r���	$~Ĥ�<x�Ŕ����p\}���$��}������~�m����p�dg� �ЅI>p���t�����!88D�VIU�%Jy>�v��<Pܸ�I��L��s.���CKX���{޿2��s�et�Y��%x��N�[P��V��F��*�f�͕j��\H��hK�~�Rd�`(w�}��̊���b��p�L��G����0{������� e��\28̯�cg��'*�f���8�I��q)�AU�_�~�&�K,n=�A������@cPŻ�~�qa�z&&X�.֋x:���l��ߜ�|)߾l��'���pB�E0T3'��O���'f��PJ��ͥޭ�苢��+�J!f��e5b}��HXh�3�����~S�#�p��+�J�{,
G���(W��g�A:	�}�d��C�G��v�M�#aU-�G?�j�̤7��%t���$)�d)�ڱ�o���Ez��lO s��.u!қ�Q�O��>��կ�G�b���=8^��	���5c�V���?�0:�J�uIk��9���m��M�|�q9	��C>P'���aÿ�O�� 23m��צj�� �HD�-sl�Y�:�9`�Gfq (O�qt'�����XJ�Z�wEJ7(�7F���t9����͢숱/��(FN�S��	⮣��z-�2�e�� �~���10�еG�!Wt�M�䖧�ч� ���V翌��W��Vn��t&��H<-��$��YP�&�L�R�BD䵈�Y�`�D��%����xQ���W����;mz�<�G�ȭ~dhI3�7�PV%Z��G�J\��R'��4<dc1םD"��_��~��»r�"�* 8l/��W>e��H(Z�&���j4Tq����4r�ƣ/@��S�h|�)���;�G3��$~<�x(�%*e3�)���|�����P&��"�a!�h���6�C�DL��M�=��Q��d�:�TU�\hy7!�z\j�R������z��]W�iE}\49���O�9-�cGk5�.68����G9���X8�ɺ��W�^n�h��%�{Cb��I
�q��M���3}č��W����ub-�&���+�{*��J�.@Bq� �����⯎>��eiƕ���<�]�℔��o�Z�����e�fm%(ݬ�d���$0�I�źi�K�s�8�_�1�3�K:=`�R���ƻ���[,91���2)m���_�o�\"��Vr���(Q��4����y̑{��K�G�h�V�m��OtJce�����M]h�%��o#�����~�������Ű��xƛf��x�8�����͙�������VP��F�99��=��'&��3�&i����Qaee�����ص
��]V�pݏ�-E x*ny:ur��%�!��]ⲹM�t���0����w\�v�@u�ݤz�}l����e�V�Ŕ�^Dӣ����z���> a�c���<����=`����JsV�T�J.
H {ބ�.�G<ѳ��z�e
���-��ts���%U�uD
��r�	�Og��Y\%m����G����:����b�`�a'���v8�r�ЪB1�25�u��3P�BQ��d2{�bX9���7`����ic3�a�z]��)��tD.b��Z��������~��V&E*��%��s�|W+v9��k:�O����tu��-ȩXFN������mu��3�&wP����f$����T7o��!��)�����k#b�ߒ����G�C �6.)�3�:��7�#Zɭ���R�����d���t�`?�=6�я��`��~)PşF�\�C^��p���j�f��D
�q@�;#�){�D9Dp�W�|{`�s��mE��v=�}�����Y�v7���9~��z�
�k�;1�HW��N��@0�NO�L��C�]�Ԝ��A�X�2݋Yt� +�n����q�kq&�k>н�^m?s���oS��}�.�x�KZ���l�\/�0���P�'��VM�Uwv���4�08���F�;�ʥL��8
�؟���0�ᯆ�n;(�zo���6�l`Dl�}��S��_�/|FIy�t�9$��c|�X��=m��B�g�5�R&�S�W�7��@���A�C����˪]�Q��L�q6c�L���Ii�\W��j~�D&��}1���.[�ˣW`��� ˞�r4l�\e@7��C9�z���2�GM|I@�q�:*a�Lⶎmņ�W%Ӄ�y դ^Gwbx"w"�'F���b]:��~�;��<CJ��S���,�3E�yv3\�����d�2U��q���)(-mP��^���h [e�.w*؅c�7ϝ�	�3��S/�|)�i�dn��v\K���^�"J6�#t�O�5�@ �i�V���c���ų4�a�A�3�ˣ�>��Q�p-�
s ������ԄQw�zƮL�ĺM&��I���l�g��ǇO+i�3��t6���������Y�N6A�|���8MU�W%�P�s�d0�(�0�&��4�6�7P���`f��<|� ��*ǖj�LX�ۼ�?�(E��1������6�O�K����1%wO�y��� ��N�u�)`�<H��|P��u��aI�5ݨqk]1 a���p�X1Ԥ'Jh٢�k��$)=kIK%��p�6����P��
,U�p�W��C2@�.
��'��fi4�����8�mH��ܭ"ߩE��itt�9���Պ9T��B�
~�sd=g���!�����Ag˃���s�3a4.������R�ʆS�c: ��S'pĔb��\dI#z��m< �:L��2���)P��!�EY�U���~����j�a�3��X�|�-�fi1m������)���e�$Aף����Ř��V���g�t��s�����]�}Pp�_)N�:{�i��MN��V�,��ޒJf+�흒�{�{��G���c/�.N�A z,,df�V���y� 6t�7�'�{�T
��K�$F�hگ�'�5n�� �[�Fݳ��)/�\n������E�s����JaV�����	��LK�o/�(������M��}O�	����I��A��58%u��4���@]�z��73W�����(<j*��CE�(4�,��m�S$Y��_���,ib{Z���R?,�������ٕ�q�������L�ll��|nIt{:�����,�E���$Q����*�`�F����8"Ӻ��$ދڽ��$�������1��#X����Сp���蔖��PkR�j�-e�u��{f`j�J,�p�CX�@�dp�n�����_b��7?S8S�����i��[h���zza��6ӎ����QL�dN���K(�-����.�~�N�����/;0%��2o4���P�<M��3�J��S���5��)��p6t�$�K6U-r`Bl?�R�s� ��}�X]-�g@!���n��B�N�^N��e�sÕG��IF|���HL,i���=ϳ�7V^����t���V.�<V_���Ks*����-��BD����Y�a����W���(��b���0=ejE��һ[~/�8����ҿ�A�y�D\��1y�fֳ^��
�lI\859y�Q�xw��u|��j��a0|��T��5��ޕ�Rj��׵g�_F�T��k��� �Hۯ���7t|�L���]	���p��ق��'�0��m���M��)��qh�Ĳ��Q����O+Z\m�����6�e1�%e)�Y���X���n�}��ڀH �[@	�U��/�W�*��o���BS��&F<b���B�+�Q����lS!�|Hׅ\L�L�����&	�>4��Odg-�%���8��H�䴱�l���wɟf�?l��'����"\
!L zA�4�#�p�
�#�������p $f�����C͉{�x*q���Ip�!��d�f'���~�c�7"��,#�,qr��#��|@"I��,����~�c�}T_��΋"uN��Z�O˄U�9B!��t���{�6B��X�7R s��0�F�y��N�>�圭�&
�º��M��z���`=-���R?�}�A��8I����F��cU�*Q��C��])>�j��@a��\��%��H������
sy����&�r ڕ(�Hr�A@R�x:p�oT�0�A����ț�ٷ�Ŗ���/F���c~��2�>���Vz�h�����@kJ��_��[äN�>��g�&�	M�l�.����%u.$m'�WU��j�^R��m�����N��Ar�]{%���K	a]ګ�0�����*R��`}���{��i)H<��__l�����Ы$���ď-Q�mK�N��:j]�iw�X�q[���q��y�*��_�|-�nL�A��Py�������dN��dm*Ҵ߆�ujr݅�d�b;�r��c=8�N#a�8�_h@*4������0#i,qA��J�������ﲩ�S|�j�.�\�)h8e%J��"w9�b�;�� J���!�w-��)x�$D���Һ�> �%��ݵ��H/�ke-l�v��I��V�ȣ���ƪh�G#�wQ;���	��)����=�NF�s2[o��ڜmF���c�TQ�g��Ɣ�����T��q�o,� �V��q�������B�-ϷY�q���j����Л��_��A�Q��?�\���45�c��"����"w�>*ĵ�/5���`(s��ɛ�n��dkKÚF�"F(�n����(��?I��T1yt����-b(��@-fF�6�}�V�l^}c���R����qąغޭ�v�Ǫ '���� �:��:XN��nC<c�����Q���  U�)��t�˴h�g���h�J;��wJ�\�����A�T�ﳢ�hT����T�H[W���Ւ$�z�~��Kle����t���%6Ŗ_rz�D�v�/��D����H�d&K'A�Q��"�P�s�ǽ�/���Z�c�m~��?r@y��gcv��qY�sy=1�)`��̜�*����se�N���a��@p)i5!�Z���؀u9�{����ܳbX��"���P�trd-^�s�������:�'2 {E#0%��d8���o�=�g�Z�T~"r�� r��۱S����L�=m�T?����GQ0IfE�DtTM�J�=>>�T�+<���������!����lHػ[�_)xj3�JK\����:nƃ1���<��)ً��yų�^���PUÎľ5���*�-3E���}��E�]�����!yn@��c�3]ٶ5�*�@	�DN�1τ�[㩾x+a�@8s�5�X\�1�5;� �5nF����k�ړ86;9�0*B:a������5����)�ȜGL��"j��_?��j����K��J��8Hw�Z�4�#���K�=:M	%�`��H������\M�W�s`C�����J��fK,+G�넀54'��p�AlzJ�D�Q�4�DA��/��j��[�/�A-�yj��6p*Ԃ�&�X�Or�-�l !��'�'(��1��f�M�UĚ�Ωq�!QLc��j/��f�