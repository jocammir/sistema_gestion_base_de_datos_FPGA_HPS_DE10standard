��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��Nڭ�	�����B�#Z���?�4�j��0�ΐz�A�y�[��I4�fB���_Ɛ���-����B���M'~��k,���'zf���]A�� -̭���ҧ���D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T��P�]��h�� �x��ϝ�BQ�H��B#0P�s7�D�l�������T]����[�AzhӶ�����?���9�����M���G��j��Cw��)�Ђ~��c�ފ�\��+�p�7@�����?p���Ip���r\kᯜ��$�L���i%���U��/�&�sTk�KcBu�\v�����N��49y�G�8[�'EfB��'1؏�8�)���bgǘh���i_#����ml������2k�5�-7S�>����-�+mX��(Ʋu��O��Y�a?4ϊ;G�=�'����W=�'5�7?�9���@�^8���+� mV���P�� �=��������Hg��6��Z�@
�R6��Zc�fՙ�	��ߠ4X4�=KS
gV�Ĭ�������_�rGYۘ1?Q�J�Y��Vy�N>�[��Y%����(5�����n��3Х��A���3;�b]�t�O^�f����%�i�7u����K�^_�K<�nO�|I �ۚZ��6��v��+R'�CZj�-�-����c{���3�ܼ3���!�dƁ��,jG�ж
��	TV���i!�ʷ�{�ݤ��(h!��ocA���,��_�������I�[Q(Z����R���V����E8E�H4������~�Ȇ��>�Oﹴ>-g�� q-׻j�~�σl薍j>l[�=����;�-�@��Ưm�v{1���5��&=u%C�����T�@հr�˕QΜ�^͜Δ�ܶ_z3�c�xOě�E�f�b�D����c��;fK�>����kOQi�^�A��g�3]��' 0�Vn��sqpcSړ�sQZ��4�p�ǭ#z�o��]�pJ3%�t+��3��nUw��,�Y�q?��w!�`(�Q���Ȝ�~q)e�$<�ƜRR������v]�Re5?�+��?�	�2�ZBӞ���X{�����������H^S&z�J��%���5k��vE�l$�;���~��O>�,�Ox������U���VZ+[H��չWq��\��:W�E�Pµ#.��d"�z}����˅��K����)�͕~��@D�ݑ[)n�}�g�LY$�e̏�����M7"��`�������ґZ'CG9���JbaLy��s�#O���z���R�O@e�I��r��z�T��3��E��D�Yr8���\k1�*�U�9���ܼ���Q� �MccD�ᘥ�ʯ6 Fz�a��r]\�������7xܳ/��C��5���>��߶����q�]ŮC�,��x:���?޶��e�c���c?�r�n���1�*
{�B�h+moԘ���?�̢�?�h��L��+�����-���_¨�b�"��G�4
�U�m�.�U%��J��4�e�����[�0��CF��g�����77D�
,)Y�1?�"�	v[Rf�ü���M-�%x�m�G��6�HQ�<ocwd�1t~9n�A�X�h�:Z����!v�C�\�>M��J�h,��nj!_=m�p���(������\خ�[����p�S?�qx��4�}丫6�y�넔7=�W�u�z�Z[��k��۩`�ol��N(���� v�xo��<'�}�z����M��i�I��F�=�~!�f
�W-�lCĵ��'C�?��]�ݓ��|>]��/:��h};�{���.���͸�R�K��G�W0N��&�Dh�[�<y�,VR�g�ν�uB��N`�Y���DG��O-/Zc��F�&C&{>�OB��o]ɫ�������3@�S��隼��*��^V�C�.T���@���	{Q��ue���c4���g�tFN�H���Q̐v��yX_Љ�XE���S�����WZk���"yt�x��6���`-]�Un:YD���	BC��i#��X�9ٟf�H���P��{a�eIw��Sb�e/f5c<�t7���
���0-��;}�7*R̓ժLſ��_ 7 �l�jZ��2���+\*A�C�m2�9�SA[�p��*=�惪�$4�D#O���@w��t�9k��^�12�-B"+h�h��}]����ø�>aR���7��7�����5�f�ND�����mU6��P�b��7��$G�e&� e���}@E��`�1@Ԉ��G�]%��TҼNy^���(���l�]t�`:t���$}ʹ>�LW��I�{f����J�G��N��a���u|5�e/���S����$*��ހ�ɩ���p�oq1�T*+]��rfΖ������Æ�G7[F5��jڎv3]b�`i�땲�m�V\}>#��Ji)8����7P��8�0Gb)����]��W�ğ�2k�̪dy�F��3$����1l|mw�qz�O��2N�s%o^A���D�U�#�;%hv�|jyTQ�O@�u:uj�s�E�=@����'�Xt���{3"��i�{�!��ci9��jE^�UO�mI�(�]���n�G9VD���,U>\{�S����¬r��HR�+��΅�JT��r{3�qA`�����r`P�ϭ�ַc�߮���2�3�M��ٿ��]"t���'���oi|�6�!��^{2հ��?� ����3.�����p�fT�9��I��&�r*�-ラ����k����������ڏ���>X�]����Ґ��e�1"`!�w�+��X��k�����ڗ2�*���-{�7���|�BЭ9!^-  k4$�� RZrõ�,`��t�	�"n;A��فx�!~�`�����򟶈wP΀�`Q�|�˨��pO�m	N�ˀz�z�8�A� �����}b���)�ӱ�]�IF��F0�W�d��VǧŹl��E����}F�ò&�H�hP���%@���H���
��^$��ˌ� ��ʖ�F@�6���,P *j�5��Aǎe�3K��v;��Y]�*��$�[�o��ѕ������$�IU����J<�d�!�O#�%�4S?&����:��1t�l4Td#BhSD���M*(��䮇o��=<6܋jň)���n���h�T.0� !fJ�!��.�!�0�F.ۣ�kn���'�����&�LV�k����l0S��:֮�|bX\	��i֪ǘDq�L9�p�ȯ))|�c�E�ջ ������/�b��3�a��h��)�����I�S�B���^����Xs�,g�k�]��m����7�wT���FўR�*�{m/�k0�lv�.��%���c}�El.��Wݽ]�<M�!�K>b!��k�N��Yve:ܯ#'��l���=���Wܰ��YٱE��t�;���n\۴����d~N28�9%j���k0���c[�]�o�����`�o÷���4&@��Z�s[ly�� ϗ� DT�&��v(���i��iW��5F!惂�~Vb~R�_}�?�ن�=7��̀�Kr���BD�l�����6�yҷ���U�,����4@P0P����k�^ɐ~�O��.mOA�p��%�����:��I��0�<�K��c`�� $�[A37�&�`lٻ6U�Y�6�1���?	4�*�,�Ka����3�A�6���U��ۀ\9�4�B�p�F2���1��F�#~��eT�~B҂��%�/��͏��	��RЂ��,��+�Z��ՔC01�KV��	O��g����Vv���D=���"+�Y��٨&D6��~������|�o�6d<p%;�-�.�8�j/74y�6��Y����c:�GTŭ�RD'd=V[ζ��ջ�䜁�>��u{�qIB8*zd��)�ڰ���7qp�m��6���s˧Uӯ�5[^�����3���\}�F���\�6�Upw+��%�������n��LEBǛo�A:�/����H[��)>F�Qy�L2Ci��`�∙e�ޛ��I�k�P:���� �H)�#����u[�a�x�	W(!*��M��������3�1����qQ8jbl�g*���.�_�0���C W���ug�n+f��n�t��'��P^��+/"xBӪV�rVo�������nÁ�$���<�n�bC����1���?Um�W|�хO\�x�ݼ��Exө�1�osmU��wQe-OB:K&�G�NgXk��8��6QO�jo�iY�����ۭп`O|_��ף���гy�@�����gGÓe7�e�t��{�Pf��>�9����k\�g�z�Xв�v�ս��n��+�_U\��\�����g:���@G�@�� ��XP�`|�ekG�$أ���ç~lf��\��N,^��x�n�Dbb*�j���(E��Ʃ����k��,�^�	�^��!`"��f�|i�b��=@�Q�M�xo�@P`����5�����m��P�@�vCjJ+st,���o�0�jrUt-��:Ig�Z�_u�QԤn��E�d�P ���C$\�,�޵���	���M�Zpڅ_q5�g7ȈU*F���C���Շ1�8D�"qD��`����/L����gH	ؙߣ�>��'�>i���G_�y�[0w��R����'�v!�@�+��5i��lz�|�aeW R	HٌU��Ew�G��k�l;�Ns��V����g3�������>���A��(����U�c�6A@1��h
��2U�Z��3�*�'f'��>s(8��k�������p5O�25�H�������SyD6����
�?�2�ܼuJ�[TH�*qbQ�iC��H$�G�g!+2N��!�E�&7���U��3���Ey���<�,
qS�="���l���X6x}�HGh�w�il��G�6��!C�n;^�Y�M�0�S:l-%:�<�v#)6�}A'K������-F�D\�-�E0��f�	�**�滛���w#)Bێ,�����N@��b�Uuj�?G�h�K��@���-���j'f����[���Ǯ�]��ؠ?���^��z��>)�t��1���5�����:�����	f̩QקV�m!���D������=��'��Y�p������`�.<�+�^M ���.	u���'MǛ�˝W�|�d��n6��AND��*g�R���M\>�I0��ڴ�\�c18
k���ab��+���9�r�|\�Vj�O>�?���Y����q�n}/�-�7��Rx��$�[c(��]����$�hv"�fP:6C03M���5v��vS�3��Bo(:e������l?�'i��Ц]4/�ɯ!`�!� T��
�.
�S<�wt[�6'�_]���[CZU�~�^��$�L�����4����E����M����F2��>�$�lV�\����~�:��y4���Ҿ���ƅ�a�T#�YWp�U�������4/�|��!J�����$fK�ۤ���j����!��O�+���`<R3��5�K5���ѝ�1t1((�L#��0T�u��9� U+�����+��Q9yq�r����Q�>�X"�vSJ�aX�[Ҏ��ǰ�%���[_w�?v,�hm�����䐧kԅǰ��͎:M�r��������W:�X
A�M*ɧW���k)ד��֕۰�kq�4�_;��k�Siz�*�*�]�/\R�n���+�#J�A��=�r�Jff��x���4�#[⏤ٜ��Ň[��~�����Ah���l������	.\�vY!�3]fu)��RQ
fxY���m�<E�k��qj�(�Y����ؗ޲��.���Q��f~
a�I���ù$Mq:�Y����Q�`�悐�mZ�G��� m[��s&�6ՒpJ4�ya���Dj�UG+j�t�`ikvy���Lܽ���\�Dc�v�lFjZ�8�"e��`(G�̦W�N�k\T��cg��x��1���� ɑ���qo�D��������d��wՊG�g�~M^���5�]�$���3�1��
6r�� �-\��@�X��sr&�^���u.$$�C:_����[���-�׏ ��Q]a�S���Ɨ��%]�K9�o����_4٫��{s!~_�0�+>���;�7�y!4͐�P����ʶ�E{��ŵ�
�\��R�as�d��fߏWV^.ݠC��TCY�$8�K������k�2J
��ڑ�I�[�����E������@1��I>҈�U�����Q�Y:�RY:�/?�u�3-��t�>���n
����[�,O�x�)F)�]2 �Ҹ�]�'h[I�'ex�%���D��⡧�_}l��0��I��I��}8f�1�znA�[X�&�eH��O�ȣk��}�[>(�n�\BHc�V�~N��2�?�����-��MGx��[]����+Z���@}��#���0��TS_p�U����"n�ڸ�@��B��K롐�Y��I(��l�响"�N�S:A�v�r;ݫh�I�ّ�k���(#T'���T
����=y)O���gKF����Q��H�F�{?�C���q��o�`�ˏ��=ʆZH���Q���3�j�"�1�����	�*B�~�6��J�B��N�)J�Fvzajk�|p �6�E[�q��LL���6	�����CF���7�V��Fi��{@)��m�7����O�s�I~=����q�ɨ���a�n����;�.j��&�T�'Rn�����>l\*2n���ł�8+��5���
f�<>�`��-'�{c�W�`�"N8�����a�;ż��t]�U"��hT�F�>�d�?*B�(a�#�tm�(6Ie������p��HN�ʇ����!��0w��2&>����W�kK�0M�<�E�Ge<���5迓�Z�m�����SH�d?,��S_1���6��I��R�������s:C6qG����8���M�5p<JYS���(���^jU]s�?/&�+���R��%6e���w��'@[zԢ����N�''z�@���s�^ֆ(k�J���\����K��@-���x�[��G� Lt�E(
�4��lSk��Z��w� �T�S|Wi���o�����QP�&C,&��e�K�.tPi�ӯ��EhG��s9����ԫD�!�v����Vo�K2԰7�5�<��`��v	�'�"�@]��,�n#����!��yr���Hz%��
U���/|о@�ɛS��~���)����0��MU@��L�^t��\MNQ��n�N�����ф�2�݁��G�߀3��oE].���ƿ'S�p m-AR�2S���2EM���*V��4^�=���@��R�c|���Q�	@��[���Xр+<U�a4hQ���2���������(��2��t}����)��VN7y��~�]Z5�{���%���a6V�� JBط�܊	��p�	GM�p��O�E�۱4ݿU*��>chE��N\��!l��&f�ڸ��9���V��U�
�5��<Ϫȭ;���	�|��t�k�	i�o!�����G� TDm��Q/oe�\�ŉ*º���V:J�Ģcj�l�ש6���8�5	$�x�ћ�O�K$)���N#!��&>�X
�g[�qx�U��6z�HJ	�i���Sc8���E�==y�կ7\����=����z�����v#���ͳ�0[�_5�l�>;a����2T�	�-T>v�eQ^�+�,���o�
����^���S[�˓��	! ޷:i�Fj��/{��攢�Ϧy�-N꟝4�{����m�|�¾L`�`���B����aVGp�2�Cqd&z��P�b�$x�칒"pm-]\���H~)M9ݪ��'=�^��%�g�ˠs44y]�m|��+� F)D�>�4�}�X-������y����*ʑo�~�\-�c�˕�QN~�
��u�y.�d[RBz*F8(�=�J�y�l�nשp�V�
o���C�J�۵#���|�S{���My�x�>֠�j%HYO�� ;y�ub�++����W�G�������O`[�?�"^hcč�R �eӕ��#�pSB��J'V�1͑��ZR��Y��aW���0W�9��T,�9D�MbR
�W���7�7}��$����j�_���")���`#� Xlp��{|mvb5�k3f
B��w�y�ָc��PWطN��D�á�Y��j	b���x�Z����c!Gly��H��tꊹ(}(8Y��e�6V2=}�@�����j���f�G�?����f�!���ズ��O�J��<�^�I�7x+�n��G
��h�e��O�ؙ������EZ���Rs��U�+�[];C<-w��5��,�^,o�TjXY'�g\�~)a��_�t�HC[w!�[�xע8�/b���&���IH��y�`��.���Xq��y�����⾞�*ׄ���ޑ�7������x�Ƹ0�������6_�\��ɢM�%��|M�Z���޾:�p/���S�{,�9�"��XV.8q���۝_�'�5[��GSX�l����Vȇ
Eċ���d�s��4�	���j�q<eX4�T�M��'��4D�> í�`C&(F��a�9f����t�V:R�Y}g�c�?ҡP�}��=�"�e����f�8Y����#�E�x�u�+��7�ߠ�v"*4/�9,�1B�1vCmV�h�� ���4�KpE�M#MX����$�<�AB�V�Q���4z��m7�ׇ\���ݘ�?a쎚6�y�u�^n9���ܖe�R�!������禣����\y�*C��h��D=3������(g&4_e��Ğ�������\[���m#��N�~��h��#� o�a���,��K�6G�l=hs����G�_�'f�^ӣ��U��GY>3�IJ�+u�x���:ހ:H\_&�s���u*YU�*gE7��/���`]j�2pn��8CH1e�-� a@܀a��d��V�?�f
nC4
}�hZ�a�]'�����H�V)K]\
`�������W�Y�ݥ����q#4yr'D���Ϭ�~$TGv�J�ӷ�S�U�JQ�f�I_�v�nqԿ��NLQ1Q�o�<Xἀ�i��3o���٥n;t�LW!��+��([rq�\���p�_�$�!�X�<�V�����oğO1W���4~:'�ӥ��!{(��#r^1����0�����jaz��:V��(&�R �X�	������]h3�MTp]c�O�c��D�Ʈbm��d��
z�-@S����e"��A�co�|� �y(I�y�2-�ΊB
�"n��5��c����&���
m�-�j2A�ʘ��o��w�<X�z6�,
�=at��48Ta*�΂qdb!Z�[i�[o��vw .Ʊ����I�����Z?}�ڵB��ל>J&������� ֮g�5��a�'*�v^��n�(ؖ@	��Au&� ����21���U-OĀ.�S����D
�n���=sv��Ħ�< ����l�1��V��bsbJ央���b�[4,Si\���(���$�������8�(e��W��q��f��D"�]n�y���yzS�_¾�Y��1��/��k��_Ke�+�
�l}X��Ճ�Ía����K.)�(������qZsI��h6���"���u�nͱ�+��.�%��$f?����WP�J���K'�n�~��"m}�P������k�m^)ǵBX�jjY�DF�߲��B�MM�K�?@�虓���|���[��N~v���'�
ܚ ?�LD����@z��׻�S��=�A[a��X�\����v-�/�IP�>;�U��86�	���w� �Rg���������޷���>N?�D�*�&e3HLc&�=%�����"K����D�9Nj��U��ܮ0~z��T���W�Db@�_���e}0��t�
�Ʋ�7:�Ѣ�
r��fE7��ˢôOI��<z�,z�b��>��r�F���v�#��B����wi�Z#af�/�����f̝���MF��"\��3�� q��jmZ�ƴ��v�gN�S��;oR��@���y�����9[kBZF�^P��T�,�^_���g���(N龰�bo��[i�55pډg�ǵ����t8�&"�mc|r[1�������&�u3M�#�C�*�@�j��s�&JF{��P|�$^��̕�3约�!�U\FH��	��z��b�=��нG������:���>���Em�.=�I���
�'9T�ܬv�-.#��u�
��3@!����Yta��ԅ�W,����<.�2'D���R �&־�.`ur�7�����<i�b��O󭟓F��es�5�;�����C�sN~�;��5��y�x��Iq��Krʹ��8�����m��i���y2���}s����"�9}~�j��~��$ٱ��M|;��+�;���9E����1p�a�|�SR�_
��x2 <����lR���S��*I4��<����g�����4�e����T�2���T���0����?7�����%�{�O��;�ˈ��w�������/'�ǮV�A%'�o�_&7\��HŒ���9Jwei�E/�gT�����W��uf�v���~@<��fS�u�[Ήj�����b��f��$��9:M#+:���z����� ����g��$O����xTcj������4�%ia����x���ڼ�ha�:$�/�f[��л���V�C��z`�7O2�'�AJ�L��7R��{b�q���O�|*u1��1V�_r�Ef�����7�s��^&v���L�?,J�������ިh�/��o��d��]�O<����_'(��Gd�4>�<����P&?���4Yq88 �JY/�>���r*0�e�2�30� �TM����z���ߓ����#��l���A�&��A_ �f�z��:s ꥟D��)���D���DHP~��w�S�?����T�A���-#��H�)�Q1�"��]��]m�5{�L����)����ڰ�Gp�?�|;��N`N����Ԟc�L��6xI��f�4e�k8�y�����z�,��I�qX�-v��m�o=�@�b�c�)
�y��̖�c���4��r�1'-�EǞ��G�!5^n�%>�;��L/�� �&ٳG�f��!���o{KP�d��Q�Xrٲ}�C�9��-�"�SS����%�h��i"�:?7���;�?�B5�^D��*����_��74�^!Pʖ'�m��-"�s����}��3H-�g�	�����u`�} b����
�q�AIfCn);k"K^&ޖ�|�S�����J軔�
��]�K�d��x����L��~U��2�>{���~���2��7���>ƝWv�>��*�0�ʝ/�7.b�f���&��]�p��U.�Wg���c�̎K�ZY�)�+Ժ-9��3��.�������-̱k�ㄩ�A�������gca)��I6![K(��Z����?��K�t���8}/��"�~�z?T�	�;���s�� ��Z���|��ŲUڊ}�H�	C���� ��ɴ��rՖHeQb�y���o��p���I�זfov���݌����l�����[����"�� >��f-��j����{�-� �d��q�B�n�D;��l�ߨ�
:�~��!�����ƹj�wW�Jm</�h���M Sr�3�sߗ�L�����8�n'm��J�����'_��v��,����Z���&>c�L�6�Vǋ~91� ,޿:�)����v�)u����|p�0�<�&���:?"-�Hq@y��y����2M�P������JJ�M֟�9~��;xꑔS���[���zd�(oO������������1������D�$���TT7���K��[m�5����Y/wP^sw�Wlj�)X2�Bj�����w���z;h���q�%�3í��k�-Ћg�ƂΤ?��=*F'Z��i�q�]̾�t�GM�8ēD�7��a�_5��a�Ϩ��	`_�K'�dE{rj5C�kjwC�Ԩku���M���� N	��};d�Lw�:=݅���.�gJ����Vd���NoM�>��+K)[K��]�6LS�V6�fD�z���b��q�x�����E�,��t�f��3[��^}�&
ޜ>o�����U�9dl�O����W-`C�(��]�i�"��N[x.e�d_tb�i��;e�լCTM�gK���4�3u�n!- ;%��w�`�O��s��#k�0d+?m�7�IeU�f�2�B�j�%��+�
r�ƚX�K��렄�;N}И0V`�$�D;�䜕-9�r�aٳ��z,Y�q&H#(~D����OFXx˄��+���,�b�ЗTr�.���������A�S�(ѝ+p$0y�7}�Q�t�,b7��fwsIg�t�u�ݢ���X��.D	L���(E��O���yq2ȇl�>�x�uE��`����g�O�ؚk+�eHvkZ�����>�6CYڅ���ܙ��=����h�!�����m��9ы��_�D��gk�n\�3J�s{{HH�n��[�_��;����q7ə����av�c���b��]X����_9��0�lX�(R�X�Q��Vi�k�KG��edRW[������h��"7��KC�D����|��g
�����%Er*��2T6ɥ��vşd�1^!��"@�:���.���V�U���o�?��f�z�}��x��N��Rddw&��t�����{���Z?���!�#G�_�z���"�9�c�$|Y�cR��MP�d-9�x��j�EFQ�� ��L1��o������J=�hH�Q֙�B�#��_�-#�7��	���u��9�%�ϥ��u��0�v��!��g, ����pI��H#��(y�u*���_��eT�rN[��.a��H5��h[�L�B�Kf�u����-��?��!�U�s�.���e�_�zR� L�8�FNHJý�k�J�>��Pgr(�A6KXވk'�S�)G���P��P�Z��t��j sj�hzU��y�l��3��'JJ�m��=܉���k�:>�A��K#e�ԒJf�i��h��<���<�h?�l,�T�8�	6�m��&W�	F>�,Z�m���Y
R�$�6N�x+�h�Rd�#ςɤ�Q�{�§&-��%yfdc�v8#�	 '�s)}�XrC"��ڪ�����y����@O����4�E�ҍ@��>��c��F!IQ�b�t�x�ó/��s_*��믑%�[�E�Q T��c>�6U�}��]+ș	��qtv{�(�Kd��
��L�`����8�}���-#�`fzX/��Gî��Ka�fk�LZ:h��o��t�v��|��y+�x���#%iW$5"�3-��JN��m�d��=-��kH��u�̯�[q�)��p)��˓(]&�hh7�~�ps���k��S��0ʺ$�^��p��tR1l�{ ߝ������m��m?C���"��Ϛqk]�����Ƅԏ�7Ii輝��o���S�!�D��v��pF����b�=�n�M�{󕸗YL�1ͧ�=�1Ϝ�@(��r��V��ڀ��Y���;��X&/)�m9��t�D E�Wq��@��r�����R��V���	�UH���������)6*�Cw��i��4�����U���{�����3��`�XnM�ū��v�q�l��d�����)O�f����{�2�rV�Kk}�����{Y;��x�oo�ڗ3Z�N�pU
�ߊ�,�,1�E����/#�V5�X嫕��	���o�3��k1_��<)��5������mD'��Q����T��v�t����B|�d��M	:������Ŕ��N��_��ֵ���#J.C�����H.�����Wg!'���C�ޒ����Y�Tn$�!�X"	������x<�q$d�IR`]J؂�C��D0|{�[i�v�>l�jG��$����$���E<���$�sP`�?Sv>�n��9`q�/+U&_�������0
�?��'":R0��/�%kېt��