��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T幌�%(�j(�ShJk�0���Nz��)S�1_ܻo�^]+��蚉��V��;i3ۛs��Ͻ�|��5�Y�&���%��.��ju4��oY"BR���\�N:�7�e�^]0����s94*����|�>~B�n�U���~^`_��������ZT�{��6��O����5XI{q���]�y���2.�����ך�
,I�����[A�F�rn�	BA��;��T���J>;p-��=.�ȼK�T�_�T+v�H���d�f�>�6�f�����B�Cځ� ]���c�p!�)��3����C��s�����Ţ%�0�qƻk�]�� ���4�J�{����EI4/9i��Y�e�c��2s2V����?�x�a+
:������o͕RK�m�=b5���Cs.�F��뵮ciy���~��L�O5o��@�y��+4�>?Nچv	^7ltP����|a�L�Z��^��������P;K���ʋ�}�0�-��*"=��J%���������ZD ��/9�����q>�����s�'<��G=���/�!H(A�9������I�z6<�[a����������e$��Zz�L� �a�1:����xS��ા�Ñ��1%��ض���ٮ����eĔ+S�y����{
�2��r}}!�O���4����v��m{�h��2[�c��ʍĥq��Ǚ�8ޟ�S�w�Z�8����Gp���������߿������n��<rD�,TX���yڋ`�@���ޮBv�>�^:-��Ƨ��E��l������@_�I�0�K��$��y����#��9���X��
���ͅ 6��)#ڥ:�����m��,���C;���B\3`�N���8�dƈ,|�	b+Ը�eo���]Tf�U�X	� ��:yѵ�^����J�_���b�-����dV@�9�o��a��P�����rIf�"P��,�d#��]�n��r=,��/�� �3�	Le�-:4�*z��߱�a��޴���<�h�e�Lo�\�e��V��;�+[��
�69;|8a�H���mJ�_I�`9�k{|a�T�~���Qv����Uc���"�$�����mfL�G���"�W��f�Q�[V�qA�؟�1�+��Grrb\y�^���[�����F`�,}��9k��+���n�2�T{޲̄����Tܙ�����v*�i!\iwrR�}�F�r��M�h�X�i�j YI2��-���>0��ּ�$l��N.�P�Vyfq��o�G�c��A���.LR������Rx�r���?�{�^��u�|
4��c��L��^��g0���J2�>���T���������0a{�����!�q�ۻ<nܜ@�5�6͹
Oi��kBW�4�8kӎ"sN��6x��z=Z��T�k0z"k �)'G8�#tsA8[�3��WfE�&"1�v���tݮ��Y6̌�Dh��B���?�&���;G"�7i�.h�w΁��O�hp�{�N�룇nZ�#GU�M�f��o�+�X�~��}&�,�6bScx5Q��L"=v{G�����F�QM2�QZְ�K�4�'��+X�^�}�(j�Ӳ�S�MWK��� o;8�A���j��ʖ��J��6m���Z����\כ�]f�}!���Ϝ�1� I�L���%�a'ͅ�X)	��*!DnT�":�H��.�	���m��PS�W����j���r�V&��׶� �(�B�
��}���ДL��ӊu�-K�Ц��!��nV���J����)[�D�)�rG�_'���pfp�2�#7.�py9�%]�� ڝe�p|�GqO<���T�%kt��"�GV�لcD�jQ�ߟy���y�r�������֪��c��}z�� ����q��Œ_�Z�.}��SB V�"��Cz~R�Ȍ,�ߕ�U�b�$$f�,�^��H������&*xq>����W:9�_�->�\���㍍�B/�4���2��#���Ea�|�G�:��?�ڽί��H�]d=�2����Sj�|�8����,��� �+�V�W Z�	�0���4�}<�6���	��n�v;�m�2����4�����M�f�������-�̱=���Z�<d��"h�9 1N������ci�FGK,�cX�|'0�t1D�����'��J��
$�a񾋝��)J��PW�3�h�!t^2�QK4��Y��Xg�k�#|��.o��^_�$��z�����fY��Յ7�� ���c��,\.����|m���b؝�Y*6��-��W
�@*|��&�L� 06dP�N��#~�0�"���To�
�O6 �B[nِ/P�FI7 �n��bR/��B(���E���R0<�t�����tKG��ݸ��z�L(͞��0<��i6P�%H�����ӅȺ�0*}�欟ә���Q��F�6	މfmr~���D~��2�&7V���W�j�r�M�����XgT��ܚ3B�����G)��*�fo/��٢71Z�7���{n�(�C��pgB��P >�g�4m� (�Q�R�:�f�����Z�jz�w6�C����)��]���K3�-�`A�)�h�];����;A+���s���x��?�{|��e�0��H��c�2����1�q��Y�# 
|�(&&o�JRhe*�V���9t��I�V6 #��PJ�j��1"x+%@��n�C�}s��� N�Ob����Cg����Q�s8Z������\��Z\'��
Q�r<�"���r�B���x�w	�,ap�~��� ��%�V�2{, �D��T��{-OFI��~�Jֺ�F*^l`!!}�^��Y�.���Ȟ%��K/�0�zz�GT&;t��jO$)є���[�4��\g�q�����G���E_����9�[�04o�����i{w?���ʌ��4+D�Q�#�ߠ/�^�b
@���?��*Q�3�6�0d͗�#_S(!����Z�������k2td��NH�f,yl��������c��E?��=�Ln���{�T�G�7�4���.C�PĲwp��?ST�Sڟ�x
��-������S-;,~����=�3kmP��zV�����~WC�6�-~g�'�E�喡��Pd}Q��uÎ����ڼ����U�{?~�Jr�W����BKq˯f�G�i�
;���Cxpt���xxH��<:�Ұ��Y*j�@єW@��-�j/ۍ��
�f��4S��+�S<��T�3��T<��%V�b�+����fy�����*+�}��>��S�86���@�S�~}�n?�lP:(P���{���D��Dl����	�E�����i�n*棿�V���e��t�0�vK��}�6�d�bx�Kx�� 3j�v��1�dP��"Y,����ey�n'ď�����`��8jbev���@QfK[������p���d��,����~p�,`z���Е�W��h3�= ��a:�ɹ�,e�?�w8(~���O�e��D�^�����Z;�mB��AB�7MH7r]�X7�n���8�Z-��sK��Qk�bɭ��t3O�|��9H�?��7�v�R���7��iU�ծ�J�N��6���P�Q*~ϡ]�k��WD�,��svN0��;Y�8�����=.-�{���� �S��Ƶɋ�3��&�'؟!$_��F]�%���E2��>�����:]҈]���GBǎ�xJ l_���8B9��la� 3�ZG�8�N��oVe���!�/�n�X���ȝ4�5_}�Ӻ�����7�~⽸B*W�迉q*��Ds�mvE 7�A�l#���Vo7� b�k*])O��3�َ�K܆�<T�+Z1�i���N2=���\6:�,�k+iR^�IL6��7[��w�Dv#Ɋ��k��������ci�����Ĥ�]�!>q�Y���*�x��v���-��	��q��&�	��54`�UA�t�}2�����X�UjgC�	ӯ�#_�b�)&�Q���Y؋D��r�M��.�(J.J~V�@�9��5�7m��
b��ѡ��>~o�f|6�3�_��$"ع����Zd�w����H�ۜa���x��|�'O�T-wGw3��K��7@����7�A�`����C>�
��o�R�_�ٟ��������r���+� ���?�����yUr��u٤��y���G+��Ek��	�G�QQQP�{�V<	1'�1�R�KFkxcYi���T]Է]rK5_�}�؆���|�m�SѡiK8F}}��I�Hq�@J������_��z��S���_�t��A��h �A���3Ɓ�c�����\g8L�.j��L9K"��~-�2zw�:Q��Y�(lզ�>!��=�}GQ/��i���k�e������1K�h�s�b� >��Y��B�U�LK' )�t ��7x	
U�����E*��
lP�pxjUƞF�˭ϯ�������C���wv>�O��2p{���ıM2Lh���*;�v2��ï��6�5�t)Tb�{�紶���#��CQ)����h0[��	�e��[DH�U�)󰚉lu@!�#G��@�&��m)B.Ȫ��	\������n$d��e��?"��h�φ���4EǬƴS.�){�m"���l�`�SF	�=��0n
d�s����01�0$`\�B�|�P���B8W���/&�|�w�j�T�?�"Q� ���8�D�A
�Ks>�*��������+�tro|����%	�+:�R����nz{�͵k&�=�;�O�C��jdh"I���TW��w�g�X�o˩2l"��jR�aù΃>���+ΰ:�Q8�/��kq��Ǘ��4�����X{�`M#ς��g5�2�Nv�y�Q7�Ėڧ�;eb�*��U���v!�	,�2��M/0�w�j10G��vv��[5J*�dK�f)��jb3!Mah\W
&��7ծI��Hl�wQ��r�� �h|W47�m����T6Xw��)}�y��B�E�.��N���%���������#�^Y4��K�5m�,X�/��S�`'Ѱ�p�6/��Bӕ��b�����TXM�քoU)��\����H3�0m�ظ�X���=��?1&�,�l옟��w��#ae�6���'C�4��}��Y�5��ٔI�7��d���8�iӄ�IO1ci��-���(ajmm���+�_����IC�EEJ�q�l�����o@"G\�!ن�7p�Q�L��}�)��l6zb}����J��f��M�\9��!��R�����������éƈ�+G���B�,��Iofn#픃���o	�c�c��W����E0��%�CU��ܫ���|9�0^[�ID�	�Q��Ʈ�
�ٝ��]��'Q�%�LT�~[f-D��ANİ�-{?�� ����\�{�������K��zx��HY�oޣ�Z{��O����g)ަ?���EfS(E�/��qJW���F�h�(������CMA��5D/��3�5��&2n�X���r�J�f�H�Z�j�p���r��>�����6ʑ��p���Νc�Zƥ�R�Y��MG�Q�_�uA�\�`��m�n�ؘȌ���%Zh+¼y99,��@Z�O^r���Z���Q�5�˼.�n�_J�N}���-1$a�n�f���529E�~�Q���j1�eD�Ѣ�Wh�44�J�ٜa����i]�絪�����x(�4 �x���4�$8�M.���Jk�%�i1L���`8�D4!��/�w`�E���;���k˴~���?��S�)+��̳T� ɃR�B��,>A��X/���y������wz���L��I3�ߥ*!Ӿ����ǒ)�݈�9���pCٞ j%q��!9����_8��^��X�w�i��+��$B�vrY�a��;$A+����1�3y�=��_�ifn��u.���Y��t���!n�M��kx ��H?��챬��4d���+A�}G��t�ۗ{�GѤא}��E���8]H���y��Y� a�6P�����G����xY��
��Ϋ��ؚ�ds�h�sb�l�#��d-�G�	q.�5ۋs����5L�rK����m�ܭ�U�m�M��t�Oۙ�`K�q%ZPJGM��������h�61<x���'��7ʔ�Q�=	LO�I)����I��P̋CoV/�3�w;���S����<Î��Win �k�0)g��!���^�{wSl!c��ư������WC ���3����%>ilnN��r�aY�������ː=7��\\�v4n9�����\*�sd� �,<��.��S4���hf��5��r�,b����L�8�akg%��`d�#[�����*qfG*�^'5�՘���$=��b��ԁ_��#}y�R��t,#$�gD��u ���.zw6�(�ᦉ�٪���9g�۽�����T�W���X��g��R$��L�<r� ��0ѩ���(���AF��)F��͜��{m�ۘ�k��W�p�S�ÚAf �l�_������+d���f��r��6�s��H˔猅N�_{�Ny��%Y6�C)���X�TB�sA3~T�RA0�� ����8g��~�nE����ě����	�Qu�q��Հ����.]�BiC9��-5�W�f��@���\���)T�;0�c�+�0>�&|� :+y(��O�%.�4E��h�G5V�*��˅�W]�Z�Dx��f�.����"�������:��ZG�Xp=�.G�1��f0��p�;�:���tV��[��M,�F[:A��㸌t9���������uӇ`5k<A�wgXL�&�	\=����/�;�2<i�����1Qg�j�Wz�|����"!��(�5��L��~a�J���Q�1&�]�H���c�AW9�f
���%�G9��:R�S�kw���܈���s����'e�E%��p�'j�>xݍ�BZ σ��|zz�����ΨI��w�Z�1`J����QE0��a����C%���9���&�d�avZ��7�#0ڱT��K�@��b\K4����e���
���;��{dQ2T�C��9.��BX��R=��1�v�!�U��4���4ׄ�ך��^�%��A@��a6{I�b�)<_J����d~�@�X?�'8�0Vִ,�	��c�&s7h9�#+��Z����5���g	���)�.�k]f�As�Y8�̈(�[����1�A��erh�2vF	�V�Z�;O�|�G�fn�e��_J^!B�:�ߐ�5|&�Sg��;�������ʨ�ȹu]�fھ�"'��s��J��0aL�Orz,aU��ʒ��1�a�3�ظCh������R$�[1�,Ǣ�f&<����I0t{�;G�fY���^n/�Ty��\>u�o�`d��V!]fm\�g� uӪ��`]���r�6�Ҳ�^�{�s����&���G~���:��y~@3��ْc�^�R1������ٽ��_���FJ�$�5xz�˲٦��6X˥�xޢ�0�������5H�%w�M��>�U�w��2���Fː q�� -��O,��P ��d�����2k��"�mۊ6���Oz�N�^b�m��%�v���ķk����c���>���H_�·bn��RN������e�w�.k-�]�Sd�an324�Y7�z��w����A�\���j��s!��_"hM2��J����;���Q��h�l�@�Y�/�~\��@��-��g����P�b�M���M�*�vP5��ȶ}qX-�6������:���f~­��3�������x_��>�m���C���[ěbu1�b�ض�F��f��LxHB{�PZa����;�%�:�q	�F�{dp���I�)����A7�i�of�eә����W���3�{AU��]ti�������BE�)�����u�7r�˔<�޶��Q�K�x�؟�ёe�XA��60ǫ�@:۴x�媒'��	���؞�LD�T&�-���ᘧ���3�k;G���;n�oNZdLi���fQٷ:�������y`*Q���������w��O	ρ����e�.��J��ޜo�Sҁa$hr�h�8dhB��Q�	8'P�؝��J�d �~R��-�J��+YF��A�eN��x�/��gT�Xb��5�k�����]n�5�t�dvJ2�k�Nֺ����БDG���yD�Atx���sy�б��]����+�X����ͣ�j	P��
JMA ��0�?y ��1�Re���*���<\NY�T)��<�o���ǈ�hU�UKQ4_|�� Q�e���e �P/�������>#�֙���V�v�Z\1���i��i�B���
�����Pe%���9�0��&b�E5���r1$�Ъ��EO	��jmV��=��%��.M���dA��f��ߧ#��<n�xoP��AKO}��\H�`�����_E����w)�GA�`+� fs����G#�[6��?�`��)�-�3�J��\20�͊K}W�QZ�j���!|3}��<�)c'��p����/m�B�%F=lb�h����K�
�����*U3�C���;k0+ނ���B����>�h�;�}Y|���ˠ��;+{G'�uS�Q8�'Ο*���ނ�揹{
���p�Θ��,2�"���;�U۽��+k��?0WY�Y�/!�Dإ7D���ⶍ�U꥖�+7�m�b:�A�Q��B[�\�	������K�@��k�
��kWd�̎3D�X��]<ͻ2�xDED ���/�Bc�rT&M:��^��1Ѿ���d�r'80����b��B#�>���1�׍x���Q�h��$0	�y\�.7��x��H��'�1�d��_���O�"Q8���6s�j��e:>9;O�/s%��r3&�{ +���4դ������i�]��\�'d�Y�� �{����Y��7�I�p��0edC�1\��ƌ�|����b�W��d����5q-[)�Qu��r��>�`��(��G����H���LS[������� �R�+�9	�<�$!*�3*��A�s�m ���m���6�����Ro�>����7��l�Ջ-��uM� �z��<c~g�dS*SeAfq�Տ�����1�/o�8��+^sʕ5W��;�����{M͌��˙&�8������)�؛�����ڨ� /|^��\i~���� hOk�C;9�"L	ۈ�-�p���S~�ۙ�mI��6�g���,�p�$�H�Ѧs�0�J����H7Ր������6�X4�)}�ĳ:]�������ʗ+�zV!�C���2uf�>��NI�3�cT֍H��ji��?\�q��K"�OP�F�P0plI �D0_u`պ=��g@�q݂���0%1��%RA�5̖<NR��d B������{TJľ����m2\�Ĭ�n𫻜�^��H�b�:��2�H�7��F��p��Cbhq��^o��3*���ڇM�Z����쁎��e�6�z�;}��w�2�'�ޅ� �t�!���Y���:��/� ����t
�zj��j�Ӆ�����ˠ�V��[U�/�%:z5�y_	�T4X�V;�.6����_ ȂEbc�M}D!w/E
�S@������8$�ݢ���?2��I����SFv��j��My.�p�����R2��E|V��nQuu`W!¥�L�u�ǂ��ˢW�����{u�����M�� ��e6wO0���a��J�W?0��ܣv��vZ�)NW*P��cj:��p.n+:��zSS���S�f�0��3�5����;�,N�;+2ǃM("�P�:����9����y7���B~\lg�Wh�^�1A=�p�v��fIq���n@�R~�Ո��u��@�#������=�dJ�!l����=r3}C7S��Qh/[������w��}�
2��=�	T|��M���uf���Xu�y �H�������=&�[�DSy�Y!���
��ao�����@Z�nf3�gLv�џ�>z��+6�|\���'�Q��&�e�4�/�o�qa7�^/c\��N*n�k��e���g �����̮TG��LX/P�Oh�"9Z�+=g�$�� ��*�w��P��?D�T���U��Q>��W#�F*�߇<�x��z-DP�}6��ԒX}db7IT{;�A4[ʸ�v�癌9�zK��U%#*`j�Q�Ya��5���7,3+\:/�Vx]H�wx�~�U�X��J���ė˶*�S�N�����F�HQ�[׿w{�Қ�s`R�#��9a���n!��1*�Y�Λ8IT,� ��X�ʧ��*��S��@���<��8_v�I�����s���Z�a�p0�e��tJ�i�^�ʫ����w�}g.�D;4o�-u5�V_����[�����Ű�NˇD"J�#��,���^x&E���W�{�x��G��k~��2�<��>��awG:f\vE
�|ǦD���%耶y�\BO	��?{���3'�}��s\n%�Ƌ�R���1i}JC�o��E�dZtJ���T;ų؟ɒi-sA�� V�S��2S![��d�7_�qV0Hͦ��βҖ�~����V����%�[�cC�D�&��fKP������w�KQ�3����du�f~�H3,H�U��Fc�,���4�2Z����RZp/?�;�> 2�W��𐱪�t���!HR����G9}�Xΐ%%��
�
�9E���uY���1E{Q�M���,�AŜ"�X憹�4d���iO?�[�lĽx���q-�����q0� 1w���X��G��z��]M1�ޒ�RO��� ȣ���z�{��H \_� �9�1�Kru��myj~�31Ւ;�4iG-��?��BuW%��F��͆'Uy�y;���T}MD`���'p��B%����K����_���<�n��C���S^Ùu6���[��-�;գ�*Q���WA��}	gia��U�������t�6�Š6����dV"�����_���x~:/h:�͋@k�	%7�r5w����Q����u#��NbPâ����I�(e	T{�SM�R���5���קb�1|۲8�`J���m!�yz�J!=��Z��u�e;��O>÷��.�'��3i5x�g*W��lp�Ў�A��`��Jou����F��L�Q��[���[�E~���X�H�
7�����TN�&�}�'�R�pS]3��^`Z
�H]�0h	����p2��������z�%A�}=�!x�Y�4 4u��G�SG���:q�M�z��s�|D����IPX2�/�H�u�?9 ��Q�V�x)��j�M�[.N��}��F7M�Չ�K��䊶�+hn.�2&�e�;e�`떛̶������>U0/k��
�)�7�S����4�܌%�.�-��G9�JF\�M�K��� �1 v��Q���P^�7t�1���
���Y�9v)i�	�_S^'��M�%���Ku�вx�S)�P����5+�)�R%��iݴ�{�z�"9���qm��w�"����-�Pr��U�v[VW|tGu�߸q=�Gі�^9��8z�ˆ���k������!^p���$qZDf?DB��/q��o	*�D��*�C�?\
D����Ƨ�\o��y�CӃN�k�mu�#K�H�#ʔ�$���s�Ʋ9���!�%�uD��/suű�FmNa������+n���{1�XQ���J	r����Z�d��eZFp]��d?z����c�NRY�I��b��JU0ߐ��+�< �o��l�����ۼP����Z��iԺ^�ʄ�?��'�X6v%���r��J�CӃ���o#
?����f���5 �A��2d	�wТ_��qE�b�=}���\zWbO��o�׈f>�\�|���V�_C���٠�0�+�Z�k��k�{t*���(o�,Zꍿ�T�E�{��� �y�:Ӈ�9�ۍϽ���Pf�j	.c�q[|]�'�~�Oډ≱�z�d�j��gN_zY7��!�/����t-jU1�aYt�갷���?�<����A��� �p�Ȏ#_�b��nّDnA���_�P�$�p5�HY�ș�/�{?�˝�:!�B�|-L�(�BO��\����}�:B�厠B,`�U�P\�� �~��.�'�� -���������]�"`�=�"N�؎u�\~��b�,BA�X�0�nƖ�c�zg��c������R��� �������7d����D[Ɏ�e�=�������aq$��3��������~�dL��b��р/��X�w9��/��{�[f�z�l�U�V�8o�'�!�7�����o��_4>������~���
�����>|1l������fe��#%��H��Xu�u��@�#KX'��aQV�"#�W���+��W�:�:w��T_¬��'���G�������l��E���=�rw��&�Y"��Zju�:�d���5�[0�l.��];!CǙIwg�ԥu�;�[f��0I�̒>6�7��P^|�z�Χ_ /N�Fp3�a�+���$�c��ڝ���$��v�D�jgI\�b�h��a+I~cs] ��þ���Ӕ�W�3��
+:�Z�ف�#�Y�\�v�[g��/8��s:rlc��L:���i[0����`K&�>ǩ:K��ۨCh*��}�(���>�Ӧ]<*�Q�A�V���^��|g7�0����Q�x�51
&���m��^�b����E��^�)FY���z��C�B����#�� ҄����o�H+J��)$��*F��b�|�8��*�S�����{����5qt|+�Y!"NNPFn���eX��eXt,X�Yk����V�ߕZ���ж�i������:� -��c��͵�H�Q�(�&����T��J������э���"��4;��a}n��1L��w`����F/��V=�g��q�bs� *����8�_�&�ׇw�K��{ٳ,���9��s)�������~�{�6
'p_�&���O\i��'E��VY<�Kh���ȸX������]S�ָ�;�)��Wy����A���=���+U�}��t���}�]����:�@�i��oZpD
H|1�XXr�?w=?ZH��n�(�Σ�bhk��A��R�va��A�:?����.��k�K��QT�?Wi (S3����ȇ���d@�)�����Wr�n�2�m�c�u� 1���Q�}F����cKJ{WM�ܡ�bi/x.`�+���1����*t�㘤3���Kx���c��[3?ֲ�{���.��QC�J|�o2a�7��k��"�n�ZR���9�ܸk��N���a��/�v9#�آ��w�����= ���3'��`���aL�7=��n=G�`R�A[P�=Y��6P-/h�+-߳���cx�Ņ��{��d�/�B�[�9\�5�"��f������-�tm�w�M��!H:cO�j"Zx5c�UJ����\�V�Z�u�@�F�<g�	?�s�w���q���$���Gk���M��͐9@�o:��f����{���%�|�� �ߎz��y���I5'/��
�js�b7�t�Ct����g^ ��:=7h���!bc�;Z��o�����OU�~�]�i��6u��uH�]RU���7������v���Կ��R�O����k$�;�'��6��`�\f{��ͷ`���|�Y��qq���v
���Uq;��v����n&��]����S�����Th+�y�7�#iW��Aa�J��S--v��\���}W��@9[k��`\�5k�:�~ q*i�[�d
b�����^N������>�?.,�#����h�<8Zs��9u[�cZj0�t@�4�iF�wzM7I�ݣ4���� ��X�9K{�������E��J��8��f(��S�z6䄧"�0��L�h�!����tWG��\p���j�ӫ���P/ȯ��zN�u����r�)��_b�X������j���at�i�	����
�c�ϔ��͟��'������a��F^�U�3؄*6�+��R}�d��v�+��P�Z?�4�u$��T�!��n)+����6]�_ +�	��6��@��;Jp�1e?IƷUM��E{)�{+ӵJh��([�c��F�RL��[����q���#g�3C�3�X%1�ʔq�n��ho�:4��1`1�l���.�
n�?��@d_����{�$�����yƹ� =�i�|~S
�W�Hd��0���gs���q�y����/� �t����@��	�Jw52�o�"xVH�����1�8�����Z@�'���c\�-jZ�[1�`(��i@L.b览Q���H���,f`�עŌHSC���������m΀A�uKԐ�K���9鮘��A��~�zHX$�i����<�����@�fk� ���[�
z|W����#��i���j��q���*f���7�K�G� �J_�27@�1«	�!���«�Y���F�k#�N�@���U�Hҽb���9� I��U��Wh�u7Ɲ5l�xS���نoK�nf��l�WVSj2��+�OZa�eD9eHY8|.�k��*���5S<{��T/�h�?WYnmR���ex��HH�P��t=�ȹռ�?��/V�7mi��:���p4&i��}��j��Sz�mp�+��U�=g���-�
Q��Aڬ�G���<�C��q��"����{u�|�(�:��?��n�������LH���waԑ1r��ƶ�\��O�3
�_3D0� �o����a*�ٿz2a����M�Z��_��L��_�$�A��f#��N E��?Ju3ҍ�'_�Q*<�X�DD�͎��/��$	��Uǩ�_�(��s��xPT��G������=W@���ĭq��49L�?	O��}��7٠�������W�%E2��;�oW �K���N]箚̸�A���K��#�6�6I9#���)��O��W�8�
����f�d���c]�/jJe��dˍĈ��+�K+�R1�h����h�S�������"d�{Õ���6V���av����ȏ��}7gK����)Cg4s|��4S�Q�T{�h�G����hFL�DIƄgQ���$�A��:����pCm�Z�@�"�����pL���B�kd��jl�|��Qn[��bA�y���rfN����������� ʀz5K\R��ь��ܴ�o㣢�b�I4�
�����LI��@0#� ��%6A�j�[����d3�QM ��V=J�m��/��D˞��syƉ[^��Y�v* �q���*��V��q�����J��v���#���:��r�f\�M��`:��+�_�*��A�ߧ�]�P�۫:xE8M���8�v�a�f����=a�n˓��	�����DD�"��6�� kgņ���Tζ��w�"s5��S�
 ���� Z^}��#�gM�d�^�JS�' F#d��9�Gx��U�3<]�X�+0ݍh��)A�$s!�}�~B�F�g'�s=�ou,,$���Nc|�T�HgQ�2�L��A��܌Ȱ]ͳ,
v#p"��*���M6pv�z<�$�o+���^9�0�X�bl(L��iG���n��`����N�����_�A`�)dfn	��;���.�"oV����<?��>�$���mM�2(r !��ЍPlo7�|�4g�;���kB"����L��p�+���d ��IX�瓹�����8�1���O4�c��I�L����֯���&�e�(É:INmi$.��7���A�!��8��dxR��n&�Q�H���d9����+a	� �����hz6����Uo����c�Ԉn�9�~SŔ0m�NG4�㤰Š�GJ�7����op�	a�������韝/%ˢ`E~F�y�޵����|��:iw�n���)mV�М�W�;�N�jf�4A�.�p�U��@�}�,T��>��V^�~�5���7�+?22�ܶ t�0,��|M��]��\gv�iרR��!,^��[;�T���V��Ͱ-���m�(ֽR���>q:��(�K�!�D(q\D�
aݞ�A�x��:gk�&!�v�u"���'A��:��/��}M6��F�yX8<ʞ�	����LL��#<y�"��1�*C�\T}}���L��E(�̊PƏ����f���Q@!��qP��6-'3{�t�M��Yo2sT3�vϻ���Aj!0��B/E��[ݒ����r)�#�=2�+�ZyY}w*d��ʌ[���7�QW���N�:�O8����.+�J��8Kz�AFWJsb:�$^��d3�>��q	�0�N�D���2��H�yx�Ϲ���RJxf5��\|mq�OL���Gr�C�y�{/�����͗>����6�%~���Ǒq��X�iM$Tt��",q���!���#1��� }Z�ߊ��w1���ڳd�٪T+�F� J2eP�����H"� ļڰ��C��K�=L���v ��p�g�ɝ�j����%���T�j�u��6���lD�5J-��0�i|�$�T�l4�8�G�%�.�^�Z��7��Ҝ�7?R�4/���-h�(���p��W.��	 Т�zK�i]u`�^�����smc]�js�]��>�����{Y�i�������,Z	s"����G^'��\ù/٧K��ٓ�!n;�G����TG����Џ���&�/����R'P+�@ڟpͱ��;��KH�`s�s���>�eH�����N��a{��M���M���ep��ĤO���:��������2�s4����)���+Rc�e65��g�#nU#>q���Rҿ>���7���ם�	ʘ�l���ْ��h����!(Z'CY3'(�+���Z�Yz�� ���B��ҸM	M4�sŶ��7�[6�&0��G\,��r]�[Lۢ�	Y"��U.�_=t;��L ��]Y*��Ԕ!�b��w�`�;��k���9^r�y���Q��{�ۘ�� �l]�mǧ��N�k����?�Hqkb��L�Q-n��jpز���V-�� m01�#�VU2��T���z�����#l��Y&�,	�d�'1�%�q�t~b���C�Ec��B~�:,��ĚF��LH�� �`��B~iۭ�%k䬣��YWf��\� �J� d��j��h-�[DE��L��3V͈��U^�S�K��L�+Ԅ�w< �wP@'���짆��#�䎓����C6�/���Ƽ/q3݀�2���f=h�qј7	r�Pa����E%I*xXĳ�8��5��ZXg���|6vV��3�vUK��%h�a�(�׹{�A��A�pl����F&p�Z�"�(%�@P3��Kt;TX��e�Bo@���I�p�����뻵>W�8��l.&- �~��#��<���:����N�]e+2x�����dI3v���x)#5k���
�}�ʫ�Q+dBl�@pG[�8�U���"�l^O˰��.U;�c+(.b�T�j������+��=���K*ViO�W>F*�O�Q����{[��il�U�����qq6�zV�zIΜ�L$�T=xW������D_��z'��+�$y�o4�G�B�>�<���F5���(��k�f����N[���[P��-�w�Z]��E5i���J��5�&a�r�9=Cଔ�3�z�5"��.��H巒�y�׊�	!4��Ű2�*�Gۦ�<�%��pye�^��V3HY�A_�uO�t&�ɘL�$0E�)[���0�X!\�-wв�'L%D��<�XK���T��y ^o�<t����)TQ�"w�ݓ��u#{Ć:�M�3mʏVJ\�r�#	"�����Q�E�O|)KVu�ޚz���Z����/4��a��^�z����E0R_�X���#SO�n�R]>�e\H��7ߣ�w��r���[Ȋ8�J;t��k�Vb��3�lB�F���P�)g�����K���������������B�NA0�������G�
����++P?\a�ē`��a�Y������N�C�MxJҎ�O	VL�YC�����'u�����W��|����G?�b �ϵ͢������$�,U0&S�5(�a�!�7�������S�e}���m�[�ⶎ�g���Qd�á�w�R�bs�J�ks8�Ѹ|�2�tu>5��6dr���}�@����ɛ·_X��^5�͔j�4��gW�l9��?VeḚ
bY0��� �����!�`��&�㏖xK�,xMm�aPfd�]5.\�����8���������3Pدen�?����8E53D6�
��:���1�((��Ðۓ��ׯ�,'K�MD�:@V��x����|
H��Ɔ�3�:�sX� 2Ծ���.��@�k� .K5*��IJ��L'{�,#ɽܱÅ�~����>`�qN�cGn�<pe�u���l�h���FK�ꃞ�	�A�����'/�R��<��K&|4. ����%^�.���DC�qWA��Qxa��ػq�ks�_^SP>Ս�'�+p���*��<��&� ���A�T҉E�L�-���k��
A�@�����o'(0`��B�-�t�VH,�LeO�pSM܈�{v.{��>��U@�%�ӏ��v�,�؈��F���>��4�o�Т�k���n��*�۶}�s��+? �a{��
J坋�֍W�|$� E� <�(o�C�L�5߰q��KW�,��W߾W,挆����ng��|���xv7��#����D���L|���}P�E��'�#���>�CVVW�##jq �!	���1{�Dpxe���x gD�t��ɂ>[��n6��f�����za֚�"m���$	������d�9�$�e�@7X�֯�����ϏGs9���wEHC��.g���i��t �9b�H./���a��-��f��$��Z��)+�s+l��!jF��d��[rY����`1l�c�,L�@��*�Q)6�c;� y�=� ��,�JҊ��̈́��H�|�b��k�'��;����S)���mǉ��L?܀�X�-�L����2�c\JR<�ed�}�8}�W���%�c�ӱRܑ6�ۖIb��4|�F��8��>�'d��ޱ{y�u����)�p���$%�`뱁zXAA�9��S�*����s�v� '�%w���{ɕ��6�[]ۛ�P�L����0�Էq�h����|���.)��:�;�\EK�8B������28,h����lOX���,�L��YKU=��ʰP�yT��Nj���rr� l�|���_�0t�2�����s���Ei��tp��ٸc����g����ZJ���j�Zl+�eQw�^���ch��\� s1m�˟(����K�H(+n"��<|��m�%2����[�Q�L�Q���P���"�ϐ">���ɵ�_���bt��V>H���8=�R�F��_<�r��舊��h%<`~�\����?����y��Y�"p�V��hǣb�;��a�mHZ�'Ҙ���Ƣq �!Ϛ^�U���?��)��u���
L�M�X�S�ۈ���`���Z�z�,�G��Iq�Cx�����ֶp_��ᴩ8��(�1QW�U�CX� �ω�_���J.hi�os
��v(鵵��Y:|?�6Cu�U��OF2��>eCs�J�l���g
V��5��я�Ǩe����ݱ*�axLЎ	w�gQUE^kX�Tԟ�/��O,��쉙H��A	r�A���A�������oSسE���:Y�n�|`D����R%b���y#��~�!�8'4���귁i�ɭ�� !�% �{iq�L���6������3L����|�8g$9��ٿ� N9�s5��x��]�k�[�e��Աr�Ǯ)�����H{&K��?�7�w�l(�V��\0h�S|�^�s�y�mB���'�����v�泣;ҒR�ϼ�0W����t�Ÿ�W��e?�x� ��7�����y���*��5s����Ʀ�?�m��r�71�a�AuI�[
w耆*q#\��IY��Kϰ&6)�Q��eBkk:�}(&ß�ˣ�����J����< ��V79N�P@��6������6
�~��$S���G�x��h�}P�L/�Xr�t��HH#�z�
l/3c)�N�>`j��� �D�,<>�E�"̊�Ʀ��}�庸@�[Uh���'k���%�[`���.��>�+�A@���MxngDd��(��TO�������M�.���֕��ۏ��������m�&�p5�)���!��l�2|/}��h�����QC������<�?���d���>�v��Ŵ���ee��h��p�gw �" Q�����~`��/i_��`�vgB#���Ix~�j+*�<P�2қ�-:�V���n>7]��k1�q3"�x��s9t�s��D%�r(,�y|��N���d�^ڀI���ʮ�4���?��%H����&�7�Iɴ��/��1���K�$��*؊�5����Ea{o��l����G3��H�d\r�}��`g��C�.x�E8o3�,;�[v�j2#7SP��qh_�����)��j3��xQ	�)�[/-X����{qb��WAP��̧͔~ K�i0g�����ٻ����=����nԅ�����wS�f���
I�3��D�4�E�Tڢ콬�qJ��Y��<���@�ӣ�*e�=ڌ=~��Қ+��g�*��!�Dz�ި�ʿ�#�;¬����Lf3�?n5��#�d	E3q�y��ų̎��GI=�Vߪ�x���6��Q3u�0�V��f@��V�g�
͓�M>©7}��ݐ��e���0>����K0���;�A��*�?�3m�b� >�,H��`�'��}����2���瓝+xc�X�yȄ���6���Tr�aS�C�J~1J�/�����A�}9N�y�d�ҕ'fU���B%{Ο�+����uʦ�<������D5���qYMz��._���/}�J�x��N�i~s5�^��#*
?(ss-V�[e(F����w�� z��v�1�*��K���㕕���q�s����ʣ���� �"Ԋx�Q3d��̙BzN������qҷq��E�=�^��Rp��8��=TuwO�i�%=�N���`�,s�x��`��X�d�;``�Cs0}�Xq���O�H������k�+������o\͋)s��?�:rS�םe~��g��$E�r�v�׻B �}����_����r���q��R'T}�#�oCJJ��n���De�p@9��~5���:�����_��vt�gc����^�/�f�
��;�v�S�+vz��l�{]f>�ܱ #B�@˨�L���_�(�n�QЖ�,�rlc�q�Z��yN+�A	a��ۓ�kG��ڭ%�y]�H�;�hJo�*�-y��`�_�����c]�D�{��,7�~���-���P�	��y]tn��(߼��b-E�	Za
��f�;B}��w~�����z#�M��NK���R�u��Y�簗���,��rb��8�6�dӻK���.��K�ǒ�P�́��Lr�7<�=dI�v+�~�U˅��>��Sֵϫ�P���%��uX'�&�z���,
ð͉��B����CP�;ĩa�B-�b�R�	����c�Ս2��`*��;B�s�qϊ���]��n:�J�o:kio�*�Rᔣ%U�]8��M�V�ݎ�Е=��-|�6��4t�����#�׊g����{:]�^E�����ӴQK�Za�
|Ts�K��f�H:����d��a�d����u&�����P|z��"B_�kAm�/��ނ,���И!�ԛ�T��C��j�<���J�����ܧ�S�4�B���8 d�mr�~���׊���\�kVu��FS�A�I`�O'$�U8��k�=�b*ǝ�3���`k7�u�l�՝ڪ��޺�
KY�8Z���c62�I���f����cph$K��@q�6NY)��]?E^Y�i�S��v���J���U)�R��e?���"�l���b�Q�P��r*f[�f`g� �y�����L��L\�c��&��$S��o�G�-J�#����sҩ,u�>���˪�e$�c~���aif�Ab_[���ȸ�#�����tJ�P޺}�E�� �*c�yW�	�]�?T,Τ��`o�Α����(ka��c���g������0�\�%x�-�b���<��}���b��y������*���_�ÇH���W��d!H*�(օ�F�:�V���kq�$�W�8�m����4L/�ʲzW���� ��0������L���!k�+M�V�u�c�&4����m�[� �(�Ta�c��u;�g�=)k�u���n5S��� !�A�B4i�e��(�����o�3�XA�3a�摠5�6�	�a�6�)�m�T:^��{:L�D�{��&S����Yq�_ԉ}��S�Q\l��V٣�Wx��K������t�Sڻ������U���Z��g��+�q�^^�i�O?��<'c����������[�����)&���I&Hj�⽝���rS�����3�(^�m�ۿ���<����v�4���/fh���AK�*�\�K�e<���ۨI�I(��":x���u[U�U���߾H��z
��b�,r����[j7�@��d�%91��\3��JhTҵ��hq�z�U����aQ��=�ϐ�)���.��H.�����Z�+���e�;y�q�)��>"��I-f	! �  �-�M^R�%�x�~�:�c�ȕ��jI١ :�DF�z=��t��G�e﷝rA�Or�+�pIOm*���)�	$���Ɓ�In6AD�G�_��1����)�V��{�n��<�=�N�OH۬��l*\�.���Ua(�]նi5��I�a-�2��֧����=}^������>j�7�$�!����c�X���#��)>���˦��?+!�U�m�f@,�R���Bۛ�ާy�-q��DG�hZ�� M�DK����k����sU`��[铁v�zD�2�t�.Ӂ��Kn�Y9_�MP���O����#�Y�����9n���tg�v��߹��\=���M*9l�4�FRF�**�; Zi�	��=�]7G8H\z$�We���_]�Y0P�� ��;���?_8�6جԕy��O�#�﫱AbUy���n-�������uצQ�[C�;���+t�d�;�F����m#���ѝp��j��� &*�0���6�~
Q��,s*Q����Α)��Wx&.2�� ��ؐ#*���Lm�g��à3�����Y�<!.����|���qD"�(��6��?�f!4c�����>WX@����9ZѤyV��i�5'ѽ뚰��:��s?*���-��j����7�m��>X�r�0z��o�i��M�t��-��];�Y�g+߾	�|]�^x/��YY���d��e�&�W�I �{H��$�y��*�`uGF-g�����~�-Ŧ���iUZ�U���{Æ��x�E;Q��s��zK(8�[�����7�K�w1�]LûP>5��b,7�Z|����ܳR&PǶK���SF ����"��sW�I�Nw�Ë�Z-�u�0��o0���Fs����� ,�m"��>�נл�t�ZSz�%i>�r�~��Q$�!�{��������s%֩���6�}E����������ޥ��T�"�H]���|�����_�ylH��.��<W�Qsuu�5��
��3�Z/a����dΒ�V�ˁyq��4�q��N��*����F;�Tt��a/P�}�$� 7�ˮʜ�xRcnb�j�5ἆ�Z�O��.a�I�!��hL;���*�WDP����"�jzao.�ꭩ/��k��r�N Y�|�o3��.��<�)�P��Eof)��ti�yb�9��!��832T�Q������S���utL����2n_2�6-p��ЕP���.Ԧ��l#Slܔ�����G����_����GΉ]�3O�`Q�Ӫ,z���\%/S�Z�`/=�^	f���+��m[@�d���R�b^�羟B����}麰��H�3	=Av����"A [9����PA}��UO���g�Q�\;]��9ww�x�z�p�% �[�a������4�*t�:љ]A<M|?|��)QpD�s�f�]�)ҹ�e�	���F����5 ��<w߃åwh��1ֈ^�.����;KP8|�� ������7u��^{ÝU��}�'a ��_ޔ�"8:3���=�<s��=�(������d(N^T�����ޞ״%Lu*�))Q�fH�{�{��Lb¯��N# l��ϙu�#�U�dc�~�*A0�G���t�J�ޑ�6���)�
��Wq���^~�MBݬ�P�.�뉟b�F�[ߋ@O��YP c ���c�+�F�A�q@>����n�k$��P�����C7R5�[��"X�sB�Z?�y�������.PS�Fc�TSn`�Y��D"�%�J;����=�X��>�
����Y�;g�%O�y���8%�DO��J�|H���N��﷈fف���۱u�X�_<��-L����yت����9!m�=�mm�q�c�<������N����=�D���/^~����	و�J2�X���L� ��ZlЧ�Hq�?)�W6<��+��|����B�T��g�[�@]��R���Yf=o�G�T�I�\ԩ�p�E�}��5lȿ�U���(��9E���תZ��/Y�?s2Ṩ��XD�%�"V�e~�8h���S��
�$R5a�;8���� %:K�Y�.^�?�;����`��B�C�3>0���t����O��Ek��<�Uj����-�TqvL��7�1<Y=�&�����e�X�r��@_��+E&Ui����G8��oEk��F��7q.P�~V	#�����έ��B�b������#����N*Dϱi(<�0���������y�gZ���'�D�xC����o(BXMP�2ٹw3�_�+�*��[���%Q��k�o�~ݤ$M�������I����nG?���R+�ܣ�a��i�0kC��TEp�ō,Z�s^5r<۾,�:ӽ&�c���pO��qs)ߣB��m��r��ǃ���D��Fk�~:�Jޓ}�'2a�s���ȍ\>KzAHz��o��?�.&��=bH$ue��	�~#�4gY�]Ji�trF�h6��>\d���qqn�(EF�m�m��lA7��">��W�̉��0�.�'4�����]��B�LP�e����V�����L+����F�۲�G�X	' U�ˁ��I5D�[�/ߎݤ1e�ϑ%S���x{Bk�E3f�!�OߊH%��
X%�`�ק��H:��������4H����z���0��Q�!�7�����Ϭ���E�L�ro�>5����6Þ���.�6��ڥ��%p��_E-J�u��͉����o��(�r~c���3t�P�p��9���r�UH���:$4w�����D&>2�I���ƫ����tW����b���}�[h�|�E�h��Ⱥ�	}�ۇyG���AB�})и�9�/�~t8��Fwe^�Z��n�����i4Z��y 2�8�b�އ�"3�]lx|Īda�cR�%J۱#<�t��be'>AԸ�2�:-�4{��.������娲���vU�ۉpS�c@��Q�K_0���"��A��0)�C\�V��E X�萎��x�|ߣ�lB ���랯�ΈΕՄ�s2��<��ՙ�t�oi���y�r�8ShNL0B�>yg������L�����/��ꪔ�8B���|�ǜ������)k�l	�k�Ӧ����;��#��Lu�>J��Ճ���h��	[��T�g<O�x�Z4+z-]�~��T�i���_i]��>2�q�9�)�&;g@���Eᇲ�8�PQ3���p@���%��<�z���p�ٗ�\��e૊3R�SPD{���F�ʁ3����j�7�c���1�+N���g	/�EA�
��]j��gi7^�$:'�w�ğ�u҃� �J!�\u�M���%=��{H�8'�^�iKC��TSв�-�"y1c��ݪx5�W�^�5mt��٥�$�ME��'B'{�Ь�.[ 0+��<��`��6o�f'���!�u��vZ��Ǉ�`�xQT��B��ZH�D��y�v�/��n-���6����9L�\�΀�|�R��*����1Lp�F,����]*T0��dv��
�\9]/S���%�Q�\_����	 ��9T�����������i��5�2���V��Ȝ��,E���!�w��\�d�Ǭ����N~�U$}٩���.�H�d��}ظj��Ye�^��E ǤɯF���0P�4�5��%�ӱ:UTD�]eE')�&	B�tD�0Q�����f ��#wE'va�	��=��$%���چ0���<W|,�^��!�p�����z�7�M����|P�#�Fz4���U[:��[���`Ye�ٻ`�e� C��s.�3	S�J7L��kD�k����7���Z
ẃ��އ�:Qli�(�0K�534@�������}9D0} cb��Z��7miV��HL����Z��$䈤c_,�M��������$#�#**�>ږ��������s�F��$]F��;�`lKӂ��D�+)w_���N$+x?�:�%18]�2��<d�x<����J'��gx�j�S,��6�ۘ�wJO��T'&I~8�1,-;�>�#S�1�R������g�9����
`<n��H��뗅�P���k���:d(��6bx$�>`���A#J�J-ܰ��֊����\��ӆ0
iO�M���!ϟ�>�Qa�4*���(z�P`�T���Г_��D� �=��#v"��T^ͺ[��-M�#�ger�NJ��ճǨ�O����Lf3>�� �(������`���[�oq<�͇�0��>�]���G=�ac��f�%i z;Ʀ��p�^AD���ӿ�������4z�U{c�j��
���E�m>/��r�K߻F��3B4��ն����,P��fgo)�B��7Xx_�??�/֨f�  ����綯�-��Z^���T˃B�&��A�pԟ��?]���n�������&׆�-���S��K�A8A��֥,�0��Uá�Ep���v��]��[��@�2f�x��Jp)���W((�� %���Du��l`O���o�P�.�0z=hܒ1���f�1��p1j���S�x��u�I�G�:n�k�SEyK���#;���:�F,V��w���U�E��mD(��.����ܙ�}Ł�W�xV�My�}�=2�*���j���0�nX#�L�Q0��}�[�*9�0b!B���)ˑ0k?"{���<���CC��XT-X�>Y��7f�c��U��A��g+ �p5)��U"�ÊD;�%$�����T��ֆ���]������LR��I�~��t+sg�P�r��W<��#�=ѱÓ���筥.-S��m�tuw���s�2��0�3��|8i���N�o$��2V��ϳ�Ԙ�oJo���mZ��J�*~��Qi�d���zcr]ة���6�߇{���p��͸�?9���m6�\�kz"S�ʖL�7F�Lr0��{E�@����X���� �����]�ne��V��O����Kn.�]=�"L �e͇=���>F�5�ū���M������g�r��;�������E8���1��A�1�l��a]�>o�7ܹ��^��N��oy�<�Dc#;�MV�����tO]8�T�t����;;�x��L̼[�1�6���6�׷��d��ǎQ�!��C�"�:ӑAă؁��_	�( �a�*Nz�c�f!.N#�_ߍJ��ٿp�<Q�č��
\%.8�#���}q�#�$i�#+����\��bŒ�ˀk���r%ǱX11=F�|�	]r�>E�>�V[l���6b>��{LL�qZ�#Ã�
Yr=��t���no[�9���3r��A�,�d�?;{��Qt��;��f�� E�������ޫ#:;�`:Z��<lx�@Ac~x��W�C>Q:P�*ڃ+.�H;,���[+���<� �g�S�
����������K��S�,P]5�$�i�IF	�u��\�E���Ja�b1���Y�UCT������	O<�HuL|�~/b�V&4��RU�^C͞����V���n���D��6nyo��.cn����
��M��#�\w���#� M�V�}\
��|�5���5�'u6���L����,�#)�UY�Fa�ޫ~����#�d���~�	y`ѻ?��	yk�^`o�GڌX�Rd�QOU�����OFs"�g�͗0ɒ 9.�H����x�C?SoI7!H��&�t2�˵$G���s-��7|��2���T��p& ֥O!a�eg���Үځ���
/�k�~lyPϽ��Y\��D0�@u֮�ă�����S*\�����x9�w�^�X�0�ŵ������C[�U)3���ӿ�N`�"�s��C���q޵�i�X}����7V�T��!:�)`N[����� ���ҷ�e�Z��N��J{��G�j%/-�m�\#i�&��񵐮I��0]�2��

?�*ЈH�Ŧ����o4��ӋQ�j{KCQ)��'�OHo�����c����8�Vѿ�:��7O�f�ŧy�Ȏ��b ����J"�EG
�T��1��ب[<j��b:C��m]�B����H�S@�Y*̓�~D���E�X�R�+`�P"��3�}�%���k�\V�������p �=�1�G�OYhG��J���4����>ܺ�{�3|CV3��Ѯ��I��3��d�c�Юv"���IUښ-��(�%��qy��fۢQ�fe੣[��c1�2а��u=Hz��z�`�Ch��d@Ep���{�P*i#��UG(��6��v����,N[�*:c�ҲMjx��S&���VRH(�7A�4��RJ�����(a_��D���A� k��[߁��X͹z��J����;���?W��7�rn拎y���F\-���|�а��"f�	�t��r~�����[l�Az���c �s�1Y���rIlg��(�H��ǽ"CP��xe��[5�����?p*��Z�|M�����bz���`��p��嗅�W�g�*��h�WU;z���C���!�5�\��󒰔:������-�ī��d��1%��P���֨e-��YA�x)�VR������n>Cw�6?sa�8&�R7>!�*p^��v,h�n>���W�L�a6@Ȃ�J8�`gC�xI��SD�����6����W�4 	�Y���7J5T�*�0;f�y$#�ð�V:ۂ�����/��2���$ۋ���t�Yⶠ�r��?+�
Ȳ2R������ �^��&K}�M"@\��R���:+�'T�n�ƈ�Z�%���5Y*>g���W�w�*�r���\�o��f^4���z�����6�����%���ssm�&z _��6�&y�S,"��)���*��8�'˼����3J�*��ڧyۇ�`��`��5U�Q��FU]QGd����1, �x�I"#	�f�s���р�Y�V����.o�������?c��^�PkG�	����s��ɛt��\V໳[H4�\���&����tS�a�HM��u}��2z�r�#���}�E�Օέ�:���۴��Ʌ�KЯp� 7D����C��D����'̠�`��k1�B�}�n\ ��xOY�)jҥ@�w︚CC�$HNL���D��#S��U�z���j��x>;j�HG�8K�=JD�|G2m@�!�/��" ���ǹ��{F�a��3JL�tB��s,]�;���_e��w_,�'�P�Þ�^�R�p�O��/��B�u -H�������6�PI#DO+�tCaA�W1���g��'O�М!��;���-As���I��U�C��RI�m]��4�^j?ҳ�/����^ϼET�[�9V�QH�6�E5�����n�u�iuǣZp� ��5���f𷙦6b�j	}�a�'�S_���C� I(c�}gtټ�� 6�#��9���^>
�wzW���vץ.�7{�k��Q�l���B>t�^��5m�7وaǲ��1�P^)"���Ӊ)$����w�������
����CSS��A����}"9>�o:���2�8wω��by�:=׈�N�epag��p�ji��L%�5O;�@
�NW6ͳdd����ʀ���k/�3b,[�a�QC��d�����h�]1E��i��z�[Y�ɶ���q��`�W7կ����T��/��JGo�+ȅ�M�)Ϗc� +#�Q�]� �K�*����0�!�*&�bA�5�|"oK�(�� �� 1� �
��\7��y֔ҧ�eޥ��77_� mR��������l�CF��	����@>X2e �Q� �KhG��T �O�t`U�L�2��z��c��ͭY�g��Zd��Z.�O�f�ą�Y�����t��K�qV�
�k���^��P]����I�}w��e\#�_��O���Q�`�+��p$�y��I��8֕'7#ѧ¡�T��c����{Ƅ�E*�j�٣>�z8�0 w��*�@l)/�����GR�y�����ɟ9�UuD�`R�����_����/���M����0�>�&LH,�7&�;���� �%�頻E�Z��
�K��Ω���c��0!��~Z ��$���2��(d�]�@���?U��o8
]V_�4V䜝���!�<-2�������ʘ罬��VçQI�v���X̟�"���sAՏ���fB~ [�?�/S&���;���(��K's�ڑ�vg��N(j�Vl�U�pO ���o���l��U��?��$&vf�d���ЛQ�u��>��"������vY'q��
�q;J���qc���iE��Uذ,?�ً'��@p:;q�J���C����G&�\�k�>��2$�K�dYiI)���c�%���Y������_N�P�a��UrԥT���5����n]�,��M�R��u-�+�Щ@)������[�@ҡXn������a6��i �L����W�T�\	�ib\�=�|�F},1{78�r��%#oBQ��J��A�S�ZP�McfQ���������4a��u ���Ḉ���vZ��,�o��a��{�;�;�}27���W���1w
��[����Q,�єل'��ފ���J���r����*�3�Q����Z�����9�^d��CIR�7CP�(���r�G?�s�̷���^$�{��� YD�2���L�iܣ2}�H�o�N×���o�kHY��4F��X6.V��x�D$�����ۋ|S�$��S��5�y�:0o��"�r�/]w�p���ow��� @N�F�����t�.�Ɣ��j��q�r�N��^�u��'V�O�n�l���i�0�����f�S�N�� ��N�^3wO3�,��Y�A�
���1�5HG�}���:�j���؀{��ӻ��{��U`On��T������]��������
ď�gP/gGo�ɥ
�0wu��i���gk���I8�n���s7�w�D��j�$��X�u�x2ƤD��Y6���T&��,uH�p1��`�D�`?���m��Ԫ�k/�{�F>�9��?�w��"��`P��L{y�D�י)B�'3}�͙��`\nvH}�>Y��%7�7K��[�f�% ��H��B��ԧj�ޞ1պe/��������!�x\B�2I�AD���+&��>�+��I�/��s1�@�c����;�V���ȯ��ߟί����Th�:��K���� 3�?����J�NV��F��7z�������a3zt���4��Ϊ�,r�˂�,ӖAT/��&LE2��w�^r<���2�w%����4��m�P8��S��=�sW�����Jcu5Nc;����g�lP{/ľ��������U��&zPԝ<g=HX2�$H����'{~���z	G��7we^_Q�g��6����Z��@i�9P�� 0�)H͈k�q�C*i�W�@�:#S?��/������g���� �+�1����S7��}��YU�b����2@�1bhl��vqεĊ=�R����y�?k��:��dI:�����/�(��mL9?-�QI�r��[Ɇαb�!�`�LZM��.ȩ�
��F�,��K��*&��n�ݕ+�N��`�;G��~حz���-[���K$�25�� r%6�y��3Oa�9Y�7�-���@���ղUn�F��V�M��3&�z��ֹ��"M'�������F"�����q�H�QCE�=�3˞e�:�oݸY'��������z��.UF3���/0<Bc֕x����܈�w��Ó7L3����Ȟ[LġQ���5�I(�6B��~l�\f_	�pcw;w	��L3��d�2�w���Q�8�r�2� ���x�'}Us"-�[�B�S�C�%�!�2��aė=�M��E��/�Ϙc]��<�u�kC�r���-^{o� ����iwE�qy�����������[����g��E�V��)��%3������KвԖ�jwl��
� �,�̿�\,S���0r��j����n��ީ:6�Վ}/YO���v꺭J
h҈�'#��`{�Bb;��Y9m����ф��|艚��p@�JD�,nv��ɴ?��V�(}��-ߛs��k��5
�~�fos<���x`7��{��GZ�W��k����},�#�LeN=�ʬ�����JhZ]VC~tF+��Z�b����EG���Ĺ��fٗ��7��bk�%�.�j�.Y����/Һ�Ʋ��'ګSo��/X=��n9�RYbA��m�)�7�Nsu�p��jD�aէǈ�����l��g��I8�٦��\�w}`�o\���ڛ�=KNњkxS*�F!L���C�ABj(�XD�I�gD�}�wXj�%�E�ΒlA-��kM��x�Mx��}��+<��/v��Bd���Kz��L����νq��$)�H)���߳y��8E�)Mr8U�"�Go�K\��G��'�~��T�%�`���[��������H��D�^�j�����ZS�J,<�Ĩ\��cj}k�}D��eqA!?d"���G�Z��d�g���[�}K��u2�!��v��A�����XOQ��U�t"r|t�;�d������c~]���!aY�6�*wv�g��K��&�RӖ�X��̔�0��B��<�f�g�L����r�yήc�L&9'�}��5�S�n�hr��l�m6<�H�߁�~o`�G����q���թa@OA�I��8Zn�j��9]��*��~0��v_��q�^�Lq֭�X�p�I=�s�V~�q�������C��/�Qf���D��`�5���*�j�N2N��}J`1��d��vWrX\Fn%J ����O�|
�
��e�1��Mk�H8�6	�oҢIZ#�sB��<�R%���m�����,?P�71��_��i:X�߫Y�
r�N����wLW���OSNV��z؛��*��>�?����wA�����ݴ��M"��p��TH�y)�ˣ}NMl��������-h���i��|@I�^7��oY��hb1�	���2>
������*�ߎ��aY��U�!�U����99����u��=����XQ�� �Op���=�̪�P�V��!x� q��� ,����Ocצ"��5j�J�;ٸ�I�:.g��ݚ�	2�K�bW��$wXB�@s��4��vKd��{A���M��Ww.PҌ	6�����`š��2x�\��eN�Aė�~���<hFE��wvG���P裼U�Kh��m	���Ϧ�.�O�>#���_ ��We8.�K,?J��|���|���,\Xm�:�G��yH1�7��x���'�iᑠ��dM1*&����|Q�ʷ�YN��$8=����� �R0!�#H�9�1wh�H&K��t��p��˜1���" /17fVo�&q���d�r�}k�
�M\F�i��_&�Q<@��n�?��s�Sˤi�@]�0��rߢlۑ�����m��NB�M8���c1 G��9Nn�jG�҄�$ɉ�Y��ǚ1�ԫ5�N��ׁK� ��jC�!���I�1�焊0��j���L�	м�\q.������_g��&O����т���&�ɣ&��b�?șr�|N�.�~�=͵�k;�'� �!�ǽ�8U�{s'�{����5PB�;S �G���9����z&H���T�#ȁ���OsȳO5�48A�o�����j���ر��=3c��	ܥ�����3)Țm�B�b����'��IQX�x�C������?��o2��1�Y�L�վ��J��M��7'$�2��~��d��p�U�]�Ca5���4@h��s��o��	a�p�O&�IŦ��:	�mm	6��� ���{S�����AΙE�7�wCz��r:2;S3V ��=�u��wS�7����+���$(TÏH5��M��d�@.eC��[)5�������#�c�X� jR��Z7z{�5�Agl�y˨�/QcɃ; 1o���%{j�S�?��s[�&[T��:A�F�B�5/yq�@�Ry�WQ�_�U���hqڏ�&�<t�4q�l�s�
a�eL�3��]dm��(��CZ�A.��V���OaJ���:
����`
["Y�	��i( �_�&��&J�ji��(܆�����"���*��X�r�!�^��L�!���b��Xu���	N�
ݵLwW\*$���㧔�8�_#���5��׼�i%���4u�:���2��'k�㝞"�쒹�FA���yg�r)�Ä�d
�#
�',���ݛ� ��r�&K��4�pϼ��E��5|�M�ؿ�|����O�Ԁ�?�#�
�+�rs\����k�b+�9$�ur�^�N���%N҇�s�6�O��M�$p�T�.�$�Qp�ɡv��-c��
�yH�<<�,:��k@n�_ 'i{-L���%Ar�B%�2�"N# ��r^Wk�e�P�_�[��9�}�ؠ�cð
����B1Mݳ�rԜB ���K�z������i�P��TI.vm�K�����+ԊH�C�Ě�J�a̒�Z׾���i%9�!_
�'̿�T���l��wZ癩c�=��K/�>���]�S�q��^Bʭ����d=��޾ڋj������6�w�*��٦� Xq%tx��2nRu#��N�5����m7]3'9��D
���3���NxO���E��9�1ҹ�Y�D��nV�L���#(��K�����Ʃ �����a�&V� �\��v�O2#��f�! eI� ���i�@��,�ѧU��VIȗ�dB�������U)��a���÷7�fl�E�"��&��i}����f����9g�5�e��l�@>�����$����%�E��w�R�(�:��#?�p:pE12�F�Y3F*Њ�fG	���7v���yL��8�)5�U!�[W� �\�9��u;���&o�Ԣk�L�~9�U����_� �G�G���bnT� �u�k͑��AG}m
���KH�L�r��7�|��Fv+!��@�%������H産h�Bt�.�����<.@��k�Jyy&#gH���7�~�/>��"�B�fW]��L,n�g����>!��[�k��ɥ[o���T1f��s��~��(�c��� ��x��b����5B?�bnMVy��m�O��("3N{&ν���s(fIs{�ln��J+ꏻ�1(; ��~ۺ���C���"�_�Q�Q��f�3i/�<u��Fp�ф��mq/So1	HYz@�\S�q�/)����Ҫ��~ۻ��U<7@~��#m.�+tX �VH)��V�~mFGo��ܪ'u�2�'N��ꚯ�����HD�@/��۰�*�R5T��$��4�� 
�:�c�c��b-��c|�S��Y�Z��J�/��BC��ڋ>#�ǥJL9,o�
Q�D�`hl�/�o�q+$ ���+u�I�ޖk�3�^��m�C�\0��/�~�͏���b8��Y�IhU�<�}oI6�k�Xhq��l`���,��y֏HcŽ�<����7��[|����p��d���J�=;G��$�Ɉ�/Ԕ�S�Uy>�w������"/I��$8���ۮN�9#�Ε�{��.Yo�ùi;�c�y��ء]HX��w��}�vB�ˈ�e�B���	Z��<i-g@M��Etz�����W"��a`.}�|h���h�*0S����G���#�Q��%��̄�{��	��rP�獾��Z�Θ���k
�n���M�|w���Й��Kdd88�V,�ќ�l�n��!��:�����_6W8� ��)EJJ2
�u ���Pp�/�?2Ł��tp���	-��q��dX��n#�Y��7#C�~oL�2�vT%����tE�"����� �;��M������
59)a;ڽv���6�$%l%!���+L�a1#WF�P��_t�����w"����0P����6cW�0�|l?��E�x�+"wN��4��"&KQ��: ��J,�-t��.��� j"Vq>�,���I߂��uk�)YwWa6tP�0�1RRI�f��������V�9�H-���ڋ#W�]�u�}���m����)�Ӈ�16 �-#��N�ps���&�h�ق,�Bmjn��X��`!�����4�r��
�-y����n8�WīϋlY˯=I봷U��8�C�K)����+[oZ�b�.���Fu��&��ۤs�����b��h�DԤ�(��{Wbx'rW�r�_T>kyIe�!���Ee��<[O-�UmZM휋�W�7��z�{x��p&ױPϙ��h�w+�b��䍣B���o���S�{�7��U�5���'�M���G�nf��)H���h���w�=F�v�n������1kFk�������8'e+�y�!�&�s�d�]�p�Ŗ�����DV�-�w}��LWT4X�2n+=7q������ A��-W�`�B��^���I#i� �3�
����:u[X�C�Y"ZX�|�%����n�0"LlU+GnK�+F���[&����}V�I�H\����b���rs!3p^~ .�ж�|��Ԏ�i-m��#��~+��[�3����?�]�n�3�^��h$�A9�������\ �t�� K� � �)��d��h�,��./�&ve���.��\�>i����~��ZS�N8�g�K
 �$�-�@�2(?�P�Q) �2Uw-HJ��5.��I��̋�Ю%>�-��T�	B��&��z-?b@Y6ł�+	�ْ�LWyEw@߲�%���CnMF��]>k�n�v ���\T>)q=�n�MvQrUj&qYca�h�囥���x�YB�\"h�圤.���E*�4���c=[\�+s��g	W,*�fqЫ�-���<�ډ$�F�Z�/@K�	��0��L�sm,������}��ڽ @J'�Y��I�Nݭ�W������#�T�l!gq]H��Z�Y:U�;�C(���S�W���b����c��N�X�ҖcmbA��n�KZo�t8��$�(&9&�&:9ØYt4�%�ֲ%ۂylB��p{[��9S�U:S�
D0��BZ�+��� �a� �j��>S�冥ci��**����[�q��ޣsv �`�F�HK5$V5���� ڡ���kc��u=�	�O��a�H�=.R�$�,����r~��&f��\��د������>m]�X� 0A3Y����'�$�K���͝s�~��2mr��p���6�1`� ��1�Ht�=hw5�T���t#�{��F�=چ��T�Ju6�Ԩ)�_{�9�+({.3�OJ�I�*\>+��8ϧa��̠�u�>j����l,)dk
���,@~˜b���Tn؀�0�+���(0�)D=��oL�G��/�.���]�8�x((/�0
�C	![x�}���'e^�� >~�!8�v���}�����{�I�w#���9�ό"bƧ4����`%�D�D�t�Dl����(Y֑�����	�t�Op_k�gf�b{�j���[0�	��U�9�ܢkr�4�8kt�7�{G33��S�p�����C܆�\h�����\(�Q#���s+R}xj��]��ϗd��y��o-䄧{o���6,��ю�X�{���JM������g�b��6i�m3��"�J�� 3��AhT�E���'������e�07{���!�EE`Վ�=)�ޗ�Ա�Jv햒Cu���K�P	3��D�ܥ��I�w]�hO�Y����Z����|"��X;�qq�����C7��&�͑(1�� ��=PF��{E�vd��rd�|�(JU�~i=��$ZГ�&U����f���=&Eёg|��g1�Y(�j��g)����EZFi�Pd����G��Q �
��x5�D8R\� �$��4o�2O/�N�*pc/R86��Lyp��E�.��*^���^�S��6A�xG$��<�_'k�_=m���ʒ�B�V��$�&f8p���^�v��0�`��f?P��/լ���U`B���asV�+n���ZB	�u��Nh��i:���������BЯ�qS19<�g����	�L{�@^>]+h��l2z�Ŭ�{sc� ֍S�c�fS@�ܦ����S#�����pX^{EC�~x����1vZ�;0K�d�eH�qPSk���D������!�B�kp�Y�\�����n?���2���M���L8o����M:i�2:�Q 	�2��GK.���3Xc�*��4A���r�0���Qz����>�B�k���옳d#8KYU�j��=�˪�}�%|�jА�= �C;�߯����VvV����品��NeM	��tC��HW	�'�AbOFX_ޥ���37��㻺���P�̼ ����P����>.���U�f��60�:�!�8�
�TNtW�ⲃbWA@��f��y�� {w�W��I�\#��.�rl��J�
�Ԍw5wح�f��T�V��f����RZ��ЌN��A�>��qQ6�~A*ي��h�m�݉ڵu2�(�F�랒��Ѡ0���J��)�ՙC[E�Oo�O�0)#�J�<���xE++oi�{�U�j���R�m��^+��j��I���d��`�T������N�`Gi?���/�y��ܑ�|g�y�����в&����}CZHoO�Ԣu&�j&����8��܍2�&�!1N:�5E����*	��ki�qpn@\����C �Hڑ��;%��a���r�?�^71��Ӭ��:t}U�,v*��jڗ�bT��o'Έ)��8�S
_���[ �9��"��L���%�t�O���ͅ�׷f婅�o�P���t��5TH����@�T�7$x��O�1���̅�;�Â�����q��^O����ǼW�sR-$y��a���g[<x����A�=���v�WS��N�
8��L>�'Zy�Yk�l�\ɢ�=�)2d���,�o���Q�]�{��O~�
$�zF�:�eA�F�=S���Ě�_�~ �\�w*�|�t����%�
�$�>���H�9���8���f���~�줗%�;c ��bAU�����0�ɗ{��$��	C�ChF�/�yIF��YE��4eX��~ش����5BP�N�v�ô��"�2V�y3�)CJ���`�`2�k�~Gxd97`X��G�闞�LUcꂣ~�5�a��V�����/s%^�%��#�A��H�6��'-�+��O���U�*���=gI5��*J���4Z��f)]��=vU��3��V5��_P���w�g;�K
	�!�T'��2d!h�w{\�n���D�ʥF�G0�2�ãf3�g��#�1��t�_\圩��q� ��X���Ǹ�Xu��j��s^�Dm4�á�U�z��$0v|��>�KU�ٜ� U�\��@��-��V����o�,�r
�FЪj9�H"��x���.3��V�2`�T #����	���k�q�82��JS)g;������`u���`g��ޒ𘃼��rt3� �X0N<*�Ƚo�Ӻ�w,���?	���8O��%4��y��g^�y���%�T�e�s�K�g苔�:
f�c���݈�<�sąY���=��bG�c��"�ty8�
�Ͱp�����w'5L[�B�6'�}��,ݺQNbJҩ���	`h���b�*�.V���/�u���=u�rwrB{_^��AF�Y�a�cȣ�v�N�.��ؖ���C�U���^Wώ���Mh��4�8U�Sظm��HHL�VK5Ɋh�i��S�8�yr�Gn�.�Fr�iN"���`�*��=�O�C��C{�	w���Î�?U3��Cu ��q�c?B V��B� ��ܬ�))���|�)Pڙ]$�I�ww�6CC"�n�.!���3���X��R���t�ͦ�U�_3�*� �3i ��m=ScGT����=]-~�����i��bpL���3�FuV��orsOm��]���P���d*��ܠ�w���U��k-}���Sa�z� �B���t6�EJ��6�r�,�834�"��2�ҹ]v����Al��*�f�AVą
����	J��/�W8
�LZ�9����́֠����"��b��̗���`�߾�ٱ<`8�"r���6�B�^w��0t6�����+����:��T@3�i�|� �C|��_HQ�i�L�_`.�����G�A�Y/u������1TY-�Ћ�n�|����e���!���O!%K�az>��h�������7�I�M�N"M7���.�����+�1�h��'Jg���.1�N���^��x�r���/N����Ց���_��<i��Y�MI>��D	]��o~2n��#A����s֑��7�2|g�w���E9�%����4*+g��<ոd\��1@ buT����y���:��g���w���_�wz��W�Ͳk����l*���(�s�2�R��?��79J^r�-��������M	�j�!n֚� J���jS�l�%�*�֛8v0�Lc�Ѷ�: ��W�?X��'،~j?�����ٯХ�(�!�i�z��y�:KR/�6�A_��x��쵴�)n�m6��:�2Tu���6���F��� +���$�.�+O|������@��(��?�?�<��;O��7`�E��9 F���,�ѿ�wE�q (Λ| ����}G�ҵ�+���48�+�A��
֬h̂ܿ�)P��Ԡ%.��l8�*�������{��{@��FTcb�?��mo`#�/(��'x�S��w��0�Y_�$DAߏ�&���`B���f�h��F����E ��Jd�z�g>/糕	����Do�j1)����,�����IH���Î��P���֩���?-gv�p���?���H�AA����a���c��)�8�]8亂����|�f�����Hf^s�xnQز��]�u������;t����3�{F�}cY`q/߭orft��.R�(h��玒�:=<��+2��ݢ"5S��
=�a礩ٽ����UTL�^)w��l��cԪ�2�Qo�f�ˋ�!X���~7�����HL,q����į����x`�!��9���Ǘ��Cާ�(�W��hӛ$Y)d�SS,g��+ӓk�?-ԩ#���O/���U�1�Gok.���|?+� �@����k��%KkC7����'��us�ֆ�'���_ZB����2����Y�e��X�xL�]�{M��Z�%�G�w��[.���ՎwϗΟ���\����ˢ���%��^c_��>ܨ��L���B�	�ۦ���� ��AvL=u�[�TJ�B�Y{-L*�u��S�rӭT���M�z F�N��M0ڙT���ʈÎY懸�ш
�d�3lQ�+]�2�T.����fp�������W|BP�����6g�|�	d�J߈�`�VmʧxԄqH��?���`;�4,��.��,֋������L�ݐ�Z�j�I��}���[!��n;��?0S�3oaj>K�VB�L�=�N}�`1�[U:v��-(D�ݟD��% �╣u��ޘ��ӟOW��2�=�	%0��n�J�>.�WF��Q��
���Hi((�+����d�b�tvD�73�b�3�����vZm���3#N��MȨ�-��{5�;�9KY�cV?AL��C���Ӫ�K�@@5kqP�o-��ĸ�ޭ�0��� ��O�pB ��M�TcV�J>{{�T���_�����7Iq�A]"f��Js�x�[U�5K'����]H�<��NX	��@N]O�SҴ^��H0�4ĵ��E���L�o�ķg�t`���
���o}�����ש4���\��M��;6J���;����* ���y�\dCgh���p��U��|����,9ɫ<J>�#���K�v�C��eD���k�v��й�`>VM�ND)�� t�D��Q>ٿ����\��;�=2���P�O���lv�O���"�J�?����`�w4^�n�%�FǔF��g�j��uG�dU$�L�YIs�Ӭ]��b+����ǀ�iq[BB�U���s��	d�0�t����f�	SL�.�8�}��W	���%g�fK[S�:�:�V2vץ�p��.}�Q%�ƌ�^�-J��+$j?$pK&3��`PM`b�:�h���"�Ù|���_f�fqj��Y�x�������n&Z�/8}C�$��s"3�c�]�Bs�?͆iN��d����NX��'&��,|0��\�'��,�Ʈ 5����I;?��(�nt
�GɃ"lv�@��̢�Q8tܟ����'���1��0<
Sck����>qo^�U����9�;P�"<}7�[vn_ӗ��n-Pm����_�S״)/(� Ok��{`h�{�����J�������I52�t�t_s�{}�W'��P�n#cR��75MF�>p�[nu4�����|k�C��f1���!˷Ԣ.}���e��"�<9C@��=-�ݶ��Q����A�:#tXM�q�x�D��N��y��*�±5�%�A� V{|�]Cޢ��F�{�i�yCD��@�[KX~v���%�9�]iZH�ky�Rb6������ϩY��p���r��Q�p�[���s�?����&`d���H�~H�oR��)K��\�y�->ŕ���U�y����}�${��9 ��,Ψi�����O��pYHZ;Èp�׫��?�G{��e:�yh]F�%���Q,���c&趸ᯙ�%tN�ѱ�z�f�)=nd~[F�r�|�{�*.��QS��U������l���������GU�N ���Zd��CTҦ�q���#'K,,�O)���ם#S�P�A9rgS�c�E��k����Mh��Rݎ9V�4��:���8RU�}��z��K�ɠ�{g�r�XW_����Z�?��w#�_�W���1�H�Te���I[!%��>��~�3���)a��5h�TౡʾDp��>A��d�I�����%�s� ax*�=��?8�|�d\SV����õ�ֈ���+��k�N*٧����xx���{�)t�Y1��,~.��0``:�a�dh����`�Ѯ�ⷍPjp������%[ا����8+����G�������IR$E�u/*e�	B�����i����G���||���`W����,�g���7�qѽ1^ #GX�s��Bla}�D韚ݵ�#;�!�����hez;��~L���SS�ߞ��8�8% U���	�Ќ��P��$���7�k`�W�Xjj�8�ؙRg�X�R���N��ICbʓ�,2�``�\D�5��6�y��k6�9����{!^���d��h��t�O* _Ȣ�6\v�(�y���LЃ�[�ΙY�!6X�ٔy.��7��FFE����������(�FC,�b�^���k�Tc��|�}�a�B�c��Uxs��Sj)N꣸19w���W����ި�4f�|��$:��.�+o�h/���s�� A�&N'�:Zn��u�2��ZN�/�s&w���䵒�[��[.�k�B�Fejz����#ý���!Ϻ@��~���m}�[��7n�H����R�����īD���?\:v�u�qc�2bM����������x��O�p�[?�o�L�ǂM䫴 ��Y733*�H�^8iM��Wт
PL�B�cL���NK��Ìb�߭5`$�7�:1�
w�E��eз
���&|����g�\Μ�y��Ͼ��s�4F�í�wwLn�Y���e���:�I}��K	M�ai�}�х��
n���V�o���Xvw�� Ų�K��P5���.�캛Z쏿Ӎ�V���Y�-L�5����Y���
����#������'#]6d����$�O{���Bb��:XxDJq���O�ء��+B�o�3�9�>[�' o�s�K"?�j(���H A��q�^ͯ�����4��|�Ib�MO���hg⣥����$���\���ڸ����Ο؉�ȝ����u3t�׌���]Mfg����0hG({���Gl+��53̴��8��i�T	F���rq|�
��4]򡈞�����w����
�KI[����D�I�?����
�aN��5�lA�k�Y���
����c��sY�;R/R ����#�l-&���_ʌ�B��F!�����֊+:.�����h��ׁ�:�Uj���� oyo�Z\���j=/
�4�h4}�ߪP��g�V���+����:�:j��/�m�*ND�w�@b@�j�F���y0Q|�8|iP�f,!��[<�"��Eg�ƞg"�R�aJ3���~�+`(��R���;��rN�'DÒt-����ALq��݋齃E�@�x��d����;�|��D�ǹ<��&�!\���/�L���H����ꂺ�V��;�4�0���H���d�~��(����}�*��:	]�yEG�+��ph\���?�����:�Gy�$��j�`Qw��3zR�u��@�������6��!}?���=�g��kQͯ4��"�/j�\��a���q�hːu�vl?�Lxn�E6� n�XM`�ڀW�섊H$B* ڑ�����B����l>*4�F9|�݀����
�W�1��aV����ۏ��5�T��5�Ѫ~S�������ٖq9�|f�� ����!"a�5��-�������ߢ������p˰�]������ܷ����E\FgG9r(�-o�'\���*�`�R!a��%�7C�7[g�~���9�0���\n�A�G�b?ᒆ4'J��#f��$Id?��b���qc[Q��^H�#��Kq��&*��}�c��P�J}Ƕ;<��E�P�	��R��Ϻ ��Wn�^��w���}�ši>����P�C�rkj͗���Z�$��u%H�0�}���IU3!R���9���^)ޔپ߂����@"�Y�`��v|=��A։RY�����e_�;1Le<�oQ>��u5���-�+��-51�QQ����=��G�U�P��bБ��U.(�*�j�$B�
 � y�槒�"ܺ&�����=%�%������,�}�h#M�A�����0����kF��W;������ѯ|�a�r�p��yÔ��c����(�@��f
��8g��a�Wo�]����8y�Ԛ����N��({���ʱ>[П��RC'K�ig'� *��&�G ��.2.*^B����;`D��mEt����������x�j�ѝ��jo�|��C��ӴOG瑿Wv�"��*�_u��Y�������c���y�c+
[���E���g�'�k���u�j��W��{Pt��4ͼ;��,�W��	j,ӭ�����9�fQ�Ҩ�w]���J�����q
H�� j��᭒��B&��h7#��ʐ��Hl�l���F��*�*:�R��qQ8�D���/q;��@P�k��� ƚ��A�� Z,A:�T��S=�ô���ϜÖ6/������ ������T��dl�d)7�،I�]�]�%�P\�^V)��N��	ߛn�ŗ�֝Z{�]�:$ .sQ@��3����������?��wR�C�&�/q��=W=�+�e��4�;h[�߫#�f�5�B�HQ���NV��¼׭O�ㅼ�<�~��"�c�t�ý;ԝT�Ppp�/�3���R��#�ʭ� ����׸Q�eL��J9=ƨ��p�x��o�R��!�IrH�����]�,�5�,"="h!1��F��n����H����
�Hu��r�cC����"�����L.�t�@ػ"B��>^��Z(Ib�R V]ު�6�D���K��/���֪r`g�W��$����&l��Ȱ���E����g`7�H�u>�<�����R��w2����E�Wz��5^�z���ܞ���lL�>�-Pq<���|�D���
U~���[��f�'?���̧]4p~��i �B:)�M$� �Ėf���WPhf|b�p��|t������d�0FAA�
�ԓ������V�8���㩹���W���ӛX���?�Y�E=z�V����Ȭ\��X;r��|��*�j�Y#��CT��2/]A�I/��f0���2잟 }�=�+�*��3�r	{!�VN�ʣ�c�:@\1M�ȋ�&�G;����*��+��z���'�C̙KW,7�A���!�{0WK��<�f�k���?w|�|)����u�/����#{A��n�mc���GG�{�����@�J���d(��8$�SD:/�Mw��~7SO-��Rѯ�5�7�MJ��Tpv�Тa]� �	����c�z���yiM�Zh����	�U���8ėO�=�p�Ou!��m��z1�DÄ�>���>o���X��]�	�2 �v���V��
�GF<}іMDX#Ӡ�`]_�_���OZ��a�isi�6.
 -|���Pܐ#9׶�K,ư�5�,����ӥ��b�xJ)B�2�ݖ���'b���	uFLJ����1�ϔ;��w����GR�����8�E,f�����w�;V��-4(���QU�'3ش����u�i�톟�\Ȍ��)ڏ\�hP~^�m�ەB�1�1�-��Y1Z̞?c�_P;U:��n&�m����j�[�,}��2�~�	�F����à��k�w=�G�s\�,g�T����AB͝T�1���#�A�m���$��s��XP����5���	�dZr,i!�'��s'n!>4+EA��2�6~6y&��'	��&�s1����x/+�HǕ��$�rbm�����(4��N����Z=-�r"Ks�%�,�R���p��X�qn=��-�㹢�>U�'��[�&� ᇄ�������c�������h$G����{�Q�s��l�>zb��晚��G4$Z��o��*���Cb*�כ��%��$WM/�/����5>	9:L�)�fͲ��2mI�L�$�P�����(>_	��;���r��ش�@��B�����F�+~s�B�HECg��"�����5Et�1��y����!�C�|@�\��"��(	[W9�ɨ&��r}e���"X�:7��=CɗUw��*v2�a"�L��W����y@�7�GQHe�>T�g+��=q�[�s�/*�jY�-��J��⯁�����d����V�IA�N���������97��m;�������錈+_�_�5=�h�����d��-O0��,��#��9�*���eFr�BL���G�s`��]t��mכ#�ഓ�?_X�~5`!2nW)Y�x"v��DE�d���X�ե������z��_hFN�ih�R��\GKϣ���065]�O�w5����o@�J.�xJ'�)!�Zj��%3���h`�j@];