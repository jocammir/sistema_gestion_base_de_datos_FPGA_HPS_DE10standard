��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0���p�?�gu:���@�6h�Bzt�7�{zC>r7��n/SA��FƓ{��1|]�ӿ&hf"��ŉ�z�xz9�����������~X��N��l2*��XҴ�qV7�QAy-���Z�5���
W,�T�=C���q�arm)�Sr��������)�Y�y���'���m��g��f_�̡]v��\�	ڐ{q�].--y����闧(0�Z��}<�.�U6����B���v��W�\m��ǐ��N��9ZBJ ����U�\�VAߋ��%ߕ�gsQ�1��%�em�L��W�������U�лcfZL_����̊o�;V��=��`,Ah=�\4�D6��`d^11�� �x�D�a)�?�&� ���K1���,,�~�4�n������A���q��&&��dfh*9�O��r"�s�Ҽ��	p�,�p|&Vu���k����LC�2�����#�;W�T��]N���Fɏ��Fd 5�5Sz�!����4B;��ψԑ�Y��FEI�t�c���jy���o��l3˞�Ba֫�����׸�xu�;���a�t�~�/���+��6�YYrY�sь���<�|?���cNK%����S`��%��RQ�;*�W��􈯭���'�ۤ'j,m Zh�š�ez�����Z��sqLCkVc���4�8�$�F�aoݵ2/�d�dT.=��~���$���Ow����B����]Xzbի��_���k=�0/��V,��+l7P��t>a޶綺r9d0��G�Б@o ��l�$�7����t�'k��A�t�
�h�JҀ��� q�Wa���"q�5|���ń��=�8c�$���>���d���Y$�I�0NX�)/d����@�I�U *���xJzQL����d�}O�����{<-�T}-a*�tr���/ê����?D���ח�_�J������r���DB�I����H��ꤢ
�t{F�l��ʇL �Hcb:�\� ���_���ބ%r�C?��l�<���tjc������ձl�*+~�h@B�y���Nn7�	y���M�2�1XK���yD���y����|7|�?�<�hv����t�K�Vkg����W
m��P���ô���Gu_�d��H �xT�����r#�!�#˕	�v'�};
�NUJaL�B���3b�Ӟ�6|1:V��TR��>��3�`�S�؉���N�i ����*/^g|/"ч����Ȅ��&V[w�?W�{���ubf��蚙��Q�hWgK��<DB#�(9�Q(9E���&^�����K}�\��ӣ���N>19�d�"����C��HD��vW��8�e>CO��Z%�vz��f9�]��~Z����II�׀���O�E>�~~��GA�#�#ڠ���K(>�6�M���M�	�5�&�b�S���h�SX���qxt/�s�,ɜ��|��
�;DmpH{���ͽ�^r�n�����K\���p3sR�|� �������ԁ�#Β-�d0�O�+?�~�:aH�A��q��Nj�R�����߉yĻ��j$ήUo����]ׅ�>�^�z���*:�ip��RcW���S��ko�'<C��i��|���P�-��Pۚ�J�]�A��A�*��l��YHS��R��撎
S\^�|X�HE�Dm)K�C�ko�bћ����=�W�B=5d���|5y>��`*GZ���/�SV�ꖿ/�Z��{7��L����?�H��'���G�U�S�[��%l���E.�p�>�5�����5b��sg�а�!D2��y(��_^��/�M��#��F��`M�������xE�W�0�	(��:�N���~Sְ	��;��\
|��)�ϴ
��'rZ|�����?�p�p�'�7�R�'_�F������Gh�C͟�����u����;'x�qR(�4�B�Z׆�m�8�mO�%��m�ڈ.�\M�3�]�[��x��4+~׍��
�c�Oj�n&ǸD,@c��Dt��bE�����)�ݦ�0ߧ:e�pOF���J���L0z�p��R"Oʫ�4�����h�)�?ޞ]�|@��(�.�6�G�d����$���۝�=���3/7��'}�N`%��3�6{Y[C�6�r��j�X����$U!)��ar�5��A"(��̋?���t����3r}�φ��֚�I�eF��ҧ�(űYo�s��H t�F��JO2JӠjY��O�!Pq����D�%v��ؕ���3��b�0� �劯Ӆ�w��L�W9��.I�����KE����u�?h��U*`^[��w�D��S	�ӦP���/�~l����ߕum�]�PԳY�f|�E��ݼ�b�,H�O1��Yva������lY\�>�˴>��LIt�]��/8��k�`���c�W����{��p̹(�A�;2ogI^��"�!<ҝ�g��=fHE*c�?�>}�jO8p�!d橩��V���#ȅ��#׆a��`ީ��6FU��b��q��*��u��o�f�6�J`/� 3��\�
kww�B��o��!����qe0�� 99X C6���Bw��>^������[B�����()�N�3T*z�L��m<�ᗒ��E^*�&�(z�?0�g��B��!�q���xe���Z�1I�6�`#c��<Y @½�j���@߯�i��+I���n�P�:��![T�&D-�����2{��4ѵ��s�
)E����>7�h�0ۉ��_�Qm��F�iMg�����Y�<�q�`{�z��co��	l�_��Z�y;�i�8�
琪�>�j����%�M��D��(a"j�^�����7`6�M!i�dr��8<7:� l!�������4fl�e�#fsJ4u6p/7گ/���N�`}5�/4o�8��4k67?륖4j�mК2B��N�a���h�}*T`k����6�1V"GKr�S8�?�hud^���.�qOؙ����R�ȫ�4�o���i��3�X����l>t��_O�����kKH�2��.!�1Ϸy�k���\����J>=�nQf
�i�F���+����f8�ׂŔ��\��ў�k�/ld� ��O%~�I�8}l�Nr�f>�J�J�i���c���%��Ų#Z�C�����͂POo��;j�OHi��Dj�NE�=�57l���a�Z� ����B1�Z�Qɫ���
�_���!4Y��%ع�"�M����Q�>a���`z3sz�g*�X�_f�R�O�
�b�����m�p����i�-�rISI�F���丧��8(�FE�I��eY�¢,���hcVｩB�qɘ��� ڄ�Hr7MD7��ۗ���-St�W�A����b�j��PK3Z�|�Q��-1c�	}+�WE`�&WdY�#v�b��4ؘ��ĸ`cg����fahncK���\[�>��jΧeי�cR
�����"�M�nu��?�;|~@����ze�Z]�����LT��Z���m�G�:C�I��I�ѳ�i�FC_���8)�����`踁JݲK���P&�m:��q��d,����gԜ�w�n����W�
�(ܫ��_�'�gr:�q��V{X���\�ň�����g[�d�cUoN#�?��}�(<>>��E<5H�&���?��hK@�Gk�V"��X��B�&��5�
�r��~�@��4���GK��a�,�I���J�e�mV�	"�ӳ��hL0,ʰ�;lS���DY0(�S	^��|B��O)	�b�C�p��ǫv|r|m�-�f�*�z���1��4�U|�v��'� z��(>�Tv����|Ӥ )�� '���)�X��u"~yO����;��{.��_~��қ��|��4�3dYYb�������D?S��|L���C� �{\ӲN�4*����,�L��ݠ�Dm(���(�= N+ݶW�Qoi{���\�~1X��\YH�!2�fxU���bϘ�.�P=S��,��'��f� �����'��7峦:E�0@o�,� ��J�o�"Jʳ�e�3�g�IoD�dj��f�3;��ۜ;��#�k�
��HPK����+ZĐ�X�X�5{��U4������ܑJ ��Xr���%�Sr|-~ַ�?N��a�#1{�|L;�(`��I?Q��%\�\ң��
��!N�#��x��	gCpj��Hk�@�Ee9D@0�h��e��R�;�ӭHӃ��O��զ����N�j�T���.�ئp��Zj�W�3���Y8��c�XV���W�O��~g���8�/��w�a�~#�Eyrӊmu2|1T%�s�A�5m�1�|�
�<%(�^���$�='�G�'*��h;R7c�;��� �S�Xo(����,�ģr%�WY"���}�B��t$�.Y!�.��`;_}��*�i��b�nci�I�NW�ڀs]7���1QRu����%t�"|O��0J�����wKg��R ��j+�p�&2�Q �!�`��6'��|*h�B��>-��.|��v�����5���b�QWd��t�Na;��>��d��QA�Qb���� w�jjfG{�Z�O���ǵǌ�D������Ԫ�F�0���:�at���P�6gV�I4�zh0�L����ƨz<���;���'"1;]��s-w6��f:�����7��K�tÁy�j�sy!��Mr&����R ��A����(�!�QC��pu���;o�3c�	�	!���x�؇�u2V��8�n�3�)���Ԉ�3�^^O��!��<k3ox���\,�-	$�d*��.J��!^�x`u񈧕w-��/��i���؝�����%N��u}b�����PI��]|3>Y"^1ˀ��'��u��mY���,ȃlhl��R�%r�/l�N
���Bk~�򲏁�4٧gb)�VJ!����\����ރ�:�=�U���\���5Ǥ��-�ˇ��k�Qӄ� �u$6N�"�o��6w�~l�u�]o��b0�q����d�� �*wr�V�䢞���{�NX1�`/��9mZ�	�g0Z�uYTj:�A�޳c��+ �wP`�}�AQ��	0�Ǚ��з��ݭ���b[R��Fd���B(���-9΄,�WH��v��r����^��>n�p�"u� ��h"�����d�4v��>B�?f�$!���!4m�<ᬞ��<,Zs��\| /�o�T����
K��\�+�,0`2��@`�F\�1��[���ܤ@�)���� �qD,s�Q%�4�!!>DvI� W3��W�>�w^	;�RSgfL�N�#ɽ��b���%���ˊS}�#�_~�����!��QR�aG�ծ跈h@��o8� �Mw�J}�Xx�J/�ؒM��|��<�(���.Z�����܏�k�d��J}�GKI��h ����$��I �	�^�ry��E~@�c��Ì�YX�W"��^:����7FGdX��յ��e���O�ܟ�D�R�;F[L�gݕ��h�����H^�VI1�͂t`�:�n�­#B��D�:�iI�D<�������o��:�'On��g��֡6���di�#�_���J.��J���y��-�A�<5�PF" 6(�s�i�sG�qCtXn���E8��쥂<��+ԯ,J:����8n*�r�������1Kr t�3��C#T�aťN�8�1�u�J�o[x���;Ou��8(#0Qs��� ��D���_ W9h�(��"��1����l�Iq�h���Z��u�b�Zl��*�P/�I#\,~A�~D�?V{r�uT?"=k��_�j�^ײƑQ�F��h�F������Y�*�d�j1)�6��eu=�6ч�*!{J�2�+�c�H1��o.�R��n�,-��|;@�s�;��'�}%�1��϶�8���N�$���b7���J�<H�B�ā^��ʒ��ޚ��0>[�DOqL��vlȴx���D���u_���,Dk[Gmo̜�9�c��-1o��m֓��Ϟo�nHw
Kw�-8�A�{CD��-��vI% 1����y��"&s���Ӄ�|RK�.�)�quX$�`꫓D��yt�w���xd��g5��˩�����iJ��A�����Fb�_���-�8����px�d����Ā���y�6�2��CS*->V!�.���8�������t�z鹊��S����f�mW?%�_�^^�q����$�~g!�TW��U"��������F�2��Υ��~4R[Az�iK����t/vb~w�^�Q�Ҏ'J��f����@��֠L!&���:���nVZ0��o�d�mw�=�&��ĭTa�����2W�F�X�O������Y@��hG2��3"湎�`#�=� ���Nfƚ൧&Q���C���XT�)�4Z��z~Οx���ɢ)���I�z���#g[�Q�<�A���[�MP�v�PY�tO�|���ط�tW�3`�*=�O�kL[!$n���/�mn������X�Y��p����"����ފ�֩�)ZP�<� ���뉸+�ުZ  ��ȶӮ�65Q�Vᛧ����1�5�	�k�5���E���x�m���YוΥ�9.!|q���"8�����~�ݛ��B�iZ�_� �O�/*�F�P�䔜���r�ڢJ�}�������60�Rf6�я���%c$�=1y�t�	@�(VV�}��[K:��<@��-��,q%	�ފ���J�jkhgl��/�ۭ&8�b!��}O:c`©_�g��ܗ��"\_�㽩ݱ�=���3*Ϳ����Q���"z-/zq�]^���IM�)Y�X�l[��;.�J���ABC����Ʌ$��kʦ��9�2DA�C�0�/[�� �Pp�JE�+A�A+n޻[����Ҽ�8�W���ڥX�>��x���Z3q�fwnP`S6����?2��#�& f�c�Z�V�i���>E�@�ߩ�G��Ŭ	��&��}m�3��Ǳ���;|G]�.sN���A�9u$==q��\N�n�ꔌ�1]�ꁧ(!�.R�ھ�7N�9���f��*�=kPEvR�Y�y������W1��aV�=�mB���`jJN������Bh��N0��ym�i�S����rK���gl��[�Z��:d���p���=nd�ڡ�4��^9�7�.�筨������*�_��6�c�>������ϲ���h̺� =$��D=P+�N�y���<�0�
�]��c��^�A�s���E��֛��d�ɏm`�j�k�.�􃿽���|�[Jgyp4�>�iؓȢ�ֲ�i���I��
�W���]��\B�緅/��q�7��/ځ����1Ҩ�V��n䥋�N��`o���u= ����c~A&� ;"����%V��@���`l�S|�<^�	%�*�R`l����lp���L�i�����Ճ���:=<�]8{������vf�� >^���3(M4"۝�
˧8�Y����ܦ��3�n�y�h��Ob+�ڡ��Ed]�<㒨*j؂���W��ɉ�@f6��߻��D���Gt��]��\] ��O)���,�6K�yq��;��@��O1@|�O+��2����X)yb��ҩ76��	%OeUk�URe��o~M��q��,yѰ�~I���VSD� ��A%w�
7����֛]�
����I`�<'�y���ֿn�Ҙ�gpޡ��������<ضlCk��Fj�g�4~�6&�~�%GJ�G��s�DV5����6:��Ne���D��͈�e�};��䂀j������i��ic�dc>�&^i��C�D�R�U�ӫ	1�"������O�;8},|O\�-���N�-TkY��׻+ì�\����2�ٙ�FI�k�QX��a��Z��x"N��7Dɟ�ܢ�
ٲ�z�&�x_��$�do<4���������a�����$NS�Ȩ*�]�E����K�^�m^5hb%'��(�b7�s���-#X�烧�ix�������QN��hRnq���K�h	c��i6`��s/�t��<#Yd:ހ���S>���D���~+�ͯX�$8z����x��W?�5�
?ԽbN�2Dx���+<x�>�nT�I�*eH9�Ħ��~����xG"�>�$A�	Q������%ɏ6:r5�ֳ��#�\�&Gh8R
�)�@J�3I�5�cS�u��pq߭{���2H���!�� &���Um�����s?�V�9��T�e	\�6�:�sȪæk	[�K��C��%�i
����tiZ����|a�L�=�=�/�;b�i�{��7���I���c��a�O��#k(�r2P��ϐ�cVՠ���m�6?��X�\�*�c\����g�⩕}�.�}��{��0C���@$��.|q�"�	ʱ���!DQ�w�[iu2�ǂ,�$`�3�����Q^���\�|�mn$�O�N�)մ�1�Ck�$���V�	��Jp�1ܳXa��q'�R/� gkp�!a`��5�����(��'�[V
?G`�z�Jhs/�e6v��t�kq�Ҷ����gb�	�t�Y��k`�2X%���&�_Rk��^C͜m���"�F�(`���em�ژ���ʢ3�B��i�
.!�M)�Q���?Ҵ4X|�z����Dv��LI{V� -���	��� ��9���
o�;�1qs���Ğ��Mrn��}ݟ}P:{�]:*�AB 
��'c)U�*vO�����HgY�#�!�h��Ֆtn#���7y�,b9�ɺ�H�:n$ �jdF��Ơ��|*b�<�NT��9W�6�{�u��l�"{�>91��c8+gu�K�3��q�-y�U�4�=�u��˳~�=�t'��h��TJv������kcI!˄Q��R�ZE��SB�."/���J"��Gn���Hv-�LV- At�� �o�������C|&<P��""�̅[T=H�v��������/�Z�y�'V��ː���3�&�)�d���A�8f�{�Y���}�l��\s�I1+�7�i�32j�0�˯�u�N���S�T���W��H4�/ ���jN��@e��;�_2���L9?���M����eN�P�E���Q;�VO���e-%[���So����Q}������ƀ��4� cCL�� 2a�:y� A��;.�m�$���Q0.�6��h�E�(���9Q,6�5P,|�=zU����@�[Q:�J6��({�VQ/ܼ�a��D}:�����hb�-�}����]�I9���_D4���QK"���ǈ��Gs��A��'�#�g,�l��������ȶ�,s�}rs���]8�����KX�k��U`�'~l���#��M��չ�w����`a����fg���Rົ�͠�U�m �\�`�b��;�\dj{Q�1�4,Pk�Q�h�yDG=[��,�律D?u���Fx���J�(��~��iu��� y�
x���b
J�u���:����#N�SgV[�$xD���n<t��Ҡ���"�"M���7�rY��� k�.t{<�Ƽ���[쑹�;d&�p�,]�B��y%_��7J�i-�S�r�u} ;�.��O��G��Əmʿ%ג�R�7qiC�E���(�:S{{��o9��C���Ď��6;.����0�@|��*x9�5�AH^`֠A�g�ܝ�(B��Y|<��>�		��G�X���R-?_�%C�O�}Y��Q��E��	9n��77}�E�K��À]���=`�c$���

�������(����A]3�7/p��"FO��/39^�������&�F6R>㋏9���5A?��Xc������J<SJF�%d$ۿ��2O=�$����^B��i`�NO��]J�".�(.9�h(T|��Wºc�սܫy>�p;Q҇B��}��i�O����a�&��3y0���e�����A�f������'������ q򀯸��W'�^[4���o� ���;]c%L7�����yQq}�r&�.W��ve���i�n��7��<7C)B�j�Z;Ēe�[DqT��V|Q�����	��|'bV"5��Q�� 0ɂb})-���Aa�%�@�ׯ�a+�u7;�6�[�����̣%h��E��B�#$�GSj|Pd�v+������E(.��
8D�o�>��N7��?MY��.]�b��&�	��m�+�S�}L��(��iIyC0gv0E����A�0s���-�~�/�`E����Rt�c��`�QUp&�`,��gq���4a�X�Rhwpo��m�Y�Y@Ոo����s�eNʢWv�M4d4��(���	�'וc� �䢄~#L�H�����Jz&�	6��W�c�˒�O�*�)V"�C)��M�>N0A*d"b�w��Q'\�0���'5��\
��V:�t'2�hv^$�6|U��H��A*y��(�}�K���$|&�^CI��-ݢL�Res2�NH��Ϗ�s`�K�)�-*�(�ԇ�j�ߚ�q<�`�{����fsיs\�F��!�����
6������_�8���8z�%akM�#'�QJ%��J��o�u�h�J����2pI�}8�>Sǹ�>m;g�r�����><�$�>�im#�a5���f�cSx��b��Er�J� b�����d-�C����� EU�	�����-��OY,/�/�O��
~��p�P�Fe!�a�O��A�G����}�i2'b��9���+�BV�*r �*��@4 �,�tL$�0<�J���Δ��o\I1_�1�63�.�Y ����b�rgd?��x��l���+(�=?�� �I�.�����eT�+ඏ�'D=f5�Ë����#6/vj�/����Q4�M��Z-�Q������{蝢�{(m�HQ5�e��ʫ#�G��7��gu�TȼW|HX	�O��#�*b#��.*0Q�h���ho!R����駎�ݫ*�
Ρ깰���Q��,�մ�!�#�S�h�Tq��L�8v�|
���>�� ���ώ�*�M0A�~�//KT�.�q�T�g�Jb���O��L0��Xb��?�����w�p{��Q��3y*��P�e��u�����ɛjj?���a����H}x֌��l��M>�f?.�9�R���Hc��"��("wMs2)ns$l�s�.-@�+���}q3xe'"��m�^�Qj�;�2���P1���T�	���#�[��m��E;�sN���?�;^�n6�G~b�r�;2i�0._߾8u���'wil��Y�x��T��!��(�}4�O�Oj�tgv������� ����q��;2,�Q��%o⎫+|�R~8��J^��	q���"�%��f�a��_���0��,�4���Ǎ��`(�6z�U�1�G�к�����!�ȿ}���e�5�L�^��U}sA���o�Z�Y+l�g��]�����ΕA����
�����x9��)���o4�O�|&�	3R[Bb�?cT��p�o��:����"~q�Z��x[r�<�RR�⯮���2��|�]�N�^��%�\(��̯���@�ɞt&�����/��d�����&�7Jr(��V{l�C�:��(��|�گ�����%l�� ����`����7.5w��~���j(�Z�×���ks�����.�t/���`һ�@�e��$ק������e���=��>d�ruG��Oϴ[�x�7�>��Lj"7�[qIB����,kz���5DU6��T���W�9���?�5ʙ�Fla�b!w�`��*Ϩ5�+�Pw�ُ�Tb�z僜�g,��[G�f&I\�
tn��߲�9w]2En�k$Ș'���l�����8<�K���ӄMuy߃pP����+z܄� �'
�sP˒2���S�ʒ2�3�
� ��$��=���X��ɌY������m����@�ib4M���<t�U�\���6`K=�9�kAގ}�D�oy
�6��Jˡ�탄���6� -"������7�4X	�_Y�l�X4�! �7�/ODKL���`��q"5w�8M3e|��yG�{���.��ʧ�/ �C�_s�*ȢE@i cn�W�[@�<��}�R�C����Oe�dB��r�V�����=�WQ�Jsĝt�
Xb�u�>��s�y�f�m�:��n-g"4�m:}�3����*~y�]����^k}2��!=�6\Ú�0�� �*��`�X[r��<V�3#����*��V��K��=����{����k�Sު���Y�mZ���cw������#�X��G��w�.,�ώ�?��x��2��#�e��1�_ğ�&�l~v�Z���D";�p��9�O�./�}"��O�ҹܹ�~?l�1*5T��[�0�A^�R�[KѾOԋ�
���&�R n*y�sK�z,k����?a�G	��p&�'�َg�3+K�I��2��ؖ�y>E���p����3ʲ�A�Y�f�vHg��� H�����T|��6�\ή��}�"I�]�?���>��(��9t�ϏS�R�k�PL�Xk�^�)�
w�����_5�@� S�'ꛍo�\�!�(5yVa�3d�� lH����Q�nC�◕�+�-�r'���#�v�Q���M��%ya'���]�t���^{�CkE��e]�1�Y�8ҭ�&��'���@��HGw�_!�s��.�^\���+;B t�r�.�sce_}�F΁���uL�#���#���"3�\=0�!>�L����4FU��JL`oYA)a�W��䒡�<�3M<���\����ބ�9�s>�Wki��%�:�"����q
���
�-ݞt�q���d�y^�ԑHb��3᫇gj����+\��n�'.�h��Â����t��d0�y-�H:{5�%mCa��㔈�֫���z7x��*Y_��n��IN�4��Q"�Y����K���|��-6��J���vy>5˴�爻U�~�7���7�O"�3%#�.~Ư~'*a�w��)K�ag@���`.�xG{J��ǋQ��A�������zG�����bgh�S�s{�"	WK:���a��yUa����Y��P�C��4���ʉ2���=%��d�u���)��%�\����:K���;G챦C/�T�k�D�{��[DW��s���U.oڮ����m+�G8��Ce�2�^@�t��Yn�f(�M	��Gɵ�
��|+0�p�n��Q�x��x˷��xK+��ېKB�#εwa9n�}p����E�$����J��+�|w�$���l��ưz�p��ߗ���ր^�� Y�.��U7/�%K&���'�
tQ�K	sHYz���@F�N�����9~;��2}�^{�����f�u_#+U�7G/=�i0r>%�W�kf s>�93Y�?��eڲ�V5⍯�+ͅ(O�Aq���i���^��-J��S�2leP�:��5�.<N\�r<��>��䐫XY����A�cĨ�>��$�����������2�6
�41���Et���vY&A������3CC�KI?��p�L���*���d�@�������Of�	�z��C���l��`iZ�y=��gPڈL�B�����|)L:=�?��)4�R�~0���@�6վ�f��h>��J��{�l��V��~f�P%���SAY>Yn�36�"�[�ݾf"]��
�q��F�۰ޫ�5�w=7��~߯SȔM��_Y���	���L�L,�#6����H07q�rИ��>ayy��KC��3
�	Cv��V�����#�	�O��6k��b�Z/m]��A���n$�! D��oD�ʗ-/�xTs��ڡ\�ж�@�q�?�<�x=��V���vҊ~Q�F�QJ�W*�-"��cް���j�u	���\k�����	��x�e����~��o���n�e`���"�+�6��(�F��S��vD/�&�=��I��y���Q1'�i
�A�Z �/��{��-'{b�O�RB���EنֆL���l{$C	j���c������J?D�ܲI��Y�~���_/���L�T�����?������9 �+M�
,�b��5E;��r�f�c!$ۛ�<�K������O�*W^ɤ���P���ʐ���z���uf��~�^��^p�4zo��=�=<�ydD�n�8�,͘<�w�۸^���)1H�aW��bpR��:���8c�@��4�>s����r�-+�u+�ױ�������^:��Y7�������rL?��G���z�Q���>�[-7�s/:�P�]��.���>Z��ϛ"p�@�%�@: �R�Ġ�啝ՠ��B6������Է�Ɖ>Y�*���X��g��G��5��Ա�O��74�S�[u�j�ڂ��
�'���֢#����pޙ:�x�B�NA�3D������+��Fb��Uļ�簸#`�E�I��z�ǵ�<���Wy�ɸ�����X�0#gOi�C�����6B�G�����` T���hY4��2���%J�o�+�z�b�IӧD7�ߕ��D�k�
�rB�����4�~NČ�=Ƒm����q?�aus�i	��+� ��,�}�2�<X���k��Ε5�'8M븗p��^�E�@�ł���S���1A�����Rj�
W��Ԓ��[�;�"vS
�є�u�Ȯ��#GdV/��~:)��o�'6&-u\%��w5,��f�e����;����Qq~@��!�
B�3صȇ�v�y�� qrp�A�0X�P4`p=���|�(v Xq������"� BƓ�R��~R1:�Jd��0�}���\��Wz�
������ɓ%�G�I�Um��!���HR(,讣d�Cj�w�
��TU��!�.�J#,�O�ʊ�~:8Q�e�t ���)s�D]�s}���֖���)�2���{l�XP��@�1Jy���ͷ�[k�:܋�}��n��r���������!��[�3w���G����!΢.&��t�P�O:���
M9�CVP�S?+ok�J �Ql90<�o�����`�Q��-�¢ o/�� �7� B�9n�00�� 1�		̼R�ߟ���В��[���#Dr��ַ�>�`y��N �1%"y"46K0��8�}�L.��3�1�$A��WwkƐWu=���ȉ����Tb�p�q7դ��x�m�g��N��|`�YpK����8�i��׽�sxp5�z�?L\�/
��ʇ��3��#$Lh�j+y�i��{(� ����m.):T�w����C���s9���X���1T������@h�-�&� ���+�`� �.[
>e�+��xc�����j;N�6J��;'�o�l*$$GZt�'��o>@�ҕ0j	��P]�vߥnȬ���`�A��r��
��g�$J�r��r����R���	�y��я���X?�3�(�-���WB�J�ZC�U��o�E����ruW�A��	���^�JluwL���ZJt+@�4�T��g�^%%�6Y7ٻC�	�Z��c^=XR��o�W�u�����"�Kܻ����<U@��P�@j���ڨ�t	C��.�_���͒bm�������v�ѐ�/~���yF�&i�#rI���e�7	rAd��V	�@�&��2�e!ҿ�7�C3S��F�m 9S��^,��P��:�K ��E6��@�D�+�H����s4v�]	�q�7B��9�<$�|h��ifkZ7�"�nw��[�>Hc����U(���o�B�`�z�� ���S�س8ɤ���0>r�e�s\N�QF��xB@��M�+#R (��퐵��W֪�2?��+�~���lX��S�u7����q��c�_W��=G�%����v��]Z$�:�c�����m��ω�"x����o�޵�Yk<�_��uH�j�v{��଄QRZ�S!5��{�΁��L�?�k���4�9��B�����|�P��c��
�a�8<C��G^֣��i}M�|�����1	�;�n�XLx��pQU��[��A�����y�|f
H`�L���Z����v���H���Z��x�����`� ɮ�H����;g,�=M�q���k�A�1��H��dDtO`�0�qe�jJ���$�p�/5���bW`$������E�z6���+$��%�K��M��1�� 6�꟫���CZ���ҷ�*k��#�J$:A�r���B�_��aU���B�i�Bz+ټ�`g�E =�ܪ �EϷ�-���7��F�c���OMڊ$��qv�b�X��n.��8�YY��걵X�Ms^°��r��Mh�	�2�>�u���S)���5B�-�~�ZH������o�iY��b���TR��&#	66? '"�uj��#g9��NY<R��P�C�p�bh��Oz�n���{�=�&=���p�<ڴ%Y�fU6�sҀAYpy��
�� ��3��7�B*{-��z'!�."���?��3�g|f4L����ܜ�����IhKW�N�i��{]B�r��ߟ ��l�T��r��'i+�^m�桁�bJ���""�J����E��u �_p
�c<��uT>uJ��h�^��g��V͌e#�Wqw�h@�@�G��qY��ĭ��y6ԍM���1D.�N3�q��HR��&����YSGjٟ���wi@��(�[�j�ua�����1��Se4m1a)�A�n�	4�mX��^����I��� i�7� �.�^�#�~?������J� ��n��5���L$(����dkD{A���<���ǜ�jJ`�j�a5��dk��'�5�+��w�����>��/�#lBg�x�"D$ I)������~���/jFo�'j��;�R�U?�� �vν����x��@����-@^�o��H'�6�v}-�5��0"��9�yB^@���t2�sҖQ���C;O	ۜ�\Yu��6�+��e���o"S�ܔ�=��',�\� �r���vB�w4:�m����q�����}�],�gѱ �P�\�Z4�!��_�����)b/�2����0ߍ9�**�^��$ߪ���N��� �0�3�VD�٤
�b]�������S��-NY��\+p�*�}�&T&-$��9�x/E^C���,*�m���&Ԫ���2q�#�4B:������jd�=�Ϗ�Aة?6����"3<W �/�͂V@d22�҃�,mn��)�UR?����L������c�~�B_ � Xm}�|�U �Kݯ4pi����l�p���U֊�T�C���n��'�W����(�>bz�/0xꊋ#�U�Wp����}��-h�.�+�i7�^^�(bC���߀^�E�������&��g�
x�l�Q�u^|杍���c�����b[�ݱƥ���!E�5���ο�M�xZ.+F�>gu�]��Y_��4�$F=@6�˜#���}�Ev#�x#���S����W�V�)�hc�EY+��gE�����ä��k�p�!79fV�#��4�\��DvӦpC)����q�!���D}���X�H@�i�����#b}yE���O;�Y%H�U��7�m���wAbZ�פ��)�lER�Y�1��^aM�Q�7�b�}|�B�3y`�l�R��7S}Sw��� �KY�� ڗ�7*�ָ!��Y�ÇB�g�.q���8�;- T^gY6�OkדJBm�]%h�A��%�`XIV�b	.�&
��U�Q�؁gR܎xUH?��j�u4Lcv��}Ӱ��#C^������#&�-��:*Y���<~��*�$D�(A��2�"���&S�E쫫CD�I`j \J�جH�N Z*���O��tF�͑J�oL���򛢈�cR�	����r�!`�� I�Y�W
�F���K}�_�O��I�ZfWg���BlMJk9�u��3%4��秋v��z^M�\V ��쬵c���2j��^�yO%p@m��,m*�<#;6EĴ��z&3�4�v�g��c�O�=�瑂G������%��-�ٍ�(��ֹ��� �6�f�臔<�r��YK�Ԋ"p�e�֗ES6����(��eIb���F����ǽ���:�>���U�����kU(U7_�Ը��P'�^E8���D�o!shv�=�^N�I�I^�n�
�y/+ �%N�����p��c׋���쑲f�u�Uc�a��Bv�,6�TG�-�<U$ؽf���w#�%�2����U��vB����8s4N�t-�0��O&��«T�����&JU�~��$�J�x�,� ��6���BZ�����o����U��Ͷ��u�/<U	�4$�}��y=��6C�O��q�+�a%Ġ&B�2L�BJϮ�E*И�E0���g���Ǳl"Vt$�C���_2��IJ��|�l�o8"�Wi���
����> X�_�2������c�s޹�%����G�}�w�vk2c��{=�S��*2<+�����f������	�Y�*=��4f�!�B����.����.4�u|B 0��V4x��<J���I��,�`�t���Mx�Z.�I�Є��R6 Yos>�Ҭ����f+���l�r�N�i;(p���s�#��'I��;O�1�Q34�^�� z�[�?;��s��4"`r�Fr��0��v���?D� ~{����
,sG�׎.!��q%���⌮	c���-Bf����&4[�马�n�N��C;���`�1J�˄��[�aE��@�<��v6�P-�]�^��*(��\����7_�s(oy,�x��Q4��P�C��70|1HV��f���ؓ��0.- �Q�Q���@���""�Is�����ǎo��EF�gP��_���r ����̃�+(O�NG�m"#�������lZ�L�9��L6ǁ� �g+^߅Wb������7�Q�!�d���~3��gr��=�+^�6-��.{��o�V�_�K���Q��;���{*Ӽ �*��/Or����HE[���;Op���[��Ăm\A �3jk�lf��w-޿�9����9I��%�>^��+F��X�]eh�Ti�U~�+�������S�s��VU�u�/Y�ϵa�"YUvA���[C�0e��A�Q�uY����ґ��F���դ|
VI��	_J��W�~���;Rp��
��V+
�B�̃"��}A��GBd,��|nCm(�YD_bA���Z���"�ȏA�0Q��\�����i�J6�f͉�hU^>�"�����/�m|P�kPdB��e�����~�
h�O抓0ܷ�2�56}���!�Nr8C���j���	��o���!�jC�S%bjm���|�n�TF i�\��1s����t��g�	��t��͖����w>0S+�z9�(�����A���қU�&BE�
�@ ݒ��=����Ӄc�	Ur���^E ܨG$Ǜ�b�4�؉�u���Cm�-�{t7�ϛux�K;���c�䊊{�����o+_���!9V�Jޗ�n{�3ݾ��$�D!�g�}F0(�p!���@2�l�|ڝ���]���M�"�\�R���PF�<98�道UCv�A�wH�#v\����W�e�]L��|1�(("b�Q}i�X?�%��#�{rF��5�A�>Ym��%Ѝ�Ƒk�����(�l�%E@�vF�C�;hu�,����Z��{"o��b9/�D㋚���q��88��x����TR	^�ˊ�[�X�Ȭ�=�n��w��G{]�i�䵾����hE�!?-����u|	�����5�Ǌ\��H�"qد=�׺U����D��SS01�E$&T�JLu{��/�y��!�����W�{rnG���*ð����E����m��jA���3���Q"��FD+vr����Y�����[#��ps�1/$pԦrj�c	���'�*��}6*�,�n㻭*��x�a,;� uOpș-��q�믓��C�\�W`��J�-XH���w>������)��	�I���)��Fۂ�p%�Mj-`�~zѓs��{7?D���S������Y�Y;��[%�g`y�c����`4wc�����[M��y�H��g-{��1�A{�[�ݘ��~������N7A(�-Z����@U�5!r�\�����p�-��*,A�J��Ww� �
�2�})M�ݟ\���ɑ>��@]�&�a.�\�50T�ݓ�Uuqe��nU
"9�g����D�o쨈�d��Lg�I�����0��1��i�m��Y8�;�JZs�.�,Z��+�%�%)����T�Q�I�m��|?�	Bk�ãg��я1�B$��I�)2@��3���� �� ̺)��֝iI�a�\L&ō腯�%ڃx�r��$��g3���  �Ж�>�k
�ٿ��_�6ӌ��N�vD�\߸zB�n�q��� �ݫ�2�U	�ب���)6;�+�W�����O1�ɠ#|�/y�E�p�5��1V>U�dN�@��B�x�7=�d�!X��EҰ�>�R��t�ً�B�j����[�!f�A:�{��	�o_Qj��\TQn#�sx��eQH,Q�I��*C�|�&�S�7V[�yCشF�?�J<�n�v#�M���u�?�j>1�ڲh��}K�s��t�K�v��?����[�E$a��&R��ls�X����e�2\���*.K���ɚk�qbp�<#����'�:��Ag���n�@h����ns��c�WC��?AB�����r�M��#�X���m�?�𧗮��g��ƌ%D�{6��%�B �����?�F����nﰏ�����:���E�2q��ی�ۚ���M{W՚���As���o���_D/��uO'W����"ΖD5��?J8����4hjdk�7�EH���p��
�AV("���?�ǋyL���Kq�Vq�˺��EQh������bP�����%��$��:��΋O����§��YL}�j���ga�A������uU-a�2d5��(��Ӯ�#��/����&��0����C#	�Mg3�pB+z�F��pF��sK�?gm9�{�#����-%�,�����TΠ�~8E@��\�&����)�|zG�����&`+�_�+�nd��&���Cc�}`m�Kg��QI,�uNi�6�Ϙ^���Q4"9�A&*[��~<�E$���,��7J�[?��*�,׹�i$X�B��[)��@��p�[f�!�8�TZ�Lq͹�f�B�d{K�y�<�d�@/Bi`���.[ �#�$[A�~y"�T�� ��|�`���V-��ff	���QA��p��nP/���2��d�K	�o݀�����_x'��Z�H�4���~��,�6����6=+�.�i�Ƈ|�����.�,�-�'x�t�>���t�ɯ�8+<��u\�#�F9|ɷ�쇔ͳ�36��=��e�Ӵ�v�~�6��L�$w�D���J���/�qS/Y}��-dg�l[h�g���
\�m!�b�r�;:��J�a��g�9�RU�3V���>+9�ۈ�����Ȕ�O�a�{�����JVWT��r�����q5�m.8�<��.�b�����dO�.Τ�(�q.���eގ�O��:<��h'�yrW��=��#��KnL����lC٣��N�%~��e��C6Ӽ�b҈!��������
��í��o� x�*�W*�V�S���JRm)�:���q��ڌ3�u�&)��Y&Ȗ	<���\t��yj����7�W��0aW��a�M�*�Ni"��ڛ+�"{��6��tr�S>s�ԕv���Q_?�TfY
�0�L=2�!��Y��Q�.��fdX��Mg=�Gf�ӓ2EI�'����W 2��ۗ��e.AP��I�Wuރ�K�"�!������%R=��VECR(��G�4X�u�U$ٸO���0��\�:C#���G��
a	$�.1x�>����8�n�6�f`��"�	��lR�`Ӳ� $0P��?��Lr�� ��JɅ�3�n��������^kF�A��>�*������o���Z���e���z�B0z�^���(�#���r1����@�?Ӈ�{�'�����$���w�m���B]����rT�So|�S��w�<��o0q�C��Ɲ��̤q�C�,��6N��;����(�Vޝ�X$�f
���|��z���=�/؅^�j�h�ۋD���]de3,+ H��y�VG��e:_�
)��>-=��g�6����Ze�>ܑ�[�� $W��u��(�%C����*�㒥�>�SۭDm8��X!��e�
������C�:��Y�����f;:?�^�Ƣ�v��6HT �]m7�̈́L�I�c�RU鏪�5R�L�M�@*$k��@�����!u4C�O!XY���qe6|w�U�u(�����v*��E!����:�ޣG��0j53	��]��i�σ��k��$|繳�,�ݴٕ��\ �����e�n~�����~�Fe������h��''�B��:8~\4�V/=�z���̑6S|7�AmQ�j^J)D_�<���d�,�̱��e[Fw���|��q�0Q̧9��J|��
�"�,�e��"��cF�{;�gM�Q�i�T��!V֓޽�N뜯�[,������5)rq��u���[�w�R���ʔw��a{v��홍,�ˌZh��P��	&��~\�#��o�a�Q��BwCm{�,7hvh"l<�C���L���D�Z���?���Ă���sdOM3� Gx�{�0{�)W�ߘ9�bVChǥ&<���!r�ߡ�8���_f��QP�+�R�ls����`�-����<{�xt����.��e)�`��J��(\��A�tb]7ةXF��J5*(��Zwv�w��D�q�~���J�����\a��!�l�	q5vNzY�`�0�bױ,y�<�=Y|�ʐ�p����-%>3�fd���'�=d�fs %�v��h%����W>O��`me� �d{TAq}�sc��o�lv59��.%�cwp��pT�9�D�s1���c��Ͳn�3>^X^W��\����]����:UlK��ck(����0+�!M�	��y]�ΊV�5�W�2���Bu�z�9�� ��]$B��u�!�W�1yn�$�	��
�:^fhdB��f���E���2B�2�oY}�B��������7�Hb��Ŵ$u��u�����㊍Gxi�qgr��&��d����.���m�gݒY��h��Z�dV{N��p���2E�%+3M����Enuy/�J�ǿ,p���ME�FAru�ڋ2B�pò�)�5��e
�u"����$Y�����6LY�c!u�Q�j���g~����0_�0����)��ݙ�D�%�`����b��vz'&��g(����6�Q��>����6��ғ�Ƌ̈́4� �n��.�����h޶Ě��k1[
�=S?�H�t?	���k]d�R'=Cl^�.��;��p�����KĪm3&L�N'����)JӠ����a!^�1�l�CP4���i��w�,)�.Z�۲`Ml9{;�2D�iN��B(��Y�~o��� ��5�۩_1x��E��?�m�3�Մ��Z��Bbo 7%\�}��q�]Xڄ��m�Þ�n�L�<���*�h��E���r�Ѽh�~E`�iZ%��yJ��?��ھk�ϋC��6���[K�0�!���k��d����%��gt4�J����V��7n��l�HMn�s������	�jI���g���^�©p��rt��%!�$/���Z�����y7]�z�� �Xxk*����~B8��{�(y�mV�ȑ��?�d�Á�D�\�����?�h(Į�v@���l�7�cL�p�7E�#��r�+�xɩ@��un����{��g��Œ[��rKR\w��2��Kw:������M��W���;>����ϖ�ъ)���-$��h�Y��"۸.Z�O�/��v��x��Z<W�����wU��YXz���q*`|a��E#!�kr˕�`�	?v�_~���g��r�� @E�FD��3�S�0`��C��L�V���t����l����iv�h>�ޞ?X��9�7��6���Ε8�(]���A���5�}�$h�� �Á�݀�_��fd	�ߊY��]���T��ke|�V`�5%����ؾ���7��-�>��d�H�C�X"�bP��XE#%L�}Y�r>T�}�x�R�8m�p������������y�tY��\��ﴕ�i	z3��H�	�Ydʵ9ݲ"5�v���L���h�G\�I�1)�����aԃ#v|�ٺ��=/Ap&�UG���[P��[�ے�&�EsQ�8��V�~	�hT��V@�
�������"�~(ubD=�3*F�S�඼��Ҧ��HE+W饮G��p�������2�g;=G7���}+�.��+fc-G1"���t=�Y�hKX~�<<X��}��dCgm�R���UFibNg����1�қ!Qo�����8�_��n��}�Tfk���l��p�����c\ �$�� ^�ԏ#Oف�a�Hd�WD��.�y̡��� ,��Qí�Ux���' ��Bd�D�m���%(�":s7�U��ن=���v����)���_��P4��RD�z��L����QR!P3�3z��]ԟ�7�]41��z>r�n�]j�~XbfEtMJ�S�/���p������W`�܍O��T�}���+6`�-o��ЯW�����K4�MY>�Y)(B�-;3W�GU)\ˣ�����o$�1�_�NR�I=�֪!����R�v�P�5F�����#��X���L9-��-+ĸ���,�+���?���1�i(��;'Т�ݪ:�B#1x�g!C^�*�*d��H���v���U\�cFg���.Lb�����:�~��t���K}��~�/O�ε�� zD:DtL�Ri�"x!���[���e��~�*�}�~f[�|M ���oQ�R@6@8�oZlA��5���)�nJ�	���/
A>�ݲ8��t�>>�Kz�g�i�1�1 �Xg�<Oobz3ˈ�*߅pO�
t+����s������9J�
�%�v�O-(+�ea�>�Tx��[ �ً�A	B_!1%X|Ȇ���(W��9�6^�����r`Q�E�Tei/N��@B��oaή����0��G:�.e��<�E�ʱ5�U8��I�I��:�2��l/��lq+�C�w�f+��1ҥ�:��T�M��d���	�����C�ؔ� \4�]=:��oቤ.����s6=J�J	w��R���9vzʌax����4�ջo��54 �3B��t�f\O0I���,�~��W��t�4U �O~NSB��2�Ӿ�iY� �4�<R�7oYѡř?ﱇ����6إO�(ȩ��h��j����C�
��{�#22��@�<J/ A�����YRq����hH��^�@q�i9OF��p�}����׉�!:m�f��F�a,�rP���-n��$�ş�,c�]H�ߧ���Y��T:�5����!��^h�xSזB��v�[���J�5�yG�����s�V$v��۪Z�`�&���fr�ier؂m8e����`*��99��E�ԥ���Դ�?=��Iߛ%Fٹ��5r���MJo�f�����+2��)D�?��_�T�7�{�)B��_�W�yw�F�_t���茋�\�xT5uE]��zf?��=���>+�$O�a��	W?�7M+����Ώ�+f�;�[Mm�kp�ƚ�bKE̚$>;�6��F3l����d�4�>`�r.��/�A��u^-������Z��۹��4^O�+r�F)��x��[?�g���D��7Ξ���I˓��g��RFT��xF���7XwW��x����
�˞㻐�����@����Ķ�~����ŗ�������9�PY���o4�Y���a�����P��@��{ut��}R{�%��b /�L\�[W�h��vS��5�1[�@��8Z�et&r�6� �U6���r!1��b�Ik�,E1?���Q2+Ѹ�,�1����H��������)��/��Ì_�E�)��Y0���b�v+ݖ�'��iI��j����j��=r���]
*>%��M� ����|-����$)�rbΈ:Ҹe��*I/������v5�+qt����n^\������$YU�&�}�|��8b.ٚUu�h����M�)3�4Z:�REJ]b��Ւc�B�!Y��+F�H�*:�,���5�S��O���,��Q!�xM�T�n��d��a�c�4#T�a�Írow�5ϟ�y�c�6��S�����?���EC) ���<!�k���]��� [C�bTCYY�f�g������W�l�,���	����D�E��D&��`��ڹZ����c�����t9b���\=,�=h?
���#)y5����H���� K�Oz'
)��V�3�C������U���$�O�t����|���N�G2*V��ƣA��Y0����s,_�	�,=C��-��@lS�pץ��w*�҅U���=7�"��NSx��b���o��r�v��t{�sݛnk���Ǵ�f����n�2�i��oZ�w�����X>�Z~lX��s#��N�A��gJz��kR�<W�n����͸U�k��Ȥ�kŤXטj��W?$�E.f�ls��n�\O�tDouԋ�|��K;��6x���aJMq�|_��w��QQxU��}`�&P#�y�
��&f���)1�h�Ҋל/�Ҋ	Z��� �c��k�2Z`�4="�E8G+�����EDE������S5O������铇Լ/�2v������W=���s�((N��*�dK�8oQ�w���rvb_�����}ӵduAPƐ,+��i�l���a�Fa����I�v?�����D6� r�he�����	_&cE��S�m��JmRy�N�!��EC�/��x���1I��3(2�j#<r���/g����͋���y�Ů.�ux��,/�650o�G�����i����pÔ���Gv~
,��f���O]�7�Q�MC��
��"����o`V��ІAB>M�h�n�>̩��fZ�H���3�\��>�d%;���t�Bz�"��¸�����>h���=~|`�P�@=/�BX,�1I��wN�+�ԕ!.�ߑ.8�9�^��q$�3���G��h���U�03�X�Z=�UŉT�h^L1��塈{A��`IT���w �$�|5݅Dz��}CdzA���73�آ'���aX8��:���2�9(sܻ ��I��٨��tϮRt�W��ʓ���$��ϧ�nԆ�oЎ��m�<���<FJ�ݏ ��%�J�؎
�[e�a�'�5�T���d��6�����G�d���G��;H�����{���^�}|�s@������:`�牲�g��=���\�r�4���NjW�	�V�˸���{
w��O�X3�qgl&M2g���@�2ܫ�nuh�rD�`3|0�94
B$ �{&xŦ˅��?\k�ٻa~U���RPc@c��R��SϘ��R��\�,�|kߴ=ꁁ�SY����`��#��8t�9��X;Fse�sUD`+JE����V�z�ҋe�Ũ�����5���'�J��8�D���+{���jd�hy���)�.�Q�N��׋͔m�׾�Nq�sFD�Iڡ�{�[q�F��ƨ����v��_o<f�	U��J��=9�
r땭ZlS�wgds�(Lf���:� ˟U^ϼ1�l	m���xםS����+*�_]��!C���H7�)�,ك�'�'�L����-_��g��I>�I$<3����|7��s��t��y�j����:�6��O�<M�5q4���%�[i�S����vז񏬥d�6��L��Pa�m��Z^����ny�i(�;&�� P��J�Ex1%��{p<�sU34�p�+6������t���(_�㡌����A!Q|����?hT��yg���)��6g�$>��-��}��&�L��L�oEH\.w�>|Z�rL|���+u�ӎ�� F:�A��Ҿ/͡��ԝj��hq����z�@�$
J�u6|���S�l��@p�$-��3�X0K�3���C�!��ZZ-��:J�E�p�����d�c����}U~����c�e9�5.���O?;m	�D�4u1�=L��>��wD<������X�N(!�,3
q�@2LT�G&'2�����	�j�28N��$]@q��b��S ����+���߾E�"pL+a�	`�޶��+}���Â�x���[�QoZ�B��"�����U֠���B�ב6�;�}�㲛���gB����`kP"�x�������,!7w�{�/���U8���y�]�'S2>�.�[3�*��09xЄ�zu��З�l�^pS������D �+�\�*�q���
1s��r�},�z�w���m<Bl��j�޾9Z�T��]N$���g��/]���s��AD�O�����{�	XzNeK0��w5�Q�D;�0�������cD2��[1t�_MO��]Rr��B�u�G*K&`ء�-�b٘l�b�K����tP���616�:@�>�?�W�VC��Ξ\�bݿE����ߍ2:3��n��H��Z?� <SQfM2�WR�������kx��b���T
��"����%�^/3~���T�����B���E��3��º��],���&+@�s���r˞����/,�Jر�Q�羙�߶��Dd|&��V�{��	��)�g�[��w�O�C�a�*�X���	�\�T}�W�i��U|�av�/e���>z��^�#��P�þ֤]���Я��,@3]+�˽y鳍X��p���D[`�~����EH�|�I���پC�'v;�ѐ�!d�禱��QX-ś��wR#�t����9�o���~ڧ��[UZ)'4���� �p��>�u&�b�z4���גA��eO<��ik��e+�v5kٌν��[���J�C< f%�:���q��R}33#�eDb�Cc� �n��:�43*�gtb���3�^�i�=���u�����k���*�)��[�Ԗ������}�	��{��ӲP��S���*yahۥB�DP���z�k  ��@Jn��P�'(M:
����;��4�݊��&�\P.��	s���G%�y��E����d��B辒!1�ߧE&hjV+Q]�)C�o�v�,���F� �E1���RΞ�h�=R\}w�Y�ϛ:�4N���@���lqZ'</�̧:�Nɟ'�����b����֬`uZ$9�>x�I������Cx���C�t]�`J��o0Q��M������"So��eF^���mFQs�&]����5�bwl���j�� E��t�8�Q\����e��!EK�:i^�e�"lH�KZ�c�X�|�9Ϧ��n!�
I�jVg��>�ܴ q�X�Q>������N9��Z� �6.�={:b9�9dx�5�ݲ���Ir�9�RU���3\���0�t��iֺ�>Xw2�p�G��I��-`O���+�w�O�A��/�B���&X��ʛH���?ON 9����6���t�{�����|��hM�����E��
2�٣E,%�Ү�y�}�#f�����Jh�̖�6v<�)'��)-����P��$`�C���72�P�\<�p���5(wƿ���[�!�O�@_N:q��\ew�\��ؤ��q�L���@R��YS6~Av�v�A��D�Dx�g�ʂ5��\�J KM��L�I��i��9C�\�ۡ>��rL��@��Vm/n���[�i=��̀��O8CU�rτ�1�B��<��o�#$H�V�0@g�u�����<"*����b����lz�p�D�Gjÿ���!,d���q�f�g�V��i���~y��E����(�4I�X�5^\��T�$*>��Wq���Y;����g�`�{L���q7D�HL�QuA�0N�IH#�Q707F��)���ٗ@Ĵ3;�G��O�{��˳�i�)�n>��X6!��@���ՙ!Η��-#y(�im{5�� �����[e���8푭5�	�a���9��$	?�A�]�`��oQƊ�ֈ#D�P0*��Rz�B�nlp���~ɁKj��T�22ι?)�IV�Io�{NY���UH����Q��p.~�+{cWI<PfR6'T��re�7�9 q=+�c%�bp{����41�!o
��:; ��oЮѭ�x�E�i�m�(%�ۢ��{.J�w�b[���g[h�t's�!�*��z-���&�bʴ�Yg���5�&r~)�`=/�pr���,̮f�n��;��D�f@���ȵ%�C�N1�C�p�.�6�7�]�u)-��GT+C�V����X��FSĴoY�Δ�'��OR\{�q��Ҙ2	�w�j,�,/�ɂ+0����2홠b�~A\����c����+�ڲ�>�sd�m���r���0�E��d�ڰ~�%U��i��h���SR8KSv�:^�����J�����������o�|�El��6e�c�Ҕh���ʱ��3E�>���=?� !�����8����R>)a�N���q������zV��8�=�{\陹V�ӵ9F�j_�dT����F]��ZԽᚬ`<���c}\q	�o���S^����Xd�;�3����s�@�7�P�Ű��W�q�!�(<TUu�</ GGTqҨ�?^��d�Oe�!ӰR��H�H����%���oILw8Mk�[W����#��i!�d�c:��p�y�ZT*!n�v�����0���J'B�{��ӕ���L�KRB��Ť���8�HFe��ӹ�D��~�^�%4�b����D黛�֮Y�CW`��e��Cv���b�Y
�C�o�u�[�W݅����u��u[���k��D%G%I���������w��1n�-|7I�
�x풎��v�/J~w*�w�����A��	y\	�q�;A'���0�a r-����A�'����{�Ҭ���%}yK�x���M�V:G�ݨ]�����e�d]66�S�+p�!����CC)�@T&	ұ.b|�W�!r����tȇXZ��#�??��eCC�tu��Zl8��M+1^<[}��o(b�_k8 �>�8���b!O���)M�Wx�^���^����EFo�G`�2D�Ht����ωr$�!M܂��_���ґ,��+ڳ��i+���m�E�;	�џ8X�u��͌��.��L9���*�:#���..4�3 3��җ�R�Uzg}.������Љ	����tЭ��Q�1��ڌŹ_���H�C�,b;�Ӵ_|�x;Kn��g�\�s���Y,��4�(L��m�<�ϳ�4|�i��2�� [�^vQ<n��e���BA5M�\�o??�Q}�4OU��ވ��w�4�����ϼ1�qs�O�?����=�Q-&�5h�4@i+�C���#���
��+�Z��S�}C��yd�
;�|;��|a5᜸�W�0�C=�~���`���ϯ;����=�#���3�Ṋ���6YuGo��Z�ݙ�}����^�%4@9:
�JI�JL���>j�m��;%��
�!!ԩ]L��:Fg�̠6�#]�	y����3*�	�`C��9].#���${l=C0BP��x��,/4����؛WA.;1Br���LC���e��;���Lϸq�*��8�0>��i�K*�7�����Yz:�p����Q�5�zZE�\/��k�:�jU�(H�r������]�L�S�d�3�`���L�]$Zr��}����8j���~����,8>�d�:=�k��h�)��g�!9=�eù��B�u"�����}���GMRh����c���t�#�Vx��@�M(����[������h#]|��(�hK�nx�]�i�7�R~yk��S�KɌ���~Oݙ��=v��6���3n�}OL�}f�%��	8��;g1�L���2̇qӨ�paX��c�\��q�;|�,%8���%ԇO-̀S����������zC� ��1\}P�Kļ͡���p��.�Gz�!���A�[��W���脫ޭCou�~Z����-�q�u��uG��R4_���į��q9�
�_��գD��n|��EX`H�������wSa����O�������of�XX3���:Eϝ.�U���u��#��5^��V.(�e!���'U �f8ק��1����d�a�<�o<��Q�3f����$}>žJ�~����W,1�/�L,�9zq����|u?Y%��kap�W�k�Uo�ev4�WE!��HoY�||���#�������7̗у�i
[<X:�%���ia&�Z��	����1)�s� �*��r�)S	�i!�&J�����$�`e�lN3sQ�M����@�%'(� "�Z�(�+�Ď�І0W�̃B>7�[iwY��Ht��{p��[��9[��Ϡ �xR��������=E��g���o�U��-p�r���3&ך<��#����c��(��h���n>#"3x��(1/���/E��C����R��$JV�j��"�&�ٝ�}�`����,��s���Sh�Xe:a�v6Q��_,��'��و�5B��~���jJݜz���%UB��C3m�F<����Mi�?*��;�!e
]�����= ��B�8������0�i�p���P!T�t7`0!� f�E����D4	(ŵ�T�zK4�[!xC�Qw�{o����K�q�K*�]P	3�AH�苎�'��;kJ��n��dѳ%6�)+V ^�9h�.��T�����	�Y0�D��U�stc��L�m��3x�+��P��jLZ�I�R�	6A)�%�Gh�3׋���H�a�Y�i��;���8~3�Ypi��6�$�
�3_���+Q/�q������I���w[���Mk��J{+p���x�.�j5���k1į��g�o�cA���n!Q����6z���4T�fJ��0��A��\H׸�DZ�c����b�8�@�8���b�h엇��Z�B+��j'���դ���z�����6Α�h�H��B���]/�= � ,2#xFwEci�x⃯a������B@#I����sU4����
�9��0;�e���K���_�>J��2��2D@�|鵿J�,��U�Z�m�3G>�6���_��a�_�M���$�4=�\)�
��|i���	�����b�bB�r������##[�"f�p*f� pMz����-ŵ@s�{:byR�Q}OCNG��4��M�]���4uߔ�=����}!���=������/���4d�d�bkpq�)�/����Q�Zdr�,B�Vč�~�{�J;�3ԻR{xt�!�n���Wj����6�1QR�����iV W5[s7�F���P����1���^�ŷ�����p�Ti\	#���ci^��t[����}m7��U;sxr0�� ���G�Zb�����<��������F�#���+�R����XEl���*J���$�˫2n�5�]��p����az���������l�<�1����Ү[�m��l֨E]Z���U`fՈ|w�?#��S#m&�k�*g��ו��A��{\u�-�
t`ǘ>�����l���K�Zj�[���YC�h��C�Q�����x*���!�����%v�qKyUD��3�@���:��w���!I��ъ��J��_�?����|G����L�ӴDb�C@�0(F������F��|�	C�j�Α._�d*m��Sz���,������l^ԟs�-oy�0�����~���1�Q�)ri��G��N[��xx�[�����I�7��b�ȁ�*O��6�/�|2(]_��Ş4��/�H/w��62��B�d&��zh���ަ��6Y�)�,,wm:5|�a;T�c���a�@�Hɵ|�4�N
K=9�������E�au�A�d�xG�RSoP"���ڭ�K��r�-%�r��N�`��=ۓ�
����Ů�Ǿ�<�����O|����g����=�IX�|�� 0�VxL���Zv̶�
_'s�{�W@�/���ݙ�h]ZF���|Zߤ<��x��]�܎`�6�l�J�/��xڪ�
��N�ZШg�)�5$[_��1\���N��ݼz�B�!1�Ҥ�s[�_e�$k8G#��Fp�D�6n�����<��Ue��.�&yܛ�s��dq�*~�홿���,�uN�_қ6��,f�ipْ�s���f�u�'���/\��p�&���{�َP����fC��������qE�<��F3�k�h��Ϛ��itr�f�R���S��t�;|�ɻ3���*�}�+K1d
ma��ۮ�@�=��c�����������3�$��]
�h�GP�M�%X���C�hX��B{)�O3M뺔��ˑ~�6O�Ѥ�y�u��aj�3't�}���a��$�k��z!_�:�3`+t��m��=E0�R��W�LJ��T�6P��>��k�Eo��1	�k�o��+n;�^-��1�3���z�:5N$0��[O���l��36��$�6���gfA�_�1�u�	���O����-W!������SD#������o��!&4 Y/X��~���u]4���25QH��1���
��tǨ�%��6�{:AF7]�:��a�)o���R���Z�=j�u����G��EX�הض�3��C�8��Df� �x�2A
mg��?��0M@�{����Ez�WK���6B5��T�7Z�r���/W�K��o�=v�!Ʊ�ma6��)�"��2�96V��.���m��PJ�;���0�>���L�����9J�_���ᵅ���M��Jo��Ì�2Gi[�1�}/p�P�(LT;q��Ake�ɯ���\1���ϰf��+���&����t`�g<�6O�HsX��p��x���(��[09{Aَ�!��VV.n�󱳛rH=N�/��E�Ha���N�17%ۻ�#����k�ƳA����\���+X<n��7�KL�u�:)�r�@�ī��	N�\�jK�!�kI8_&ʑ3���`P���`�Bh�쮢AU7��s�9��ԲuJ&~G�kt��L�S��;0�0�]U��ޏy���xe�L`mJ��!�L�fWfT(���3���m%r)<��L����k�9�0�b�U|9�R�n$�k�?����uN���Հ�F`��:?�t���lR�)�`�A�\+!	�y�L]��Vc9y@���(f<g�]�~`p�Jf��j���V��g��Ho�����]�~��t�+h� _X�P�'q���,�(�LS��	T~� ������k#�v��S��Х>�b�_��w������)���	Z���R1�t��T����Vx0�Q�m��>TX��1iTl��‼?V����6�{s1޶��f�~�͆��h�H�숍������f��^�$������A{x�V����a��}L�w2���ߔ�������]��܄�+�cY :�R��b�r�_��$��~�pa�/�+�?Y�����`�Ԥ5�c ��M|����w;I��a�L��2DJ�B�Λ<mD#Q�t�:!��LO>�|�u��]mOO��LA�A�tGtp��D.!�����v����3���{[����;1�K��rmO�z��������ʲ��1�Pj5�ia|�Z#����g�8d���ΡAw����:��x�����-��w�xus��
�_0�i������V�d�u���8w�[i#"c�T�l�Q�W��ң�ԩې�1�=�� Y)A�t�|�ԣ��9,���K�vi�I�Mi����,�rPA\�ka�����<�����������yf�{�����C��k}�xCh�c�2�;����<��J~��p^�j���[��X�%��59�'�����7]�p�([7��������;nW`�+Y]z���M]�����\�~���4��X�$�?S��T:��N� g:X���`DR �`3�6��
��]j<�+y>��.^x*
�u�T~�������;<�`g����KG�4_��nC�AV�_>���&��#fi��Ad/��s���lUv�p�1�-x�'�>�O~��
7��,N�aХE3^��ϑ����n��x�ܪ.��G��;��7NԚkH��q�<�|���,�ϛ0Y����/�_d�6�6M3����o�^h&�{�2�Rg",�	����+����J��E,���EL�P���HI2���V��P�q�R����|�4 �������Ex�������f��Ux�q�����j_��0�+��Ky���3�R�]�j�uMV��
��/	4��}����$�����{
�1>��:un˷�y1�B�=Ȯ��,��-��U�+J���O�M��*2����t��6ϗ'�$E�W��SZ��Ѩ>����9�I�nellH��~?gK�e0.�E�$ m��O���N�묩v%ww���yX��ڗG5�������M��ځ?c�g�ԇ�T�h蛸�BO�~[а(
޸}�?ZM�Gr����.UI�=,*K�A4B4��I#z#~�M��NY��kaXh|�����D=*b$�{V��M������<��O�>�_!��@پ�(K�6G6��4�2jj�z#*(�CDҋASt��/"5S�.E���<�.־{���;�L�!.j�y*+��ۈzEd`������.8#]����q=��51���{�d|WZ��[o; u8�>$��
F���*�w~�,��> v�`���8߮X%c��|�,dr_��D�\��A:��"���׻a���xo�Xߡ=L)]c�͉ҳmy��x��p�ĭ%��?h&���Mo���G�Y��<���H_�"�#"?���?;�céI�W������^�K��ʤƙ�"4A��햁N�Z��K���3y{"e��#q�v[S�	��xu������kŋ]�.q�' �n��S�&I}Ӌ�(4$ ��E�v�_[�k� ��V��ۚ�.��l�oQ��	�Ry�j}�⎅�x�s��:gr��B\��¬���t���N'<u����&.$�~i�]���¼��ϸ�+x�,7��m��{������-4+�<Ez[��r�ݜƚ��_�D�r"��Sx����$�`7��&��H�|~�?Vy&)��|\H�$Jgl,��N���]�����r�u/�L p�K�-�ͯYA4/���lx��l0�T���0�4�]���Mn�>X>|E��y��xr
��l.^�Ǐ�:w?8Nм�����ס�3gQ��#/1�>'J��m]��A�Y"����ow-�>2�
$�4��
�KA�L}�x	�������z�VoV���ײA�9#܎�q�>�g6��@��k()ʞ�5��bW-|l�1E1rU��_u�/��7��x�y� ���^ԔK^���GN��|��y���`�1{�pp��9M4Cb&���`R�qd��p2�'���KB6�(��q��I0j�o�mc"EB���
�s�zY>X����H��īޮ)��Y�6���=c�ۏש��Ӵvk#�כ"�6 E��'�L�BnB��Fi��C^���"z1 �w`&�Ό��R�;�������2cô�p;!0[G���qb�m�Z��b�$Yz�e`��G.8�b;��8.*g�z4�$s������Z��\�ژ�j">������W����V�Jܲ��%�&м��U�`=~Wn���3_���b_�:~��r�!�FP�\�^���[W����Gr[��f���TQ,Vv�����U�E�|���4Ѽq ��LG��q�TVA��/3R�"ST��6~�����(�͖rO��Sc��.b����� $�W$�����U�*L'T��uQ�{_�Z����S�����a�Z"tNJ��ֳa�gѶu�Nɮ^���^���	a��=��Xj)w+E��E[�����ɵ�-y������hyƁ�zK��,���T�mc7U��{��u'��Y�44~=���Nvt����dB�A�ԓ���XW��b�$E�:F�͙D�T�s{�Ǭ���n����hk��FF������IsVXC�}�=����!Ơ�U����ʱi��cQ���[X�WN_]��4�?`f0� �{���Q�{4[�	�ا��5ȩ8�Ҽ��)��{Њ�|'�wZ��D��p\���cv��'�����R4)q����qT/�r�`��=7�E�X���2�ɦ��FB�`�0io�;!��Z���e���~�o�2a��
n:r�������Cg{=�$���>�i���:o2�ڱ^)�;6>�n�"`�� gd�y2{���;UF)���!jk�R������>㡷�D�ڳǲɓ�6�`�fi�K3�w`C��~���i�������"��0@��E%zU�3���WS�2m3s��C��=����6�x���&�qi	����m��=����]��n�&,n(��:!N����6L�9Kh-##-&R	AU[N/Ц n�IS/�7�px/�Y0�g~������,}���wC.{���d���`��]��>��ǧ�6��Y�TR]�x�y׭��k���qN������_htH��~9�~���� ��L�ۃך��G���W,�D���1���-f+��8���l]�Q˴u��	�Z�6�6�+jb~`���m�#�f �aʸ��T���xP┦���Y�2d�TKy��Ե7y�Kw�zh+�5f����}/�P�����/P&�m�ks��ߚ;�Bb�����F�D��(�g��o��ҷ���fX��SY����?*J�!~�@�5�D�,n����fe�l*�NR�]����nr!<�µ�rW �=�EQA�^�����i��{��1�{
��Q�!�V��l�Uw�8�m���c�Z�"9hX�n�*�_��c��K�ƖRܖk`�kFK�r���W$?��&1��������1m�}��H6)ˇ�u�Nf!��4f�d�v�|
ѽE��"�!H5~'�W��ǂ�2�:�� �V�����!�����e::�1�>����xl"��?'��?����a���$'���1{\&X�����&�֏����l�֢�g��!+�}�AM��+ ����M���P��S��^�B�%��D�ӿ�o���o�#-�4Y����|�?*�K��� 6B2:Jf��Y��q��$��WB�L�gb�#bQOBeD�#�)�Zħ!�3j�	v��$�+V2?�\֮����aǸňJ4�X�+m	�H\L����zz��&v�pҐMR�>������t�Δ���]�� +s"znR�q���G���e��ٔ�r.!;�ֺ�LK��k������  W���Y��{�l�W��vM������t9B#d��x�@�3a1� ��e)�㟨df�"\� "Z��ju��y���p��Ѡ�1"6?#t\�x���z��i���C/L��Q�|����ќ8��$�Jy��z�s��hi�.�>˽.X!#��s�H��G�'�X��a~!0�=����x����3�ߑN�{��l%NÛ��n�vU�\��>�9KG;v��ܝ| ��z@�N^�3k�J�
�ի���P�/A��<;��<��M�E���¯[�]s@H��"_Q�ut�5Κ�>hd��ڻR|�XA~����+ ^3�O
#�Ы)TtT@��ƽI�|d�RI��o�v��nE�`o�v%?�Bsw�B��6oE;Z����\�����SE�TU�sWi�E�v:���d��!�-�����Hn����jsl^8^�0ϱ��0!2�O�kD���,���~�O�f�C�Gw_�BL�����(�0�:�
clS!9#A�����+�;S�|�~6��3Ð%�t����_��Lo��q~�Ŏ��(���t�D�3Ս�#�x�q�b����陶�$�5 ���kw��!�@NJ�c�����o��. s�S��/���~�P�%_V�1z�y�Is]��ݣ~x����p�����6�����?:�`�IG�A��7Y������� �����?SfFQ��nW����
br-Q��E��|�>�7\eo�&���Do�ٷ�BʘQWne_� ��(��e�U��wX�Wy��p��,�gl:n�ߥ9��K�f)�p7����(�A���z��*�v����@�ص��v+ h�!�?,�\���w�w��cQO�� ��_�~�z��	��`�=�t�a���q�z��"��>��h�Bn�o=������D�F�tm�`'��XrT�\��S*��vZ~�SSd�e������}�-�LN��H��eL�S���b���;c�y,["��Q}����_�	�q�--��e�<yr�~(����(�,ZU����X��KY�.Ώ7:#l^�&��A'�,��W�m��2@/�2gs�#�%D�VD����+�׉+G�{'���l���]	�Qǖ��ةJ�N�qmޥ+�T�6�1�2��8��l,�wE�+ŚUL��<|ې�����Ě��ܝg��R��y��N��ȌJ���͡/sj�-U��@��g��ݕATHFn�f�-ɢ/�92*�>dbR���$1��V��¯B-��8<WqIk RP#<��l%���:Ka���!���*�^ixj�O�汊ɓ u�g~& v5�գ�N }��8T��Ⅼ	m�Gl���j�`�������(����梶\�]�Hh���gವ�|.���j��@}����y�r�P�n5&[v�r>��e�S���2+9"%��׼.���-�h�*��G/Ճ�s��ᔟ �7������#�W�`i�;ӡ'�Ԩ�BbO�����e�Z�b�'�ND�T̸K�Fxހؒ���l(�"p�1rn�|مq�9�։cN���^:�+��ECl@�8:\{��	cs�k5���:n�?rqca��Z�ͺ�4�G�z�����N��S�SXsc�Z��f�h��oj̕6<8j�EܯYb�u���PV`i�`�ak���%�P���X�iURU��ð�O8�� iv��=�d�V�G>S������������7��dv�{8q߇��u�_��H�w?�u������G�;�6E�D�(x�$Sh8���M�
b?���F��V��|�=���)���6��Ov:/ ̏"�Z�6�=��dOˍ!�p��U7�_:ރ8 �)���E!��&G�ud�-����:�����Y�q\O�F�=�!����S�Ҟ��ıpe�7����ǥ)ro������3���,@y97i����P���џ�1CT[&R�u�P�Ƣ�{J�����"'�J����.����.	����t�+���&yަj8��ӯ����A��X�S��/9��5�l`j�\����3���,i��f���'r^ �d�d}4�I'��P�a�z��D��p��Ԣ;���,w�V�7��ⶇe>Љ�d�*���3�h-�u�{�X���<Z;���I#�nя�Qe��( ��bP����N�I����C��ï�m�Ç埈v�	�/���i'hu�h؈)�p��[�86y�BM�0B���Ňb����b��a����;���?r�ı��n"�� ���-���jm}�P�-�h��Na�O�&u|��,\�4�&xA�=\� ���9|��ܑa^1�� 0�+���ld�+;�|���Q˒8�M�
NG���c0�&{�؀T�󔋨�M���5��a�h8g��y�ɳJδOM�a�C��9��K�LkL8 	�k��>X"�r�����" ��I5ޣ\B�v�#�HE�")��9<��r��1�����2�� #?@��/�x\�sI� T�fB~�F�-ӏgi�+�l%����s�"�ooV�xD-k��vt~��ԕxU�1/�����a%o�m��ْ�Џ*�8��R���~;��};�}�{%a��UY��7��)�q7� �ez>�A�ۇ�j����-���������@����L�����,(�����3�~�ӒFF>ցvV\��FY}�oe� ��N�OV�xz~lc��Ϯ�ʠ�8\c��W�L�j9���[��w�R���2]͌K{Cp/��d������D䖿��MZ��!{�w��#́�+�������L���5���[`E�^*�Y���FLH�D97�Ž��gA�CS�E�G�D��P�	��ķ��h~��}$˰蟢�-��:=t�Ͳcr�)����&��U\�;���GX-�Z�#����B��`���� BM� M_2͕�aovW����e)��>��Jp��Tݗ[oZI�̠�k�¥��[@b��xc,�m�X]+p����R����퓔?30����5[Y6�~�ѭ^��>O��VB�����tO2Z]�Q����`Za"ͱ�qc~U�s�LR��ʈ7J*leg �6 ��P�q�a
E^�ꪯ7}՘5`���(E��FUH^w����,�\��a��}�X@�D�y�<×�5�Ò$Ь�RG�V�&
��ڑ\_0��YHݗBd��'\����$v����q���;b���4כp���ۡ�u�^�������j2�~��r�$�4��;�a'?��,	��xH�0�X�U10�
��n���Pv�_�h�)h�EQ�`Ć��G�!x����mԜ������C���q��"��(h 
#��N���ng���Ǖ�O�f������O���p�h]�$�@�ۅQR�C%��"�L�u��E�k������~�f$$�锍PJw6Z��������"�����.��]VĈ�ND��F���4��dk������߂����)�n��6�{&��KS��̒�O�>۽uAWN�|"h�u?g��>���G}߂i�l&[�@���P?jx�%��0����{�*E���ࢠ<�~��Y��{Q�^���O�wm��j1$�e5�����
���&�/��3�T�f��w��#�
 �>�A�c;&�k޵��l����3Q�f螕�^&V)4���#��ޠ˓煰[��Jň���ѣ���f��ڢ�!}�f��a�t��5[ޮ՟L���R6V�H�߾xH$���Z�d`�xJ�7P\��� �,-q�e+ar����QM�;r�a�$���>���08(ʅ؀��ؓm�ef�<Y2����1t�fp�Q@~D���x��%,%C�T�q"+��l$>D��>2��+%Q<�paކ �H{��f�p�Hd�����c��[8 �e$�}�{*!
����oL��(2.�!#i @�c5�>_��-�X����i�E�j����o�iv��\'�#>������_��tH{j�!��A�D���9�K��9W|2)1�Z`U�?��C���xs���B�,�G��m���٥!�7�l�@~�'���ݮ��.Uz�+qN%�1z1�Y�z�;�Cl�ۅf2���,F�j���ʘO�Q:�'�Mw����_�{�j4#�O'�'c��v���T`���-)��j/��_��
�M�u�1J��O~�dˊ�j�z6�Bz2V���_Q)�b��KU	?��𾟖*^]I�Hh1�L�vxI��o�m�QZ�E�?tO,y�z6�/l�{��_G^�)�[w��X\/��p\
�>Z�6�|U�Ť��nb�&�ӿU.d�_�d�[L���Ka��1����aӬT�[5ˁ9��ѱ����%Y����4��Ϧ�}?����8x)�/��-+���A�ĦY�t�] ��6���*�I3�PE���&�'��^U��g3�Q�L;�`���<�&��
���)����=��>j��ȫ�ݥ_J��P�(��3a����m��~/�q�L
���UE��5O��3�a�X�^.�Z#\`x*���������O���;�_z��c��٨�84�x� "�:к����´�ޠ�\���2�s*�(l�x�^�T��o�"E9�Ӂ=�3c�X#5��ד���8���m�����<��G�t���F���=o5R�H��C��d�,����K��Q#z̟�	��5�UUmk� 9�\��w�L�ٗq!��Ȗ;	u�����L�m�+cx�j�Uc�u*�c��������o4.#����p(�K�C;�&��oc��
�/��ѻ�ɿ��\D��h"~u|����N,6�FX�>�.��NW��ÌzX�M� �P��Y��%�����~���y�'b>K���x@�Lt�P.�(LWS�Vgk�����װ�%"��4A8`�+d���פg�w��(^�!�D��t�KH�!�b�ջ�\1'<���f8N�QU^�S�a�/	]+� �E>����S����o�1��k�s�^[F����
,��*L��E5�Ð���p�9� �������.|�7�[9� G�?�F4�V�-��-ē��7)||&���3U1��K�b���{��$n��0ؔ���8�;zѵ�:)�A3ɤ������!l����b��|��nH�ҧñX�i7�Q-��n�����,�\����K>KY�����TL��.���a���M���2������i��NU	��0���~L<�a%
S���EN�[��i��!���KQ�2p�p��e�`� �	Ï���qL�a�Ok*�uS�5�54��R4�����󩗱�>�N�x�r��R��(�ĊCȃ5 `���-�V,s���Z�gm���3j�)���Xݸ��<�^�E7��TN%��r��QEc̱`^`�?������O��O�A��7�R�:r��T��z�z�,W�EO�=�{d*{�3�t7�H<�٧���9����:�v�\�GfVh�â�*�[��'�i����Or]Ð�F��}�w8 �C-��R����M�&�q٥ Y&9����!kS�?pY�JT8�Q5eA��%Ux�g]�#�1��T��eۏ]�L���Ȧ_�Ύ�H������ޱ"7'��q�!�|2U:�>�"���I��R����o���}�r�Ӕ"j�f�aQ�H���]s@�p�Gu��x�rp���ʤ�M�jg�E�5X�D�q������5�e�=���|�VK�y�WS��n�A���&��Z_�]8fh�@�9���A;��?� �Q����#��$��jf��
ّ	���J��s�OZ7�h�B��:󌜄���x��5���`���Z7��\��|{f�!��@�_�{R>����f�S��(��Vi����(Rc�:�z� 0[�x�.�Q�'.d��h�ĥݪ�9�1麸k�L&��X,F2<���#��G�+:���#y���[�餢3^��0Y�g�W[�(��N+��잊VV�5��a:-��6�R�'���Gl����+{�`ƈ��~.�q�A�����Q�pA]��R�<ټ����O�=2n�!���F:�[��g��<�����:(�m|���R�Ť"�pB�MAf2�?�Q�B���tE�̓��i+�m�6���B�b�9���C=��p0�0ԗ��/��4G9TJ'?v/<C��k�E�S�B�9���>�.�#�@E�\)<���.jx�ܰm��"$xPz�A>����F�u�v��l&��FG�yM7����Y�@W}\��kf���/W%&`��Y&�ӫ�N�����j�pN0���0�������ų��$B�@�|��`�=� �u{cX:�n�c�k�r;l
�ɉt6a����W��T@��d�	i�kAJC��Hģ����1�c	D;�e�*��xAj=�+�*z��/y�P/�#�n^��k��<�^t�;�Rљ���#ܓ��_K<Q<�(ȸ�-�~�@�ǻs��ȑ#���C�Z��%%�/h/��m*w��^���z��)C���a����b�E� �\��{	�]�Z���cL��y���1��c�(cVJ����S����*�t�)�AB��رd��m��1g7N;B�o"�_�,�B�>���*�� �&��~������)C+]��Z�p�,������ΐ����3�'̡dVb�LGh�R��:�>ƧBV�[
s�.Sujp@/o�a"���]��!�&q�b�!E�B�e���D*����U�:6�ۄE�U2���������[�0�kkMxo<��J�Û�j�<�hDoW������ظ�h5Ԅ��r^�}<��̱��
��j�cQ���)��u�MP`��\7��җ���H�W����5�����fM�eȶ�*2�3�����^';�G�F��k�=�%.���ZS���FA����#���v���� ���5u��~b�Ha��q��::�f��/��3��Ȏ,R�z$��c+r��V:���B�2�>�Gg"d�=�">��,,1��h4�O����z��<���N�x\R����n� �B~��4ѥ�e�6����Q�P�;N�5�.bC�i��}�ei��{ �!��rt�$;�-��� 4ݣ�t�T������q6z�nb��-�a��X[�g��C�Jc����cV�񌼥8����"���͚�'U��5;{��P�!��׽��2�}}u��rrO�g&WlK����LJ�ܣD��%�����i��"�}b���(cE�S�B��1 �`��[zA�;Lu&�����py&�&FzW}E��htǇГ<�r��L�Л�t���ˏ�?=���[�9���Eȏ�� �F>`_��YԖ�6�uV��c�'+@�Q�A;���H}$�E�*����0�����IZRc�
{��I̖J��y�n%;\�^���=��!�y-n�W��I���2(�˫�+R
�^��"�IF���L�F����m�s� ��ふG�T��9���>A}��Kc8�t��}�RB�V5?쏳��tk�S,6E�3C�p����{g��22��}iiM���
�C?�/�Uiǥ�����<�YP�o���눅��\x�ߛ&W0O�¹4o��=Ě2�#��s�
���5)���z��9.�s���eh��F����ǈ�U�7�$h��R]?_w��D.T��3�����.�^��Y�]���+p��kLZ�gR�Y��8!��%-F�i��!#}��/4�Ð�dM:^{����~�^ٵ��tsіi[ �\�u��J�R\���*�.�5��/t���/��Q�h�����YJ���qA�I�#�����b�|���Ik�S>ES�,nЊܵ��r]J<��%a��?�µ�s>����j��ϘmE��洏���9U ��ڨ�*_*׋/�-O�.$��=RZ|s�Nm	�:��jj=�|�n�ic��y�V�m��*ϑnT��]?T.��9Ϸ0G�4K��kQ�uF��[1�d������"��ys�h������4��*����k�h2�J;kpy��#���IO;�@N
��'����4��S���[�T(��-�����
��I�	���t��`�o�y��O�M1V�$p�Mm�#�/�}XwZ�����(Dt�̻SM�;�����.K���j���f$�;�}Mڭ�g<���D�j�t#��(?�jcc5��
�~E��bNy=ΝW�|��t0�����[ʅ���bi=ܝ�M�)"/�)��PE��9��s�O���k�^�[���=�j�l����;c-���C����d������`�}�z����y����\�(/�E�k�9�=������]=x�f>	���P⸑f>��:w;�<��s ���vi~�\%�ML�3�v�5vfph~y��ɯ>�?��Õ��U�38���2������~����g���F�0��iTf((�E���2urq�ps�.{	+8�	X��oņ0@w�4]��ה��1�r���*+��]�7���bgF"0��1tL�=�r�K���:�U�l���e5�&�@���|�/�`��;r<r �{1��/�ܜ�(]c�2jJg���c����<N�s'�ί��K,.N@��O�=W���fيۓ}��K�j{��z�*��R�9��u9�R����({B� fR�8*�m�^�`9O���X�~��=��y��i�o�>��X���X�����"�?�P��;�9
��Óa���F2�["-Ϭ02J���1�@trB\��
�CA�9�Hp%u���ae]gJM��}.�,UX�i?��KRR��~T�_c���*i�W��B<D~rjE���A����5�h%ql�dz��G'���v3Q����;����1�I���No*붔�K�����r/��M�SY�F@��� :�6j!���ƠƝ�g�[�|�@%��S!4D��4v �v'4�}JԲ����R����%�@+���Q�q4�*#mDUl���#����I7�#.f]L?]D�Q]��1]4*�`�B0�\u	���;8ZxV!��Ɨ�Nt��-ʝ�ӭB�U�C���F������Q.ii�<�I6���3g�/���0)<�0��Y2w8Oi���j��,l+!O��~�����A��3���3-�h;|}6�ñ>��j���z��Z2���
�ʑ����#�^]��@@�'i}Z����7�(i^x��j�� ����2���
T��#Y���>^����^�֡X�e*��*|ep�,�Y�= >��ڽZ�I0j<�#�Xf�	���mW��Y����$
��g���8�Ŕ	��ƅ%�LVa5Zaf���
��j�{���3$�vk.�ݎ`�}a���u�O�`u�	RQ�)!�i��b�<���6��5�	D��ڧ&�]�$إj��8VE���Ww�@o���B�К=�r܃��2M���Nu��b_��?`K��K��k-+���[VV\����N]�rA��`��a�Ϳ�nP����VAMn���5#�H�H���$k�p#�{bfT�m��簛���BҺ~+#_x��{��|����ձ��!�Nਭ���Cc*�e�[�;+��M�U^oJ~��S�����J�'~)>\5ҪA`���=�ƚ���`Y�
n_�4��;Nl��HZ~R�_9@�Dz�� ]e����J��+�7_�w���WL��N@ٵ�u��UJߝ�
2aL�z����H �2�-b�ٳ����ʗ�w�(������^��T�HW�D���{>� �F���8�wA�F�<����HT����Ǐ��< �ݎ��.�(],p)EUc|S��}��t�	�RjW�6L(�� �j$�c�|�h�!�^����[���Jչ�t������ۓl�-���-��pǁ<��RM"x�N�g\����?_���Ǯ��Z� ���J��'&I���۞n��r*@݁M�ѩ�ʲ\e��k����"�NG��1�8+|�e��t�13N2+��R�X� y���k���]vȳ[�3������.ȕ�6�v|E���wQ��Ρ�Z�a[���s�w���]D���vF�}��h�b@!���������Q���.��{������|XK���a����i ��aJ�ʊ8�/w�U~�yJh�Q�l<~��Y&���d�՜]��7��'�;�|A�B&�gGK��V,Y0�v����ϼ�p��?���d_Tr��CA{P4B�K)'�}�rZ��g*��Ol'y|ŝЊ@��a"L���2?���ٞNx4L"�A_.9 ?C�uT�#e����O晑���(!vl����������>�p�X���$�x�$F|���)'#�%�x,M�{���Ӌ�bGv�K�5/;.c˳=�h&��),
�Ɂ�S(�ī�N�ڍ��sJ��z��h�ӋO&��O��1�qBٻ�R�h:̵���\�N E�#�8zy�4o5ޟr�����A�ݗMG���Q���k]�d�A��:ЈE����t���Umq�#�"�T++�B�xY�*Z��z���D�!���pQ�MO��첗�W;���7F�[Þ�4}�ъ�J��ޖS��Z��uſݿhU.�֭!m�P�`�]`�~���g[�1ݎ{�#7	�J1s�.�`
��BH��j靦��Ք|Z�Tʲ�U���C4�ia��2�=��Y`���0D��ITY���
�9��q/�87$��Q�,�/�J~v�Douj�|��'(�&��lb.�|x��QGW ��\�IA�W�-��v0ˌ(\�*�[�Gj�����ˬ����</�( z�w���uC{E�p�T_fA�rx��bȣ��c�ˢK��U������k�E��s�!��^��(�h����it���q���G�� �T1��\���,Q��0�.�ӛj��{�� N����}B�6t{�;�yE��+ϋ��P�Q�uG��O�G�k�X91A|�t�j��)+��5D���
[���]e>�ߣ@r��\�0=3�$h�H=p�R��+����<y�P7x��p��#�`N�W�� �Z}֧3��Ӳ����E�!�ޯjp�aѣn-�]�UE����SB^e��G�t$p�P:I�Z�$1l��W��	#;mC#O|=��Qv~ޣ��;SkTGT��Ό؂�^�j�U��ĞxS���/
p��!c��
Ǭo����7=wA���ɚlN��K��!�9�,z��h�F6_u������S���!'1��64�I���1t��%}Q�p�!���PH|y����G�'��b,.��ڤ��v����,C��r��.7�c9ܲ#�_�H�?��[j�H��`��i)�R@A���E��&4���%mk�����U��M}zS\�@�z�\���W��>E+}�;��X��2H�{/�_�=R����s�<vS�U��V���8����&w��.����E��m]�;��e��Ƣ������0"�י�h4n���U�u�
i#s��G�G>��?�yB���,&�I���"��y+����l�\@�a&�O��/>��b)�y��h��v�<��K�5�	����D�m�� �Q�\*S��}a`�J���g�������7�0��j�c�\��O�2t�M��h�~e􀶈�8eQ�K"���+�jz�P�T3!���xB�2���ھ���A0Z�4�?W@4i�T7B~E<Z���Kht�]=�?m2��=�K�W�=�𦓱])����	s���A�\� ���1�Α):ց��#Ø��k�n�b=l���잷G���2���g������9����f%3C�~��\f�������1�w�do�V��0vA���u��,�w :h���2�j�g�)#�jQ)��L��u��R�����!>�uDW�I	�	sDw) �d������p���C���ج�Uf Z�a7����|S�}`���<�'?�'M�|�T��ŬVAJP�ǕYY� ᧓��4r�Y�cWߣ��ԃA���
gr�d!x�-�H�R�����&��hT��N�=	P�w��@0z���Q������u&��gd��"}��3"H<qxp�@��<��~V�'��ɋ=�Ƭ^n��an=�tv:�ſa����hO}��1q�F�t�@>[v��P��BB'O��)�&@�A=}�3��7}e8O������/WQ��N�(��Q3��t����@��^u4�
x!%���Q��9W̟,_��٤T�%��f[��9�±|�a��c#�I��Z���2��O�׶�R{� pȷQ�/��6s��c!�[�����2��Bs��\w���R�̅�.���4Mx���j8(���ԣ)Ԁcc>�.d����0-��}�9ִ��@|cz����&�ȃE,<��=R�PoNR����Ә� ���9�*c+�h�LT��`>m/���__A�_���)ue|I` �����t�@�+9b�>+?jn�A�e��H� k5"�ǝ1!%�i�]۸O�mE�*LdIѠ^4:�%�Cr�d��=���z������v�<Lһ�Q�_�_��t�g�J�ѺX�F3���=�2Hr3"i�ɳ6b�8�ہ��A�.&��������<�4�Et���:���/��Ep�ҏ@���)v��7�z�@�6KK��gH�n��+yn)��猊Lz� Os�	�R�Fpu"�N���hJdp���ؘ@�V��QmL�g���:3u.W"����ӹ]�!��e<�!�==�p�8X��w��<{`�䣸C5E{p��9f��)w��%�"��xNݯk
�7,�Z��!u�v<��#W9�z����g;�Js��]B������&�y�1�
�ݏ�Նz��t
�r$�AΨߋ������� �uQ��[c�5:�#g���W:��$��[j�m��?��_�ٍ�uJ~b��>�'ɇM:�#*�Ǚ8�VE�n�De�1���Ƨ3Y���_�Ҹr�#N��a�IY��>nM��n��	�*��vE^8S�~���l�³�/��DFj�I�|W}�ƙ$����-I���,�1��-��jo��dߦ$esK��ƕ�	��"$��z�5�H���t)P�]l}hQ���g��x��z�\�8;�6�ek�>Q�D'U[W�(�&�W�!T�)A�ddMV&�����/Z4$���93P��[X���;OpM*��ㄛ�yXt˥���ĥbɈ�]T�e��{sۚd�F~�������n�~,�N��ͨ�B:4��tNo�q�#������@ͧ�w�D��y[��lNC���Q��b �>�&�;��L��[��+�:�_ų^�B"̉DrG(y~�{�s�6^w����x�s���������y�FH~�~ ��"�4��QE9����^D�v3�)
�� �D�u���oj�g�1�`��m��4Ϲ�!*�N��9�80��#X%I�uykv�~�L���Z�"���a����M�qU��AR���vZM,�*3$*��i�� 
Pݔ��_r��τކ���'(�������,=�T�ݧ�DHL�s32���@���;��f@��V��]�D���v���	k�>�U��q�Rc�f���'�R����0�6��;�T�i��q�w�nݻ�����_x�)�w�*�Xʋ�n�h��t�z�����ޭ��Ӕ����6v�e�E{����Y�U�f�-û],6���kl�#ò��pz�餹~˃������Ō>�9{TYR;�'�V��oQL#=[��R�~�>����(�Wä�����q���a���R�Eш1��^��r�H&Y	�*V4�n�c�VL�Ld+����m�@��8�۱D=��&�°O&R���~�xh��*Ҥ1�+8H�|�.���$}��"����G�(�|Y�
���}�L�o$l'�V�:Yc��-�L[1��X���:Y|�bdI.K���O��,>º��t)܋�A���2EovG������Rs�`������%�?3�S�1}v��9��W�aDr�Q@�Ȥ�)/�p>����խ�bRћ���86
�Y��6��b͆i����G���zR�[��������/��53�j�AU����'vHĞ�Cq���6�4�ۥ����n�C���r?V���
r��?�V��A����!�b�ݒq������?�6D����Ӂ$0?G���ܴ��ɦ���v/x���E��ͭ�T^��陡L�<v��^#?���;A�p8k����.>�@�d���go�_?�[T����`��䃜}�%k������c�%�[ ��@x���&�_�!W]��K�r|����L��8	��`TZF>f��r�/�;�NgB*P���qϣ6�g4��	�L����>�c���I�7]օT�X��dp�)��mH-����'��̃�����UcMv�=�X���O,��5w��>umF�ѷ.<����J�X�,l���;�nug%1���W'�+fFw�u��Ac��WV�����'E�7%{����/�}�O�E��!F��LMo��M�
 ^�����-������p��w���85��q�n[���f���q�-�a�tr����:Cw�����wr��5j+�����7E�R4��sfiŠ(zc�����K?ڶ���R���7��͉a_c���ʖ��{,�A�x,9!�Hӹ���)���~��b����<X;tnv�x�ԸpʳY�\��8�V��+�UV	�RG#v�Y�ݭ�)l;ѹ$�Z��~���8��q��d��q;W	��G�R�\'�b+�:�0�� Z��R��I��Н���KA�-Án���̹Yzp�*��Df\9vL���׿F��W���l	����")�5�A��H���9~�;�[���0x�U�P:6 ���J|�6�R�vTfu���h� �JX�X�:lnM���U�?VQ�9it-	I}떇?�%x5����ِ�Y�tth�(�A��M���c��m�ӏ����t���3LD�~�DX����0���#���pf�R��������8`��va�j- P2��D0�bg��ϻ��Z�`
St�P�?l�=?�0[�$��.RU�5�i���4��]s�Xݮ�i���S:XZ���К��M��G/a4 �p�u(x����^�ۆ���9�6�\���Ӳ�)�2���bN����LAREH�q����QT*(�ԑV�}��@~O���i8�J[~���^$W�����(�B[|���� /U��������� i"�U���~j�n%АhfP
��Jr|�A%�c�H��_g.S'��w��	ň�����z�#c�����1��du.��ۘZ�Lq����I�#�xmd���Ǜ q�D�7L�҆M��X��(-��B�E� �g�K/��@���5�gi{�N=� ��� �y���1�gA/y����J��=v�E�����s�/�,���3�r��,W����� ���R���&�f���	�i+��߁hl�+`O����V%� <M�_n:�Udȁ�[�o�y}���`�'^I-f�M�!��l�)��̶ptD�תx��Gn|N
�߰9W:A�x(Ÿ��wg�4��q,�.�i���H�����P�ףK?�8��iE��fi�V,ն�~�7���8�K����m��}
[�px<oU�z���=k�8��j5���� =�e^ 3�M�d�')�k9�d��ЪEE��ɘ�/�#�.���R�l�0+��G�#�������r�ewrÒ��O������#��+JRԸ�t�Y�� ���A-{���=�A��s�I�ޞ߬K3Oש���eK��#ɔ�f�L�/�V�� $}dM0�2^����A0qJ��]�X44M�߰>�u����Zblh	f#Y��*&3^�Z��}-z�Z�ƞ8#6NH����B�U�aH�S�8rM��V�28k��Z�)+AfѰV�0z:$���q�1��u/��w�A��*����י���3���S_5V�Ƚ=
ۼ�w}& �G�z�½�:O �:�$�<(<&
�ώЭ��+7�T'쓰�N[靼0���X���렼s���II�_�St�����(�@�b���H]�)��}���E���,�.c�7���}:�<�O�~�,��ާ�ʆ�f�s^�~�@jKG����քi���g'����n%ϰ�&���yL	�G�1���J�[G��Y�N*�x�E��_hʵ*���1i��*��6��#8��X�L��|�e���rrd�$o�6�۟1�)ڿ���E`|zg�4�t� /9�+NHFgbI��F7G��C:�`�����i��NhUk4X���7�K6h�kZ;�q�#a��\�]�ZT���ݩa�'�K�l������ۿ�9h�D	L�d�!׻��9l_F�M�'n�/;Û��'��<�"wV����䆿T�`/��Τ�ZQ�K��z\�Z:��qY�e"ϷL��<&���ZKm��j���~uI�L�E�Ԑ�*�1�o�_m�2��{��p�X����9_{߇|�Ok]�ގ�����57\,����9����G�ve�m�$��K��;�Q��x�ys�Ji�.���fY�?RDX��!b��l0Yj;C9���G�*��P'��0��=ħ1_��	�])�#�2��� ��w�@�q��I���h��������:gX��m�:�`�������`i6e���w���8DE��ѬV���X�^,�hԈ��dѥ�k����/;ǃ܆�pc�g����l-ޢ&a��®.���t�Q�M�.�s��6]��y����
�c��g�����R-�Jy��L|�Oȳ��!�������s|.���{C�&�
+n'%����\�EbO$��T�4�*���(��j=V9�WP�kw������=��Z�dz��a[�^w|b��2�g��4�0ó����n��,O����W�	�����*/�=TD��{���ʶ2�+a�0�}L�{
Z���Z	Y)�r�l{�
X�SO	�Q3�,|qVP�X%��R���5J�2�`W�Z��%~�$�A���5�Q�ʃ<�/��vz��]���YK����:�K�@S���Z�ݍ9�l^�XÓ�RG��:*�!�M�i*L�O3a�ঁ�VC&
�,F�6ː;�[��Ҧ����Z3�[�f�oʟ)�Z��?f��٘�mj2��F}��p+���<Zwg�K!R�L�%�_s2�:N�ƨ,��sE�'<�����a���3<m�����,`�h�r	�Y��}�֠���������b_΂���2�- s'P����F������z|�h�G��V��.,"&��_3,�JB��$���0�iF�$:��� S� :x�˵)�����O@9��ʙ�c3�CS�=�=���թ��=;N�&���Ww9�'I�#V�CAb�L���L0 �O���3��ϵ'S-�>�w��p��E��@N�9ٙ]@�a���y^c�������#���(�@cEfd.�_~�Uk)c���qA^�/�	lvU�Ш�N?6�(�0�侪������S .O�b������?ߤ��ʎ��ʭ!��a�J;�\dcS2���1�xR
mn�+7�)�ɑ������gi��bn6�[c��G�Ov]a���b�0�U�(ئ�B����@o��z�q�	/��<�ʍ���Q��*���v������[>����cK��_"�����0|����9�" .�yf�W�t��548��j)�c���4���q0Ȗ\s�#3t���Β�X!"�u��u��� ����mY��{�%L���w�4��̝��Z��4;�g���b�U-���]a���f�%�`[��1 ���>���9�th��l+���a��J�r�$��
>�E�񑗌��5l��i�5y����S��z� �T�R��U!�kߗ������7��%@�}�5�t���4���h=��>:�S�K���3�¼FB��@xXD��Lݟ�m&Q8x�+8hqr��~5��3�P�[�XN�%Xzr�ND�����f�@��a��F�AX:�$���r��Ĳmf��8\9t�̠����S�JO4L�e��O.�'�Q�W����h�$���)���my}+���ޏ��zFOo�(zߩ@q����M��#���3j]�;)m	��6D	#p?���a��ʾ��&��g�,����B�J3U�]ߨN�b6))�f~�����E�v���N�ю��҅`�hZg-�e\��5ʙ�'.�@0�	f�P��b4���i����[^�P`��T���J{k�*S��,�H�z'����7�,�X�����eS\���
�g��6�\QRu0��:9C�����o�z�'���ߊ^�o��M��� �P7�v�ا�]��_^��qCl��צY
�yu��>+O��+�S�B�ºs�
��P�xt0�	?lmW�P�ib�>>𸣔pa��f9�^�BB�"#g6D`��+�֟s�7���(d�CC%M�1��A�*@����V�'S��ۏ�<R����:�;<�	g��7[>�::;۰��{�|�O�W���L'��k��0K�K�g!�L̃���.�_�3�&��ǧ�?�� fR���0�������V[�S�>��A��D=�8�,f��p��~�U�Z�ѯ��'c����/�rP�͍!\H�Q��>1f��S�|̵Җ���f���$<ڱY�#���$keeJ��|LB2�RsSv�1E
-���CT�k��G�Y�\�ͅ�q�e�'[h��c�Tz��;��LR��i������kI�S%˭og�<�)��_G��	fX{)�:�c
�ͅh�8�{T���<��8|~ޟ��l[�Lup�^&�aϪ��le<��1N�f<����W��L�·|��__�ן���×�z%4�T�ђ�|�zK���h���u��3qP�9��:�Z1+��(�_N��=�|;�V</�V�-�|o���ß�u(���[S��c��nt�V�Cr��ˁH�	+�u�I�U�𻐁�eR�W�3S��k��Z�,1�1�6Q�@���hK٢�ա=}LJ�O�f}@_�M��
��;@UE�en_fM	V�gi������"�Z�׶t�1)֡�=�7�Xk:F�(X�������G΅��^;�:"^����~��e���qne" #\����O��7v5�;>���"B�<�Y���{dͯ�O�(����H�#;ݴ�U��m����7�O�E1�}��7%h�(�����4����G��\,�\qn���Px�7 �0/j)h�E�����,��H[���)��o!��$z�f�Sq�@����[Sn~iD֩v� �P8��C�}�y�\�$E��R�I��Q����xjIm���Y��_q$�;�zb��=���ԕ�&�cZ�U9Z��b�N�P'-~�n�g���*㢂"�K��K*r��d���!��)}�^�ݖc�
lJz<��f��e��A����Jv	��\��M����e��	11��# nM��{�]	p �!b��m{5�FqB��ԟ��cA1ي��J��%��3�~2�ñ���8v! %Ņ��_T1�^3Qk�A�]��Q��t �Y��)I�����_�0ɯ��Uf���՝�?Qd/B�����ײg��A�J��gXb#NRZ����-�'�n����;��ۈ�!y�U�Z%��uJ^� ЮG�L�K��5$�R���Knb��=,]K{�y��r�~����f͝G�ܮ?Ձ>�PY�7�H�eY��ϽREL�G~=s�f�
�i��UD$���0%�pc��&�ܿ���!�?�U]z�Mu�`�x��h`�c�8�A�QM/�w�.e��H��wp���9ݰ��1�Qw_Ϟ- ���:�k똤]�P�4hj�8���HV�#�WjX�@�sr)�;*6?�����^zy����m��:?z������Km����~�-�ˬ��*zf� ���VKUf�$�r���s�������@ZHC��aU�Z��0T1�O���T;:b�	��j�iQ�����ګT�d��>*�u���D���9]��A����\L�O�_�� ���J݂��� �6���5iOהe��|������b�fxh���_Eba#��0�����y���A`�mpw��5w)��$"ű��iM���.�M'凜����c`f1���x��&N�}m|vv�~�
�@��8�ˆ:9K���S�X1F�ΥWyr��Ѣ�D�d�YV�b�{REr�����>�>pq��
��Ճ��/V 5�z:l�X_�r'e��Y�`jX����[-|���#@���B�R�`D0�0�_L5�W��I�r �]G�+��{�0�Sc㷵Խ7�|�Xo;Lk���Z��'�ܺ2�5cZ�^�˥,ll煯�����>�q*����jR�%���n}� ����G^�	E�`����pC������=�~��Xǁ���ˑ�]���3��*���MPT�ܘ��ҡ?���Х�j��k�-xF����/)��D�K�o�n�.Z!����p��ߌ�z�D��y�5��]B=un9��Ls��z�(7�\�v���P���&�8�U��9����a�|\_��4�Z����?�L;~�>�d6�$�ݭd#�Q�k�X�{O��o�\(/{��t�D݇m��A9V��D��0T�ޮ$��x/P���-z��̪����w��0i����Q��u��oFAf�����'��l�jC���OM��8��N��))mY+*rk��{{˜"���QP���(�?���H:ְ�~h�KnT9��I&�0q�L��V�2�T�㧟Oh��Ԇ^4��6�Ā���.��ȕI3`�GU�xW�^*䣦\��l!��@)OPXp�GT���Z�k|��N�B�H`x�l�EM��-ƫ�R���d��:	4���y�2D�L�o2k'�q�y����:��GC=�$���l���~����0�x%���H�#��y�,�֚����{�+y`�P�s=8�Uț�H�$�۱, ���.�cu�>�a�{ ,��n�఑��>����(d�Ľ�Ɗ����6�swXO��k��D%�c0������y�8���*��r��l0ɭ/��4�f�n
�k1��ڄA�b� nUJmtzô���������ܲ�J�9InHʥ���2E��ZA�:}[d��,0:�ߪ�uu�y=��Cþ�F
�:d쫮�Q��3�`f'�B��TV?D�
:ʩ(��t�%V����ϛ�L�H��l����۟ 0�����S,��������8��Z��'8���p�xf��}@K����x��
[�Ø�6wB43q�7�Yη�iZ�����E�{K��� s�V�P�^c���Ƣ�^�X�#ctئ�ˠ� �os9>�6`W/�|_�^H1}ڋb;�&����|��fQ�&��?,� ^_˩�#!���'�W}O4D���@�����[^
$WL�g|rl��h�����9�L΃�y�Dx1���	Ϧ��Ƶ5�h�+ }�����i@-:�O��t(���U���V��L*��,�L[Q���R� ���<ʚj�.k�)���/�j�f�	.�|#U�N*�Eq��7�ܫ�RK8L|���rN�y�)Q�	i�b��tw�[�U������>���?x���*ʪ0�������f���3j��}�\"���G_k��u�E�r��]jJ�+�u�)\4>ұb!7F�r�D&-�㡙i~3�I6�b�5c����LoD�2ɪ�D��&��-�^D�>�W�K3r�͘�������a��m(�?l��jVl�~߸��C��ӄQ�kR)P3��?��o��1��]b�N(W'�Q�֭9iB?x}���XS,j��(��x�3�:)`�2=bkm���d�Dw�E=��{�(��jT�P��Kl��y\���I�f�)�#��S	����\Aڟ��5��N^^�^{�8�\I�\l�_�pʈ��N����,�Y�!�!I ߛŤ��Nȼ*&Ѡ
�A� L>�%�����gB�����&ō����\�9n���#�d�_4��Nq������ǲ�u����-�N+����i����Y%Ξ�3���c�x�W�֌��uSl��e*��z~��U���LA��/��~f�UɘM�k��۰�'�l�uA>Y"�X���nM��i|I���R��*��S4����`ly�!�*���Z]5�a�la}s�2^8�(�P��ZDz/� HM3t	}K(��K��j�Ms.���X���
�ȱg�O�#ѴF�jU
�)��R	�<�A��MR_�t�:�}U���k��4w]�h�mW݅�*�j���]�6�qy����s\��)h�o��Z��󃂾\��$��$��>�o���@���0;����g�V!�Ӕ���qt� ��.[���E��F�!�I":�n�&˙�i�>��]�C�I�Gk
�#玘-l���N������!���5�F�;%WO5>bmL�v�m�z��%��"7���S���,Ğ������q{�'�Km;��;脮���V�FA�z��O�BJ�kX�z�������&ru��ߖ)7"��s��rq� ����NW͍!����/x���"�^��aR����Ú�?3��n9��9�t8P�gȬ/N�0ت���i��ɹ�:1I�C�:X�2ѿ��G:T���4p������O�{��Q��b2��n>7�x�\��9e�����[D<j,+��e, Ԟ'�%�$8�+F
�BW؈�	HK�W^��Ӊfa_g&Sի��6��W�:�# 	BS(B���g����7�2��xs 2���} ��e�)�/K1�*aH-��8��V�F��I�:7DSKSi��㱘��;��v<}'$~��U���I=Tԡd�����z�K��#��gP��vb^�w��T��6�#_ew剋�r'l]�SvT� �u��"�0�'p��{>�<���z�/��L~5�M�4l0�&�Q��XC���?9G)Y��]	�K�/�xUe+�+���V������^!�'wH{R=b݈�����>p���Kgb[��j���Ϗ��w��ԕc]�A<�<��+�[�����K���B��G��[6��g|M� vhT�K�0^���H�������[.��O&nO���ȁT��]I3�"���8WE���(��3ֱ�i�Vd��qv�/K]��SG��^�<�#.@�
��-��=����=%���C�q�r1��)��V�f)�u�p��ʉO]���͐��bK�Q����@[}=KF$��Ej�
���ZS0�bf�c(���y���T��*m?����,c��m��_��o������AZ�/���wB�G�p��j<��'���`:܋anr�<�I���j��L��D�VوZ�w�t�	��ޗT�r��]�?}�� �'Fƪ�\I�&M��OF��8��%��K��R4y�=�	쇈�?���d<FQl'�]����Su��hav��_A;��$H��,��~�x�_	�h�P8��W�p�"r�hMY�	.����lm�)�^I`�E�E(���h��W)C�G$���wVv�X6���w���6Ijz�euNx�;"E�����
uj��|�n������i{�7^�ε���1+Kh�
�|��ٿ3������a2����z�gLE^�n�����E��>N��@2��ku`߇?������q�H��fp�_�/2�x>���:[�I�r����U���75�+����녳�cˎ�o��g $�DЉp=-!>�q�Q�����Z��A�I������q��S��	��v6;+�V;wZƘ�{62����o��o�\��)�SU*J~�P�'�����+'�"ݭς4�;���g�Gk��*:Eq��M��a²�䀳!��L��)a�s�#���f�|�s�*���\��I�]��K����Q���Wf�J�x�J�Q���
}�Q� �N�q5vT���v�����'��;AR�W9�I����I]����m~6�*x/�&w��T���x7���iص��*�*�"|��g�=��쭝J�hڣ��H�P�N^����֟�%+�tQd��)��Xٔq�䮦/��%�<#��H�ye`�)���o�(V�&)G�5/ەĩ�u`��c�.`�Z�ۥx�;�4��ړ㬱������Ҭ!�Dě�H�C���md���wn��7�R�)�����9���u*��qQ x���A�&��h%�ES4�w�j���?ܡ�y��f�aP`V�HVXល�ԯ@Tb�y.�Ҵ�y2:��;71����H��L��)�k)�z�"F)sߧ���Z�M��s[b~|�J-o�2���2���[��X��Z��Pz�o';$*K�Rt]�un���|%ؕ�V1p0q*1A?�P���M�r���Ӏ ��UЁ]W��X�{�'\}����@Ŗ�'|u�v<��塺kSK����%�ä.7���2`������	�:p;�u����&�|�{ 5,�RY����c7N�"?�щ�`a��qw�^�^��݄Y#�=�0�������7���b�J%�R�_j�՜:yL���u[S0!�Sn�����xu�Q��L�f�Q����/y�/�*���B��r�Ru�3�prBr�PJH~��$��c�� �zt���k]�&��q�+���@[vܖ1pK��f��P�fo�k�~-��іq�t0�J�=P��|I��5s�j�5��.&�V��]��,!m��|�*n�����x5����rc��vNk�!؛.]{!�����G�2����!�����X^F�y�n]�U����� �M[x��qM"��k�5��GG"����k�r�[�1��G��s��/2 D�����
E�ʸ��'vo4(3~2�J]Ő�8��5�!���(P�Վ�&�
���	���2���8p)�$�<&'�c��P��ϩZ���w-���|�m�ɂ�<�9b�g2��@jR��r����<w��ŗ�w�� �����&(�-EDs�|p7���@7����TA�\���d!�~�ۇu�6�����|Gk�f�ob���(Z��O'����샴������_)�am�?x1����),�W�n��]���mw��o�#ل�|�Wy8�}-�@��z",_�xmx<��� ��3���6��D�M;�^��G��<�A?�/d(L�n�����J�̠��J��K�;��������iJ�Q^�4���D�f�D����E/Z2�j�~׌\���F�۪��C�|��JB��������j{���?��C��G4���*.ĩ�4�"DCЎ\ҬtLgE%���2ދ�ąsu~5|h/�йȢ���mh=��%����S�/��z�n�b�<BĜ�W�f�>Mb�u�� �d_C�i�w ��BD�����sr;�`�@�g3��G8��rw��(Ð�Y�B��#�4}�!�̽pǫ�;�'`^�	hnͲ&^G�k;�;R�zٽv�7{:wP�T#ɭ���V[�����}⎶���������L:���ˈd�!f����
�˅xa�G�0z=���Ї$���Ϳ-�'�ņ�9�?��1��08Zəu�E�Z|���ls860p�F]�8j��@��������B�u��h�Y=���9/X%+�3�T�:5�Y�7Z������@��{����\�,	�q)�c-���֡\�c�E�2��q��[��G��}"�ᜂ�&!��1S��߂�A�3?�,��vۥ?�H'Y��:���#�B�:]�����f�X�����K/fIYɝ��pP���3E����&-�� ��3ǔ�;S�2��W���.ߪJ�5u����ʢ���wRAu�.��7B�cҋ5bوSr��#wn�{3H!�dK��ѿ>Kr�"*DI
�呡D��,J	O/��_t�����Y�� .4���
�Xω �99E�Q���gۏi��;%��1&/E��s� j����s�7
1<M�n7��C��o��\���SZ�J7d<��n��������9�����{�+�eYä�+��+ 4%k�#�'?w6>{>�޽K�ͱ�P��U�gJƩ�?�ػ��Y�>�e[����^=���"�&=�E�PR���︾� r�ӘHr�D���|%p���;�}
�����[�Z+�����7�R�3�3���pO�4�|>��+�,R��5�^��B@����8��?&������]�%�otǍM���%���~��*�f��)����JԶ�#hn�)6M/Ό����p����2���#
|�H�����+�����r���v� �EWi��hg�ɇ�uC/��o=7���Cș��%Tm�ֆ+���dO�FՂ�(!ɻ~D�Գ$��v9s���9�Z�~�&��O�1�0�!Y�|�[e���G����,��VR~#�8�f���N� ���>V� J��5���|j�j��L2n���ZC�Rw$dB��,�5�����mi���V#O�ꮪu4����])ܙ7����p5]$�S�c�b��t�Q<�}�c�אQ�+���^��.c��(9�Y֑nu'�;<r��Nʁ~��s3;PR��.K��<\�I���[�2�y�2�uL��]ڂ�xƨҰK�&asL��Q�����X���g$��?��"��(,*+�7д��ذU�1�`����H�I�F�<p8,Tg�����F������}/
�^��܈���^�>:����Pz�����ƣ3!�%���(K�H��+��It�´��x]���������8�@g��d�����6�ŕN��R�e���?��:�:�F/=v��z�[�Gwū�\���Wd�~������f��՚��]�����1S��y��o��a))$?�P����0�\q��KC��u�J�&H8�m#�C�ym�p
n��)��=�w0ay2x���"FVCSW�F.68H�&�`�U'��ģ����lZa�����)�0Zy�U�Z�괽��� ��|�M��B�����3e�K���A��p|� ��_iG�kC.���7���dU���L��ڊŋ�~"S��!#�c�KA+悴u=��5�S�A���^#��@�~K�h:����Br�
�J�W�dp�{�ќ��e9\%��m�625�f�Q�䷀|��e'
;S�{��e�H���Msi��8+D�[N��ӓR��(��P��g��l�\����^�'�-����VI����M E�!$���&�G��t����L3���ƶ
q��!�x��W�j"	����|Ee[�SGZk)@N���'�C�5g嶐+��J��#_��6�6�7�o;Tb3Ϫ�Dv�hZ�(_p�컑.-�#�`�H`���r/y�}<hfvm�~�������d��cl�`�]d�~%pEX>�)�����$v�ދ|ˤ��:��.��ڼ��~&������Ф�jb��i;�H��-����r܀�ʜt��D>7��8�J�!�i��Em��x��M�O=�\��U�6(�?M+���G�&~f�~ȭ\��������Vhf��_�5 �I�l�:���C�5U��O�C�2�&(�A�A޴8j���6��U �eggyr�+�(7�K�T��ޫ�?�"y�,AK�)`��� � ����O�3�\��2�3K���9~ (��č?`z��E�$�v��463����H�sC|����
lY
Si�&��ș��QR�JD��PM�&Yi�Y"�'���
��	��Yd�K����z[c|I�f����ӔF���;��%�K(�C�gϊ����:�P4Oq�A�NK�L�|y����3I�?���X��<�N"�Pvi��&�����pm������w�=]ZF��aε�m�:�L�T��7T-oh�[����m�6%�TJ?�����u��F���m}8粃�fp�H�:��1�{lK��_��	���ʕ2�ݨ�{���}S�uO�y�� ��4ϫ��X�#OU��	�Fy��CSO�<k�0<)��d��G��#�le�+���.�l2���#'��uZ����D'�Ju�17�娿�d����ƴ��'���!��s��]�Qߵ�H��*��geXmCDK[nvi�����u�a~q���{I(;jy(m�a�%�F�e��|�B���o�P���4@��#���-	�ž{������O]�5����~�`@��� t�r���GA��A
]o�K�Y��x�U�rT�v��"�>s#�Ԧ%*���8ˋ�p�u�$/?
o0�k�:�3J�d �X_rE0�?���Y�l����]
�\Km�
��n��Ǽ�Y3H۰�V\
 ����K��w]T��*�(������EV�B�,|S��>�:�G�5{�y�S��Dw�:MA�E.�I�y�=G��l�kGy�F�}/��;s��t,Yz3tx`��[U�ב�x��,X�vB/.��c���J�-A����M`�p2�IW4V���7�a�:�p�Rn�5��.�٘�.��L���39Y���b^oh)�B!QO�Fb�������@���0U$�<{��ĥ���Ͱ�$e�����aKM����N&e2+�r^����	����Q}9���Q���+>�$-������0]Ll�v#�hr<Њ�k��-://}�~�O��fC�ۯ[�2��P��_����aF�/���P�ɜm���9r�E4�p����;l��2��֫|㊅	�:�O�<�!Y�k�@�H[��ur�����C �H��/�M�Wp��U2�Q�0m�ʈe��0H,[5?ld]�>N��͞E;O�:�N�ȣ�0��9f�c�E���}�,�?GXuT�����&�}/Ʋ�	��4x�����ʻ�]���3��� �a!a:?�\bc���f�(^�����(�;��k�~��I��@{WH�y_{�x��ueˑh����NW�.���>Er�v�t�4ٽX�fM�����[oJ<U��u١0ݬ~4�W��ߦ���b�����Jx.�zO��Ē���<���!�i@)�#{�N�<�D>�"6tc`|zz�{������%Q�:z�d�1�gg��?iX�vK1��~�r(5vLO��	������e�~�I�5�	��H0��N��D*����H�hR]�ӟ�iQ��!Fe�h,d6�/񣩸\>w�c{o��@�
I�G�������A#J�{��WNP���o���<�U)O�U���\9ty��(Z�M�#�5��q.h���[7� ���%Z�ݧ�H����o�.�� n+]�X-���5?B��$^��eHP�Th����6'�h��Ƞ�XXmٝ�*Gb���g��8��s��I�L���NL9f��r=�J2�yn.����Y�t%��{8 v��8iQq5��F,���B$��y��[�>>��V<�e�}������^��j�("_� }�K��ɞ�U����o�5��%L��dq+d%V�AܙѲؓ�����V�����k��d��.vF	:t򧶣�y7�Zc8�����ް�ם=��	md;��we���E���sKt���G@�V�
=���@���q�K��"*D�t*^Ow�شe^Wt �6�2�o��ͱ�O;�L�3n�T-���e5�T��#����Z�z7+�"I(_����G��d�Ϛ�΀2�j@�[��A8?���y'p%�rE���/�}7��Eq��ʁZ�?~�{�e��H=�
O2�tu�<�������ϧN߃�}����&�����k���ᅖDt�
�n��I�R.�6;�r����U�>3�C��ǭz�Q�w	z��@�I#\B��%�|y��г8�9�5��
A�oq܎*��T[���=@�PIu,��d�}> ��������o NrrMe� �q�d#�{ڈ�j?d���CwR�7�i�f9����±N�/��nJ���ל�T���r�Q�JF5��\>��D�I��o�m/��;s���7�c��Xk�qQ�=�Q������dZ�4���\q�/�ľ�ܭ ���ϪO�����l��>�7�d3.w�Yt���_�Hf��O\�����C_4����PM�N�1� ��a>�k|~�~��	�������7Vi�b�ק_���[�V�T��Kv=.�x���A�V0�- �[�3��< bHr���.���xK�_�����:��+Nu`MH�������Q-��p����#��X��kc�c���<k�Aq�����Ⱦ�(��>���!x�JJ�������i3�(��4y�?���~�u����<����F+l�J}�+ZOE3�a�X�n�G�%�^�Z���{�ɹ�a�b�PV��q����x��kO�,>TΚ�C��Sf;R����xkq�%9D\'h癎��_�zw\� �ML�`�'Ѝ��X'�	$���c�ܩ@+��x�z|����?|�+2kY�t��#�j�ȧR�ޛ��~����˷8��۔^۴�}v��!A��NG�Ê�f,�����K���n������u�zl泺8o6�V!�_gUI(��Sg�����t�*%xh 1���̴i����n���g�#��wG<K��
&���	*�	�� /m��m4_c��ndbQ��Z��F�	�*e۸�:��'���T��&��'�P���>�b����2���3�?RH��ܷ�8��+�ٻ?Y~֧��(E�n+8B"J�b�g���\���	!0��*J��D��?����8��-9�V�e��mR&9U�J��!+2]�a�k�
,��*�Y&J��򿀹m�٦�����2?�(\g2���ѠP+N�a(AfqG�����0� �G���Ҁ$W�7��a�ꛦ���i����iW��wU���?W��/�T�g�ċ�9I`��bl��
6�R�O1�"N�S�5��-D����%7�c�`�Lw���骚���%	�"�$�caP�{`$��H��h1'�oz�˼5�5镯�z@�|K�Z��v1��rr��Ty;�@}�謊�E�ݞ#k�s��xZ�C�T$B��d�M6���)���e7(�`��=s<�����䊸ay�'5�mFF��ކ}]�>���������B�4�n���Fsw�_����;J"����##eN�R��Vr��3�<�<k��󇚊a:�Wص��Xiv8��iJ�4�^�9���$��0Y����A����Uɇ�����a�1Ig�ǰI�z�9�a��S"��y�����(u�7�|�.]p�k� ��iؔ�����z��0��
h����{tYW�u���:
�+�-�oyϯk�+:ۮ��d/|W^V��o��7�z�IM� ���C�CN��F��iV
|�y:�m�?�a���I\�3/��xV��Q�q�`ytI�9+���Pyv�f�AQ�P���"�BB���j׿�,WR�g��0�j�sVx �D���� �;��S{��ـS���x�R�Ƕi�w�_m�^�������h7f
��5�a�"ͥ�J3'?RԵN*��q���1{���%>��R�L�L�]��雩������!��8�3L�ۯQ ����6��;�+Cǭ�jۖv_-kg�5�f��].��^�m�����FϷ��%���ts���;�:�эE�'8�4k�lkF������ |&z��O�>x�c��2����g�?0!O{o�)�>Z+Pbr�LGG��K�:�q*;ո��v~?�('�q��B,͟|
cJj5��3�,�ordT�ҹ;�(U\ԭ�ss,��4R
[x�-l`�� `��Z�[Dru	�& kq{����kH<�1�@����+�ժ�gw�$�/�beDr-�j��ϨX��,�أ��%���B���u�@��Ӓ��&���C>��&vw}/�͹ÿ��-n�S�ضШg29��N��=�\��+����Ѝ���-" �M�{Nq�9�}�*�� U8��,ff�vb�=�8�[N�-��w���Q�Еk���<�jRDdX��p�ׇdK��D��(Kd��a⻆��헬���A�.@�bE �W��/0B}�e�-^��סlC�
�w�~O��oy\�@��X�!��.����6X1c5�h�d�$��H[	��{��^5�iZ$��ċ�j����i�$��"������?ar9�ѧ� +���+�V҂3�ʾ�\�N�H|�u�*<�Ɋ�&�&m�Z�v�ɍ��� �U��-�SY ��c�g���4)�W~�aB�By����є���� ��T�����~�P�A�ꈋPd��.4���s���a�D¹7]��|~N���e~��1�М
ڌ*�j���J.�i��5�|L*��g�|_W?w�ԩv"7� T�W�7��^����J@5?�98^I�찃�M�S
�����E}�bc@�3�Ӂ��&���6�ɳBڗ�Q]�1#4�LF�vP�_T��d���7��:�j9�W��-�૳�Nʹ �{y�����L��z4���qI<�r�q�}C�W7�گT~8�dLr��W& �8��!�NX�0��Q�_���T�_�
�d�|�3�.�T8�e�з~`^16h��&,,�b�������F����ׄ�Ξ�H<��=��_�� ���cܴ��D��H�c��Ct/?r���Z1�L)ʑ2���m,5�����Q�7gŃ��R�vh��	�'!h�'���gq g���gJ`H��}M �AĪ��.���|_��Uy�)�� Ч?��6��!C���4-9Vb9�ͦx#Ҫ@[l��JӒ�=���CZA��j�C�/H�]ɡ�XyMo�����_�����j��\�����A��F�"A�P��|��e�����}�ұ��ƂA�@
�*��9`�l0Ә�	8����]����*��;����i>0�C��Ի� �3��"s�X�oz��+��U9J������+�tO���)�b`4�Gi����l��\)f-��֍s����?R�{:Le�R��}�^?�/5Wm���_�:�]e"��yt��0������4�l>�u�����"�m���W��g�n+��'��]p��8��q�+�QH�%X#������#%=�5���o�@/�˔lT�2<�3�uJ�H�H��G����Zr.i��:����y1�w�2;�h�z���Ϲ����B���|�5�����A½�o U���c��v�eR�{��� ��	�W�aD�k�X�oKz���a�팈��;���&Z�J$;x����8�\�'���|F�S�~q͎���`����M��ѕ4��c_���	
�zL?3�o�X�(ZS3Tg�R��^�
�#�#��m����4�#�P�o�$���#�f��p��w�ʹ��/i�@�x�_6�厣����:�(����?<xK ��Mo�^5�d�e��[�������}��7\��0�N��۪^9�����<�IϨʃ�=|tN'Q�>�F�.��l2 �j��,uأ���R��_9��΂��[I�]�j�W@�X��L�����4����|r(A��40��V~ާ���tH��_�P�j�9�jH~΁���h���̓*���
�ks*N�BFp�/����r���Kj�'d��*L�W�������9Cħrz6���}�y��Rls�i˺,s��a��qT�J��4��ҵ�<�2�ܦ��7��`E���Ȟ�'EP��{��)̳8���WQWe����H��;L	�M
vȧ���Ong�jc��}���D�����m�G���g��s�91�2C�<��<코6��64w�\��^���8���C�%\�&�MI��'3�z� #�̪�7��bk����"ς�T�&9��r����ɤ�g���q�}zc�g�U2K�ejw��:!NI+i��\0/\곞�R_�M��T�w�gg�����ˑP�
k�W��3h]�9� �2Sk&I����79���3��z��6�0}�po��Ǝ��}����o�[HG�d��+���oޒ�=�M
��0��Xz�T��_VO��m;Q�*M���\�lE�{E~�~,xIe^�[?}l�e���ִE��y��c�!��.}�] `�{ƭ������GM��!ѣ��~6�(i;o#rC�2��Oc��������w߷a1@nY��z����*�J5��"u�p���I/��Q�0�P�C9��b���[���]�$k���iXj��罅���%�vjX��>D�X���F�.����P�B-����T؃�.1��v����:��C­�sދ-Q��"���=��b�y�03X����JE0�*�iү����o�ڤ�\B���QI,���%.���zf�'�Y-z�V�P�P��*����j�!�n&w���vQ� (rڄ� ���.D�aF�C���x-�~�`k��mB{ !�P�Ȟ~�//W���{n�c�8�� ���_e��� ��Ga�o���R���A��u����fU"��X�@���Qܣ9P^*S����<�v�5�O�EM���B�;$D���w!�tH&�!��8A����;��ay���@5��0Z�����)rHZ�����v_�e�4M�9�$䬷&w���O�z]>�îq��Mb���޲�S�Y[.DVK�o��s�7�;�� M�$�ۛ���N%.��� �����dl��33�3Y�
�
�� <�M�)V]�	��ρ*�Rf5z�h�,h����&RqٯyX'��@���p�f->|악-�æ8���і�h3|�Uᣯ���1sL�7�}��z�&?��HmDY�$y�fL�ݗIJH�V8���w��.�D���T��-e����Z��R
0|BT΋���Xg���%6���@��'-R`���Uu]�~�`�M!�M��{$��f�����B0ɹ]`�B�(����\ص��E4��l�>� `���,E^�b�P\��JtC�\-[�׳�u^i���X�7�H?�$TP�Om7Ė$
Ss܉�V��5�s�R�W=k;�V�f����ШM����򮅹��-�U=�5�S2D}��D�C��c����쯎��Y��3��xw�4��Ze�QW�V^����7��6n�bӰ\|H|"�"�U�^��-���p�8��W��H��<�^���C�3MNI,���)�~o�-�v���Cٌs�<B�K��@ICD�n�Di+�s�����)��B���b��dO�j���\P.{�L�ڝdr�N�7��Y����]s`=x�֛+�Gj�
8�'��Ă�C�����M�S����w��3	��ؼ����]��� ��O�����|+��>�����C�k�d[�o�l�G���]6��L7|=��g���<\Ϋ!w<8�n�VZ��!-��Ǣ�Y�*�>'k�L���O����N5�qjQ ��:9+���Z�WH��u4}��y�W���dg��*�T���51PgC��8�1-�%
fi�>�˾ԂJ��9�� ֆ���LB[�v�[1a?�%H�%�U�������M�����@gA�(��&.���1�VD� $�仍�O6�����0e��4��y���G�r/���\.�w�vB���<������y#~ʨSN�c"<n*��&��n���}M2:���>+;�m��؅�tǇ�
��x�0��5��3A�	7�Ǥ�� ��t��*B]��ްf�P�����s�s��B����'E_���ZĈ4D����-jo�~�Yb� �C;�d�v>!��n�vAɹW���
52�@^p��*1��t �d���,�{Zܭ�N
���q_V�ȍ��&�,F�=�Ķ|�=��l�ү=���`�j��T�`WG :��Z�1�����h�3H`�g�kQ��I��Z]�_TL�{�Ba��'.=��E�vb�$�`Xx�4ON�\W�<�����X?C{�f�@�xL�hn�>��
��0�&�L��������z�]��Y��;n�ϭ�L'��R@8������JpF]�-��O�x�ǘ�QGeB�4�(K�;���P�-u��B+x)4-�{nfEU)��p��PW8]%�������	����h#j��  gśT��4��QM� �X!���hA1x��-S��e= cＮ~��bz�b�E�m���È�7�)���B5����P�Y.�
�L�UR��f�J��G���I�u����̐8Ʌx����@K�^���v��S���A�J~�m�ҿ�Ɯ�ډ�lX���T��o�u�Xe�*��0Pe�/ ��蹀gkә��O~&s����=t�[ ��l� nm�7�K���}�14�9f��?
Ȗ�~�Z,�J�G��59z���L���kE�~�ew�7s�s�!��$Fs��=O���lH���V�}��u4^�#�&}[�$�S�l��
���P�x}�Ե�&v��&�|���u��F
tѿ�a�:�S��B�d�i5T��F_�$�wE�ycd�,~�P$=}_4B���u{w��.b:��"jC�M{Iy KvL�j�����ow}�t�Hc�Z%R,s��w<u �<G-��	��q�An�3~g��hƃݹa����Op�˿^2U�k�9�1ŐM!����D_ީ�pYՂՌ���( ^��0��Q�s8j��u{<)�X�&�z��yA����ؠ�	�agW�Ǯ��8C(�

�Xϙ¯���r��\S���(�;Ij��O�-���z���)p���I����m�q?�(?��D�Q�3�v�\����2K��
"���!	�2:-��4�r�-�iS�\���mY$�R�ָ�9��TW�1�'!3��~4�f|Ž�Zy�L��ő+���W��v��S:C��m�(��0�E
$��C<�G\�tݓ�l`���ߎ�S�.Y���(K���GKP_e��L�,�ܹ4���k�	��
�K����z-%[�h��^�A7|��/#3�|�MՉ|� gj��*�ģ���l'/��_��;�h�_'����;����v(��2����^w{�'o�0��� ��}*P8�K�iә��\�Y�CH�E�]>���&�u��?Y(��{���N5��F��V��X���5x����듁��-��*��ʌ����{@'5LZ��ö8v��M�Xe���2��y��#�ૂU{�|YjP:X��o���u�+&��N���UK�>���� �����S|�i�<���]��p���t���D��=g���� VI�� ��R����P� X�+B��Җ�I����8��>�y|9�ۄ�i'��zGa0�:s�I
7[�`gk��a-Z~iS�$ �NA�yS����X[�+��!�[���A2�-�mˌl��v�Qk~� �LŊ|��ET!^��no���<�`7�����T0�{��Z3�u2�4�F,�TqFs�Ɯ�A �����Z1��i�j4RDf�;ua5�!���4�l�|���*94� �����'��S�7�����0�ו����� ��O&������Q�����v�s�<�з�M�����ݩ�N.��=��h���'��ضnV*�册5S���(����yn��dKs>��F{�{�i*o�~��T�ҳ�K(��#QXt�Wn7��Q4jY�6c%�
���{R�?��G�須D��eI��{.ò'ҏ!8�p���hp*�.>莿��U�fD̦�Ӑ��,�l�)>�0�g|���Ȕ]ć�����/�y�
�Y	eI�p�Й��ޥd�:9�������ƺQlb���G ���f�~���<�c��C�C:Q[��s�%���s�-4!ů����$��N�1̮ '�'D�%��~ I8o1Ǣ�D�7��|��K�*�0��I��s��D�F<̬��s�יkC���+QOH�~�E��;�0��l�����AZ^F�_l]�2e&L�\ʾ��ԁ�JL��ghi���h��նΕ�'4c��Ŝ���,s�Vݦ) �j�\��;et�+�U��N���Lu�䉃��R� ]��0� "u��e]���İN�BD�T6�i<�^3�}���w�J|1�n��O����$4i�6×��z�s,���̫m0�{�'p٦��l��+*;eMDP�%�����&
\�\{�<�b gv5�T}���t_��[!j�� |�,a�G����q��]�Q���pb�d^��\ѐs�����_%�eE��|͂�4�0vMf���I�U���r�'-��ac�|�b:C?I��Z-�w�3�R�z�H�t��?��Ǉɡ����"X~MH���V&�}H%d$�y�^��� ;�LlK/+�[�^0"¹C�W6�B%��$�p;����������YĢ�y�>�X�P�c/�f�G�K�����Xq�sŅ\|1��w�Mn��Bai�uq��?H���eƧ���
Gg	���`�i<����sz+�FG��z���� I?��;߼�.�&;^6�E���F$��:T�Dg��5����A��P|�c��վ��Dv������ޥ���mH�E	;��^�J����`���S�^�@���(��c��je���z�8:���ʡR�(�L:�{�����I�.��	Т�K?k��V	���n�����	0V��+[H�H�DU.�� j����i,J���3=�� 2i��� 6]���y��s��nW�̛���-�G;�� ��%�pi����O�[^��'~�M��Ҏ���8���jL�^���
d���]�
Q�8����C��@N��'�~Zj�dp:kYzӶ'���ϵ�
�$`��OmU�'������d1���!0�b2�f���9hޤ��9��df���^Cv:�%-:�;����I�b����^��o�h�Q�sK�,,��v7�z/ Q>�r�?����hK�%u��Y_�Vy�]āt�iD6	��cE,�=�"B �(��R\��-c���FQk5� ��e���<fǁDj��C�MY}���&_�t!����x��*j�ݳ��F|�z��n*��a�8e�m�ˇ�L-)������#�F.�b�[ڛ|Jw[sx�Í�]��E���\�<��n��HP)� �.������$�:�_���c�ح��1��Ʉi�u�|^\���9��EL��w(Ծ�Y��_1�g>{��ɛǀ����Xi���%��	v_붿�E��h������9F�~�ߎe�1+��{��i���#��ǉ��BAhzٹ� B���-��ط�غ����C�\X��ۇm����U�T�� yl�d��������~� }��:��d8��cs�n0*�`C��};��P}�Y�3d5-���R��P��L�cWN�深�4k�
+���LOl��B��#�Vъ*����d[e�dDm��&U�ej��ė@C�8��z <�'�	ܓ|��O��h����N���o��/�>�F��nǥѣY�dt=$HP�������lH��P�s+5�1=^M��l�j�[P�=�'�)�q��]*��ʩM	�JTp�	�氯��Gg0 �4���0���֫iF��ue��=p�l����>�V�!�E�:�����Rݮ��geâ�
D��G�ᴶP�ȉ�w=��j��BP�g'%�q~�է�j}�Y���݁��bЉ��s����/���(�*�-O��m33��9��02g�^8z��T��i�6M�������Mʗ3�Y_�o[�@��_+��d����Ƽ�ҎDA|������2�mz�VL�p6�j��*jY��K=)+N�fˌ�9�& Uɻ�x��*n+j��0��}�Ûk��j%J@�W�4�SVW➒����Cu��y�A���Q(�ͺ�6�2�O�(�L�(ǁ�u8N�eI��bUx�9r�c��.�o𣮾��[�Ġp ߪ �d?����v�I�f��.3�� ����d (�&^�B\��$I�/�|�K���-SS�s���� �$�[�E�r9O-���1�cS�S������J2��X�v����~,�UR���n�bte����[>ʺ`0⁑�\}�'\Ck:����_�ͤ&&!񒉎9�q�&��63Zᙫ0rKW�e5f:	b��έ��k$٤9�%�x���a>&o�^�y&��l�mc��I������cU�J+B@�U��z�Do��T6� &żAyb�\Gj�V�!��E���xj�\���ݻ��θ� ��RBL.=T�k|r#�9�J���r�0�W��E	���2c�+��Q$ؕ���q��)��,7���VT���}1^���Nl1
H0;�H�z$E?a<-��﫤��ƒ%��(;�.����>"�� ���m�JI����2\ۨ$r$�2���UjY�=��LKC��'U׸]����]ݙ���K4.l�j�����Y����c�.<��Rq�a�Z/�˄������
���H��eDsp���[ �Լ̄9��,+�Vp8hh�H����g~�9L�Y��zN���w�2���t"�C�J줜��~k���ȡV<��1 y�����&E$�?91��㖃%
�`��lq蒑�g��K3� oΆ�̧UQ&���!7�N�x�,�4װ��,���� p6
ΗF�e���2�i�fŠ��5ȯP߽����$}��H����?���R���C��SWØ
:H���X�����9���L5N:l-��<(R����t=�WD�_^����D^���I����t�vVK~]����j�j᝝%� H�̻Ϲ��h���)2%+3�X)}��Da��D��.lC��ޖ.T�W��P. �Z�w��'M�h?
OHG�z��*��z����Qa�x�^��/B�)QD;��¬?��o0�Uf�����ck�&{U�=+�n�9,��s�Hc����U儃/�Jt�oVa�>�C�)��.�GZ� � �)��"�!U�bx�bj(,H��ȑ)�7�� W.�����`���K����F� S՚�!`�
�8���:�BQ�Y�;���ڀ.;��@��uɓ�[Ϥ�DZ�!b�.����`/ ���629D��`�U�ƕ¡�Ǌ��x�He
[(6>L T#�ا)�@��wnr:9fWos�8K&�B�nHP��{*��*���5Z��U!�VA.2����^�J������W����M��,'V)x�G��zYjb�ZM5��.���a�*�C�k��5�ԓ<"sP���wFFy6.�|�E
k�S�DSL&��V�z.�bA��+1�1"M�AD��;��4(�(��O��[g��MyΏ�[\��j�l#���?�� 1�.�O+�Rn�Ɖa�՘�/o��*�\75��Y�(�h��u���wq]�lpA��l|� ��0���G��B�w����B�ț�+�A��E��5w���¶X��S]�s�����,(stКO�p�G�~+�S�@�TN���u2-$��ޏ����3��&T��d+��nl�?<~�����j�8�x5�F�V����-:���7o�)�2�����zOܷ�Ӻ�51����n��n�
��լL.q>�搻�hn�r�r.fߪ�JL[��FbOr�h�T�'v��W�V�4�|~y�/��|���+6�yQ����k񴲄���,�;@m`�s��������B��a �"���(.0>��-J36���K��v�J�9��n�i�W�,�b�Dz���bk��S�"�J��x�;�;�R�S=TK��%po�uc)բ���g-��m�.7����a��q?�ŷ��>A��"CI]z��4f�Pe�}�c��eW�Nt�_x��.]q'^��9�ӌ���bdu��R|�}��l)���h7��2�8�=Zպ��<�c�9v��Ͼ�JZ�lv��f�k!D�}bPЦ�mw��מ��2�^F��N�c
X�N[H��|�E�#@K� g/Y��:��f�8YKrY���_M)�o�e5��@��c�?�f�+��a1x�}p���o�l�Y2s*���d��|�d�%�-�7�C�$��Z���Z`��`P�1Tr~���#8��>/{ُ9�V4�Lk}���LfY��S6�-�~��F���Q�����ߩ�	�𒖊A�$�qȋʠ&/���H�#ؙ� @4>�َI�,:>�p�H�8 ��Xa�A�&O�8#v�2��ޖ�$���y/��=�.�c�&���*���In���0��9w�1m�~L�c,��pv��.�09}\����h@�b��10�,D"��J��B�.�Q<c�d]��8"���C�Z�4Ү�P�����	=:�H���=�z5ps���$��W��1y��!%�x`
�?�ZO����~�*��*]vҷL5����<��?�� ��b,�;��>&�g^�G�����0g2�f�]��5S�'�<�/��8/�G�aH�3ɛ��;ަ<�o��\��P��'�Jyb��K@��5���wA|�����Ho�l8\����i!,����6��H�Q�����DE	}��ei�,�b�E�{G�Y�9�ٱ����Bw���M��d"@�I�4�!c���C$:�>��)>e<q�@�L��q1UXiO ����Y�ÃCw_���AEb�_���}���&���$���!�Ϋt�·ښ��$�8�܊��랞���>��M����S.�|�T��0����c��V��M�}��{&�s����ǒ������؉�T�`,������O��m�/["mt�ӓ�f�He�K��͌�x�3p>�'��$�6�r+�J�i��kbV��D�_�Wõ9�ߒ�}p�0�^Y2�f��z+*l�A�J��ʘ�;��^�#CzJ4	&u{�,L��-mx��]/^E��=A��r
����IuD+8���yC�m%}�r��3��O�!9W�x�b���Wzaa��^U���˲N������5���~��{uƓ���/.L��ͧά�~��"�ƽƼ����d����*�ĮQ�8mNE!oq~6����|�2���[�^>_Q��:��)���V��nc��@�@�(�Mz�]���W*pA�@<�?����F�����|)��v�Ȭ�����C	��G��]��H�ϩG�nT]m�aL	�
+}��'yD�뚮��R'�؟�%����h�;��?���b���~�� �X�@ߐ|c������#���<X(n�N�,�Lg�ڜ�B�E���x�Eʆ���u3�u�2�34k�NR�\�1� �
��9$�CM{����q
]4s�;Rzͭ,�ca��^���<_�ĸ��	è����C��)��w�R9��՞���W�W�J�ÖI�c��i���i���a$�<&D�%��!��J���L��!���~���pW�8��E�ET�~�_j�[��ʋ��9J4��۱Z�Wp�{%��.!T$&���w�tcQ�?�;�מ�:7�`+i�E���Xx� Fj��&�?��C�;9�#I���@6-��Y��dEHHl)�sf��X��*�!��C���2ZA��C�Q-*T�h<\�$0����!>���&�B���-p~5��=X�mĽ��T�GU�>�V�����h0֟�{��qS'�\qi����g�'��ZN��eT�4F3��8�Z���O@���(�u_%?E��mֿq�ʇ�3�����!��8�R�[�]����^;O�"�ag����Ȳ�KKfW�Lz���5��G�.��{@f��r�[��f���)��%����(y1Ð�K{��<��;3c��s�JU�%�������:L�1ʏDHz����o�z*�eczG��J��`��r=����S�Ɋ�m{ꥈ�c��oe��Z@x]i���41�OXf�9�r^T�Cr��R&ؕ���w���w��Hn�6�3���]D|?���A7J���; ��ۅ�5�����*����($[u�]���C�~��غK�y�}Q�'�B�����w��ͯ2��+���@����2e���b����;�Z�<&˼r��]����wn���1�^�Ĩ�I��q��Nu\=M�W��J[WxJG�[/F��l�ja�������w�M�gR�I&����ݤ����!8;�����C:�o��1��Ș�e�T	
+�WD��ƈ�Onz�M��	��R�7�tT)ْ�m��}e=�mO���&��]�`�J-�}Jkƣޜ@C]=<?�f�: �Y�V+k����v�6n���[�Ge/�n]W�W���#VL'�y�H*-��,��d	y+���9{�C���-D�����ˉGxùMʷײ:����l��뙁Vo3�]��{i�r��q�j�Ӭy-:�Hȸ�1�t>$4�S�,:�.	A���l�/����D��\�t��̝�vV~g�Dy�ފ�7p��]����
����֊�C��>3�eR�~���*cI^�u}���F���(���p��=	,L������b\�j��m��C~���z?[�|�~O+����B!�$�K��l#�N������>ȼ���9���	O��4{m�׳����7�0��������krF��� L�J!�a@�k��3V�������F��_���ə�=?��l�?j��y�h���l��"Qad����9D2I���TG�x�����w�)���������������cԼ��W[�_��3bk���TM� ��<ý�˘]��`��;x��3�3>kHL?$s���~Y��0�g����(�ǐ��|�ûvh�f�: u��p�%%^~���	��B�']J+$��n�R2#AlH�q�q6�Aos���;�蝑�2�E�@kt��8K�5P�@d��͗���C���5h�G�^G�
tU��CX�S[%��i�ȍυ�z-�]����A�<�W4��8��M�_� �L�E��>t=v+�14�GQd����\���Tl`�����!���IQ��z�*�����$�Z��c���\��"�Tlg�O�|ȩ�~C���R#�a�D�>�������ց@9:V���Wx�	1q92Gnp�������dG�i�n��Va����<��'�@��י��*��s[�<V�˒'x�������n��uxO<͗�z�#5��H�?�P�?��}������T��6�̸��c�$�up^�m68'�������B�-!Vg�b-���.
(
���{�m�����)��;">_�;�ҏ�`T��m@�OR���,��hR�ޙ�Σ�����3�(c� ��G�Dח�t0 �;�I�Q�U\�U	d{Y8�*A�������_��ck3��!vR�m��$�	ͽX�sy.p�˟ED>)@�^2NC��)��F=$�+@iUv%k��"���|�� +;�8� ��f ����P8�z�I��~'%_g�*ί�ީ��L�{�u5R�u%��i�ַ�}�̐��{��ݭ�,O�+�����V�!ID-P�4-�I"�d��Ћ�8%`�:�����I慝��f�����C���z25A�L!>{6��(NP	%k�Fg5�EƧmojg�sF����~��$�g�Q���8�`�3�K�J�c��>r�K#�&�5G�S��HԳ_��pc%^�1�8��
%k]���*�]>�C$TB��F�Dw�1�����E�`V@�YP�� Y3ʸ�FB��f����[INM.'�t|���d���Ld�)A����z!���2D$;W��p�A��P�ip�#X^���q#�.��G��&��!�9β��~�2����{�69�U$F�K�k���57��z��J����9�f��U��ڔ�pS���#u&j��L� ��[oF��2%��AL@q5�2��?���5�7M5���rV�vn ^���䉧F�{�����hY8exo�4 ��.�st]�ӊI�����2k�*z�Ɍ�k�ȺO$��x�S���FL2��M���g�����o�b��."���\��S�ۮ"в�[�&�9���kl�Q������*�r��Qx�z�rG�u�vWoT�Q�Ğ]�hT�I'���V�N#�f�񆫂x&ִ}���ȥ>�ٲ��M��U���e�����>O�h�����C��8'�*E.��uQ���˺tb���<q����m�_[@�f�ǵ�'����<�������%�	ɛ>=�(����k4<�+O��\B�"Xߵd��w|/�ot�"N�H�½`U�+�3kM�(ҷN�F�2Y�~�%=���Ƃ���+o��ޭ�+��#A=��%!���<�M)�B�=�(�]!�t�F��Sv�dD���N�Qg�m��G���kK�[Ez�PX(�1���Nn����TQ��E�B����䁘��=��(m�}�:��!}V I���j������-���c[�I�ԭ^��b�AW�܍L�-�F��t���,���eTxőxo�(��r[J.�W(_���a�����c�WM9��Q<8�0	�ț�����.��0�g_-r��KB���kԑ�fF|!p�o?�n��� ����Hj��X�uWp�(DͲ�u��ƿ��]��
�"�*ڨvd|3��[��>����Ӆ�osBEy����sa)[:�aj�d}�єn <��D�NUm�cVC�&�������D�9��xԭ(%�y���
�\
皬x�+��@Í	$x�e<>��>�Irv=BU���A�xo���Z�%/4�{�����#�x�B`z�\=�\��3��A^��j�d���'�m�w�/�lCP*�g4` �C+ee�qf�*>�S� l:z�{!*�A�`N�fV��u_l#��5�QQc���8#	����@�!(k�W�d�;a��b��/d&Ζ��O���C��+ԁp�7�_�������8�;��|!N�1Ю(�����ǀ�ɸx!�/zUmO�P�e�bI9���b�o�8����6M�O�:"z���fw���`�M�4�V���
��JM4������%���%������!wM��f��ʰ+=�V休���hc&>�d?�rX!D<��ݶ����2n8�UKExk��˴��� E+uN[�v�^ϊ� �)kj�Ǉ���N�8�P}5��_�@�����/��-!�"���dU�a�J�_Q���_�'��0!HC�"H�D)�C ���n���<9�) h
�0r��o��Jx�<8f�h�!׌>���=��b�ݺ1rn���Ep<"}K��zǎ�3�{���� ��qx��t�ưRwZ���AFI���0����J��-��F�mp��P��B�l�Q�#�b~�lZ��9�WK�'��%5�F_-zD�J��lK�F��1t�r���i�5�Vo���Z$�����-?yO��M�R#�[k��T�&��F<�)?5���4Ī�K��{B-��������enS��lj#5ս��9��=���j �������9��7��`R���!׺Jg���C�����9W�kIF��ϧ�3ީ�Z@��s��5�է�M�.H�b.]2� �].�tM��*�]C:L��5��r
 +��1]�tGoRQ�	Z��~�����>�=S�,��,�\�5�T�v�&�-0%:�[�ذ�i0a��4�ubAf�Q���fgm�(�)�p �J��[�LXN3�|��x�PA�Zx�э���M�N��g%e��<PwCQF�~���|�*���i����)�J�S;���J�i��g������,.I��$�!�Ckd�e���O�4����+�9.�h��kE���moo��q�?X�>7�H"ֺJ^�+�N����ps����N���Z��0Q�(U_�*j�S��>\k���E�bA!��1��U�W;Qf�������/�k�YP�)��)����n4��?<'�@�И<�K�����r{�EW�٧�UJ�A��0�ej26��Ёw	�!B��/��/��'4�ƾ��\�)���Au��<����B��j&eJw�g�.V����a	"����H_ֻ3*yУڅ�8S��F���Gk���N4t�02l5>�TT5c��R�.|�+4�EG3fs6��N֧^���lH#z�Y?�/|��!W���,ZE��s�g;����?���1�����#���W&�w9����#�31`���I|�8�;�8���N�� #�9 FS������U���m���Lѧ5�����#$�.*fH)�]Iė�A+���� |�#��`�� .0Q�f��(�����<t7F|��Çd:�d��H���0b�b]�QK�!��bCm,A-(h}�ݫ���_��d�/���BrK{J��*Z��{�MXʼ�@F��yD�lMR�t$�
6l��D�mj�?�n0�������B������%�y�,&�bP�JVQ�~oĿ*�O��g
�d��᪮;(z���@���3
���2@|n���J�7�a�Z(2w��:ϠN'B���P�a|*�G(]bҺ[e�������瞁�f4���7X�GytP�H����n��/���+ܳ�oɗ�y:*3(fiZo�����͆��s�TP�6��2r�Yj�e���m�?���P*���S��f��՛����!Aq���/3I�Kr!v�O܅%��ke��Ѱ�]����S�����q�_6�L����{��6������؜���!���J�v��!�pvn�[���5�1�:���*=~�Ͻ�3aT��0��ʼ�����p�\ѹ�ZU���,�� (���(��騌>�ti��g����в?�t�1�2���3Ax��R���Ǡ�D�N�+�M���(V�nUs�8����sA�F���|��+*Խ�4���!W�����i7�Y��j���	{���s��h�~�b���I=�{Ϯ�)���c�V,����C>��*���@�\5	���R3�`߰�����Y��M���U���p^)&`r}6��+�G�l:Y(����26��[�= @�#Fc?�ȴ���PШ�جH��	]�fGLVք�X�K�gߦ��Дi ���3�d��H�0~K�F_����|��E��c�"�fH��  �xt��jD��;{�X/�WN�o�ls���d�� (W�G{mVSm���t����B��]�B})���4�#:a��h����g�� }$?%�Ie��^<���@#y�`���g���I %JN�>R��*��2���!gM�9(0%�C'�1$�	%-T�/k�<��2B��]�o �����'-z�w94�sN 6d�n���y�ԟ���o� �%;|��Y/���g��A\!�`���rp�R��E9n_`BW� ���_��˯��%���s��^���������,�,˨^X,~�� ����k$���L?��+��u���H�&�=��JŐ�������*�� �M3�E"(��GqN7�!�������:�3}�l\+M�3>�b>��b��Gc���H�4L> ��� �&g���Ͻ���v�@�Y�[E����hc�m\��C���]�Zbē�]�%��) )�@��z҄<���G�Q�X5S��(ǻW���Q�뾶�jJ`��ݶ.��K��h��4p���W"lR�A'����C���w��&$H���ۗ��YW�&PQP�Nɯ.]}?8�%��U3o(:u��='�F0�E���
�A*�FQ��@m9跆�Hj=#�o��l�Z��p��6�l����dZL�q{��Lx̴_B���Oб�$�v�%��5QX�d�V�s�o�I�thޟ3��a���%*�_0�9��x��a���%4��+�@�����%��C�_yyn��e��������$M�gq��X���ڀ��_t��N�j�/~:ez�g?|�ɒkl�8`b�C�h�Z�?T ��@���VK��=�=b�t]��av��0W��Y����k��H�G\n��70��F�<+;h;ώ��+��b�qy5'�Û��N��KPa��է?�|��
"�Yf(I�]�W|t�?�3���4�P�A�}��w�D��k�wv��V�D8���w�20��W�e���r�<}1�y�����h���S7��{��\Sn)�B��^E�������0��'�'ʌ���[��0��XZ�������6��C�N�T�-V47@<�$����&��|&���H!�I�@�%�,�m���f?p�K�"~n�D�5!�ӈ����ϼj�~+3�ua��+8�6��k�v���bѵⷝg���e�2�*�K
���b;P��b��N�3cy���}���'TX�4������x��,i��U�u��A����=2���g8�b��-������m�_�?0�p��w���ɽ�DwJ����!�R�&�2��
�.*N���\�`rW;�^�8����K����uMn�����Qj�`p���u�yB���Tx�} �5����a1�?�kB,nQY�ީ��Q�^nsr���t�T�"���Y/��1T3��'9s��S	?���x��'��wZ/ߕ%:&�L���k�P2��y�'H�r��8��ި�٠�5cF��l�9AYc<����:"�;�5���������K�jؕ �