��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��ܼ��e߈SU���AR�>+�y$kgG����)!"���S-�e�%]�gf5Դ���s<G&�,H��gX�
܎­SH��76���kEb���Z,��O�\��X��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�s^W���0A}�����L e����EF^��ຬ�bՃ�-�O�,Ю��sZ�WF���])\�9�W��t�6d<�3S����ii��O��CalZT�S��Q�f��	�l������r�3��7�7���|3G}����e�Q��wy(�'�3�OF �I�mc�Z;R�?����ǟ/�r��@��	ɣqP4S��}��8M�wW��J ��.�o���&=C-hSF���CF���d �s~��]4R�ͩ=�olEON&��^6C��s(�?�,�r�z*��TR��V������;;��"/ƥ��8c8s�|m'5���D��@�t4�̚O�_S��لy�@�6`�6�k�:j�.�(������⧉Fn�q&����o���Az�X���X�oMe�����F��9��/�Z5)�z-'
���A	�s�f2'Va�T��0���u��e����xIb��!!�������s�/����y��������o�^�ݏ�0)�ѝ��S{A�9�%��Nvm����l��`��㋑:$d3E��?��
⦞�؞����X,,�t�H���"����џ��1�#��ᶛ�p�Q��.P�/�������q%@W� {�a^��g���OȻ���%[%�<'�+�If��m�I����J�b`����u���c0�ӕ�G=V����i����ת�Ƚ��(�9*�g{�x�b ���"�Jg�
�1�ae��f�t3�8;|kPc��ݵ��~�zj��5`�c�dU}=f���1�q�S����m��S�nf���W�1@m�Ǝ.iz��%��EbT��{�zi\�M3]ks^�4�;f����55Eaqi�E��e3%ѣ�-��I���Ԙ���L�O�<�VIgX
��J^��k�%�����9�?�\oI���'u����{Y���j���bۀ�$έ�
�����Z���	1� �����툈i!(�f����Q3�4
���K�� ��_1*T�\.L�?�H�: s��$I+v�r��S��S�[��l�J�+��w�\�a���	P����聭�nx�ކ�����A�O���t�;��Μo��*F`p�E�H����k��Tuݛ��x��L�ɽ�R��n�[*$�/���DU�t���BÆ��yG���|#k�8�\� i��;��:��]�gB�ƒ�:NU�ЉF���	�ODF2Z-�u��
�Ӭ��0=������=aZ��5�R��I��Y���<Gt[�ͽ���B��`��"`nW]�]6����Ք&<�S1��]��h ���g>yQ�˪�w�����*��Uݩ���T��
�`i�v�s��ɝ�y��R�
����18i����z:$~�����jD����o�UI�&I���u3j��0��[�=.w��C����2�u�Z��*�{E���5�z���ht�j��!~�0�N:�k���1���%ʵ˓���v�ԏB�s�e��=ڢ�%Ex���Xr,�K���w�eU@�^�3x�+e5�v.��s Q�S)Y%b��v�&��8IfIA�e�o��
�42$��M��z׌�w�躩��|�:5�:����zT̨��ủ��6�<�0�4��,
�L|k���M��,l�%��0�=��8�Z<��ϚE#��.��?<n]���Wj��69/ gM����y�����t�!y������HJg��`D�I
��l�d,1:���Á �ĕ����a�wP3x��v��2�˷:� �J�=���*�v��t!էm�d��� �u!N�6�WV�<õ� �8�?GQ!�if�b�]P]p���1�ʁP�uʧ �=�����6���>���@(�30��^o[n��.� �{���,�)��V�e�����#��v��\=�8}��r
e� ?YI��XBlAR�F$	Y�v�!w�BJ�c����v��,�ބ��Ξ7��U2�WD�օT����G�(Gx,�����L!`:�4(�h����j�='�;T�\�O�j�c{\6��4�5��t@0�;_��g�K���_�&�)��dS�R22�l0q��`����#t���x���'<P��C�\ц
}	M�u8���z�^�bt�I�]��Y`�zc��,I��x�ז�IT:l��3��.a�zĜL��9[���@��k�$��W��()������S�,d��RS�箅f�|:"pa��v���ac�F�,�1���LB�ۧ�.V��_y�yt
��U$�ʮs�]Ve��w&�d@Z@*��H��z6b���y@���y��bt`E��W�܇����b��O#W��/# )��rp68�T)a�[0��$g�ө� 0ֱ������` MU#��z��x���xq�ٶټ�d�j)����k�Ip�т�q>���n�˽�/#�P�|��C�ԉx�Y�S}��)�LER)od������=[���@�	��u�W���[L-b�.(��-@ q`�bl(q�J��B��"����.͕!u��N�Qo����W]&��2��v�3���w�	>9������a�x`D��Mz�׏v7�b��ڡ�!,���	�~Aw�"�N��8)��H�d=�1u�����lT���D�������n���p���~]��8F�h�b���|�/Ab�NM����<&�����SV�D��\�5D��4jE��E�g� ���i���^�7�G�9��x������:��j��԰��>��,>(xb64�*�+H�C+%�ep8N=W���a�F�<g��-hj%�G�`��g)būm��/�����43�����0�K��v�|Ǉo��/Awuɓ:3�ìEI��,�#��,��bt�4KD�q���-!+k�@�
���bmuR�̱�/gj���u3�^MDb��Ӭy'й��m�p	�Q�vi��0�ݝ�U7��z3�(!b��(%�<P)���Yj���+�ĳ���9�q�ō˦j
c��b�k�J�b�GR���	�P�^�����V����˳�	���}��b<�F��Bꐠ�z�@����rq�7��
���l�e�{lY<6E^z�Q��|�~��@+���A��9����&7r%���s�?P[�0������#r���>_̞(��,s�ʷ:?6��~	�\kt?���hkՖ#3�V^���)������	��Oϵ��5x�[#(�}ч���d˽\y4������&	S��Qr\t��]S�e��j������/Qf�H۷����e�ݑ�a���ܖ�"ӥ�9���(���X�Ol�c:����d[n�Vo�ǭ)�����YW���m^Ǣ�:�i$�O(�U,�G�'��Ȉyhs� "�>0r�l�z�e�:����9�m�^�<
��볦�ƺ#SdP�2|�&w`� 33ZI`}[K���W ��7~P�I�XT��L�F��J�f�"5��R0¾pnݏ>�/K�u�rO:�C*�`�%�0cr�=u
���L=�`�2�0��|�uqL2�$��-�Uߓ�f���n��v;�O�)A���#��T{�)�˅svO>Y��J���_��6�(��ǉ�J�^^K>�<Jqʄj�}_.-_:x`(�d�q�|���y��h��Nl���4��π��QH��c�A%�+�K�wn�ρ�fk0>F�T_N(�A޵��nK+)��z&��]�3�O��cV�� A�`a���;��.�N�aV�V���.�J� �~d ��zɆ1���R� ����V�,=�@-OzCn�	R�$���eٿy��D=�gX���6c̔�%2�K[X�
��-��2��M��cC�������xZz��0u��̗L�%��=���)&\(�"oI�[�p�`7���r��V��%�gՐ#�NȊT�3Q|��C��T�(�}5p�f�Y��sD����6YiQ�L4n��	<��Y�pc��A+Zg'�e"�����M�7�2+:h}Q>\C������쮁ui'_|�b�*Κ�v0v��7"���9��i�����F��óv8ۈ|+i��~�v�1�������y��/���\���p R5@o�L%H��%�'���o�5�8�OV�鞱K��Pk��fM.=��3��C)���c��z����'?@��J�t�t�qȬ2Fl=GkW�/��}�@q��B�~?dQr�O@���1�P�:��?���	_Y�$.��0W��a
(��<�]E�zz�3�3{��\�sƋ�&�Q�!W�}7H��z�쳉Y.�~WP�|��s ��U�Ш�Mis�
�aV���y����8�!��.Nv���&|p^�d&7jRb4ӳ[�����!Da�M��2�i��i�vFu=
�YL)�0K�~��;V�5�_M� �N}ӂ1�o8:o��T���$������jx����;�1�:��A|��Ϻ��Oy�N�(��v6d�L����������s���;l������t�w����r�v���ܛ�����鵈��0��hct��t���;���건Oי��O �Ir/�L��>;>&�j~pJ,����|��~���W0³�O��/N�9 �����Оq��oC�k���c���8r�h��5V�	��Z�m��:7��ѽ�P���B�ǉ�l�e��x�y�b2��P��2l����gYcI��5��p��}wBق�4�#oҕQ.\3\������<���I�J��"������+Y�ǉ�t��ȋ�� �~<���g����|֨�<�ͷ����W`���.HZ�{{FA�{��g���DE�~��i���>�sw�����9�!*�7U������)H^��޶�G*q!��n ��ҹ���Z�ҫ���HŐr,��1�����g� ���<\n�r�� �Q�$[k���	�a�����C,�9�&�F#j�ç.��S`8b���T�7`6߽��9.�Ec�$:�4#��eC�.cF�����b2�
��#�ܴ���P�ᎋ o���;���F�व���qsE��r�SY��x�8�x���N��C�Yܣ�Q��%E&9w�� گY�r��}c5��F]�K��|kj=��#r����jسq-��������C�������2Ar�tz۵�&'��50���6ڽ66��xĢ�����.ݖ�疭26����f��U��½��};{�M2$��5���>j��J��BNS��ڲ�
�����k&�x +$����
B��,�_<{e{M�E1�B�a� �^|�݀���&�>��o��&<�E���{B�G�z\�\�jҾ�x�"8ۅk�9��>��H���p6�p��9b7I����#�V`�:�9�4J�=eEt��u�9Pe�!���`=���L���L��ڬ�4�*OpY�-Hsi���^�M��x�\���uK!Z�4��ǩ���9zR��(#���1w-���¢�G�Pfvm�q��̉g�W���/��� N��;�k\�TM�:wd�5j�:�il�Z^&<���D�mə�Ѭ�����%vD�׋�GǷB䕬`dlb�ݙG^,����>7����^M�型��⇀�q}@c_>D��7�z�Wt=�bm$�|+<)e�����5�N�sud��[^P�$r��XR ��VG��t�ϖ?QIR���Ӊ2Z�ғHѥw��~��a�+�2l�ş紼@礭��3|�x`d��ж�X�]�9�����dRY�g1n����%@���.���5`���?���	��?:(G�nb���x<�?��ո��2��#���5���l���H$*�p��I_/sQ���W�2�y�&W�bs�ꂇ�w(��;�s��n����A/T�x�J=OHGq���ޕ-��u!���dG���@՜a�[^�H��B������"Ѳ����$J��p0��	0���9B�X�v��ߏ�:�[V�q���9%�M�H�cҟC5hI;��-_��/-��m��!j]��D<�Iz^����9A��+�fe��#!�__�l�|���qƟ2s���s��ϩ�[���'��R�T���Ne�W2�Azlo�V��_1�tGȨ�{�Y@�Y��\��J��%��{R\4*�Q㾋��t�^墷�C;���b(?���!o����W�&<(j� q�e�?]�,i/t���jb�]BJ�gL�U��D��"�ns��.v��/�'y����[�ο��S9U��ؾk/�C2���(�zjZZË8��/B�������K�H�� �1ms�NQd� ���rܻ|�rV�F�#8;u�an�8�<�9]U�罋�5��y��vx�/ʽ�C5Y<^����l��H?�^4MYSi���o�e6�S��d����� @��4��w�]ʨ��_f�P �& �^����Cڼ/p�5�����\���=�v�#�K�0����*���>���%vd����t��.�F2��Dd� 
qp���z�cYd-�R9��8��6�H=އ��v��qdG'm�Dt�{�4���V��|�?�)��S��#���?�;L� �H�����3�9	h�pQ/-������9��l�S	�>T�2�n�j=Q�=OB�T�����>�2�I���y��ãaw�7��-�0t��J�e�'t#�tJ~�˙ȗ�{�hfOW�t�_�O�~6軣�Yx����O�ߐӟ�|L��Ș�=0Q���-�Ȕ�)��T����W���-'٧�~��*�A�"y��
ᢊ�^�z������sL�W�F$�0{�S�d&�Y�U��U��#��u�	:(j��A-Е�$��R���H�l[Z�/׾s��ڎ���կ9l��az��FxV�o�N]��^�j�.�g��gyM���Wyԑ�P	���x`�a�>�s�	�S�
��fs5�"``�i`�6L9G�XZJť�K��q� ��
��9Ϡ�>�6�G��{�I: QqWN$����#:�L��IN��2�6��4x�5�[;b���7�^/�3`�.V`�Y���^�(���>�S R�D�gKKj�&d��#���D�y���S���� �?DW8������E(��&�������.�(�j�qV�b8LnI���M�0��&�m�Q��Q�F��78���B��L���"-�h�,�d�Jd��c�\[��\+F��k�f���>F�L��ZC=���ﮰj��z���kNIr�R&�����;�5�P��hy��٩Ik���Ͼ�h�b3���>��(��`
as�������\�n�=��s�:3ǚ�Z�D����<!0p�2?��d
jXi�V��1��l[I��6bo-:�]�Ѭ�Q���z*��;Μ���
�H���H�:�ΣU�*,��۟)���wr� !�<��N�4pB���ȒJ��*��Agক���5�E�0v�zw�L�'��Jj���Y$�8��4
�e'��[���O�_w���g�:�@�1
�� ��)]���`���qEFy�}0��ɨ�"�{f�xZ	�|JU�����2�j
�s��<�z\lr��Q���^6�ܒ��QE��A�BF���Q�����,��I�7���\gb��a�,��&����Y�vp����H�a�I�f�C9_b�۪`}T�6�P>%V}�,X*�P���R���5xTܕ�L���#�/]�m\b)���Xi�nz`T%�m�`�Qf���~���
L_$�nO��]��nZ��ɧ�փֵ���#k�C<[�#X���1k��y~,�-�^�7yP��`�'�b��Z���/jn������HU
o
HDI|N�C}��L���ē�z�� {_��l����pgܐ�[n��I���V4@}#r�Aqt�h�;j�\����O��Ʀ�p�]o�_���nGAj�#�Yk��S�њe+��bE�9�w�r����D�)�I>�9��?�G���N4�v�F2��R���%���"�%|�ʢ��؆�X�j�-�eqƋ"�C�!�r.1�)���m�?oON��DEB�z=m�;�>_2�ߡ`�Ze��e�h;g>%�G��O�?�IT�ʜ����p!��l7��Z~��+!@~\�;`��v2��oxL�hé�R��7���u>��8^j���2>ӇD�lٮ��ӎz2������8*�c�E�C�D�YF��{{� o�n�ii\�������X-�r�o�Igӥ�&�*��t�e
�{�ޗ�W3�̹jk1�]Q~JfÝj�a��sZ2i?��쎴]l/B�
�9�;��p�k�(*�[��=i6�9.͉-0����X��[g���f�������ZF6��ĸ@lW!30h;�܎N�yC���MNuߣpV�"㍾k�mI�2�?����?��0c㏰��da�"�D�
e���3��@�8G�*A�=ӂ�*	�b� ,���ܜ)�=Z��R`D��C�ｗm*Fȝ�yp��w�cޭ�!RC�D6�f���.�+�]�	#�#�<	R�0�gu�ҳ����̺�x����-3}YF/��ޢǐ<��C�ȸ��`{ �7&9�[8j�V��Rܠ��%,�j
n��iܻs��J��=b+�g,*���ĨPfD��c��bv!��ݥatSbL7pVO}op�弱��dωlb��=�q��p!af��L�ώ�~�D߹��9�g'�J��������$@f�+'�A�G!�!<tHx*��缈}�w�!������� j��_����__��Y���~z����|ң�ܼg
#�j�2o��E*�n%/�IɕY�es��n,���_ꖄ�_� F~�hH�ռg�Ѽ��b�4���!�� h
�W�&�aA�e�b+YD�$��쩨�p�_��H�E�!�"n<���ܯ1��:��ٓ��8��
���I����+Q�K��1k��4Oc:�6]����I �c�$o��A�d���XˏRZY]����N�ŕW������d�MJ�Y�(�?�O@�N���N<k�iB\tH?<����S�cLjs�N�L�C~�2u3Z� �1J�KM�9��Y<����
G��Z���rkҩj��gE]����)5��"m���^[|�hȘ�;��d0��O��H72�S��#|H���h>�%W��	>�Mlr���P��'	�M���jb�g�6�F�)�3��o�z�~M�`���Z��z#3ȫf�s~��o��JmfVGO��Kj��p`s�.���"ߖ�O[dh~%�mi�ԡZ�X!��	�N��q �x=�UCL-$� ?�D�jb��D?V��=P�r����k!-j��A�ƥ�7�,)�V:+����X6��J�ְ.�a��]&趍p���u��Q�20w2��*W-C[�=Y���t"Cq�u��ԇ�Gt��%�����i�;���J������Q�ph�E��I[��S!�؏�$yd���-Y�:<�6�Ր�x0,������7е��`�c�oGG��[k��!�=FW����$���n ��y� ~,gV��n�a>ӵ��`��s�*�4zn5�b�}>�� ӌ��n�j�UE�Â2�N]�	\3����jT,�E�.t>PEl( ]꺱�Lcە�┣�tA�5k9$���\^�G����da���dU�dcW��[�e��&�Wd*k��^���X���[:�l�{05ڜd#���@��f���� �Ѡ|�2��6�\���R����ٮK����9Q�,^ �wI]# ���nB���'����:"&:����y��l��pHu����Y.�q"��_G��D�S�&O�s��,�'.�0�զ変��-s��i�:�)f�t����2�^�PZVWX�z�'(�nC�G��F|�`8eKP�f�-�Ga��$//Q�ҍ��� !V7�*�8���2:L�.� hg�zf"{���L�bA����^�t��g�z�1t��I�uf�BN�����%-<�z�34������r��U|c�Ӟ�sX�20J�w�ۍrn]�@�"�+W��#��!Ca�v����ZMi��F�����ƻ�jz���з���*<$q�CXV��Sз��6�:�ߨ7'�����n��T=�
U���a���6�l�8�j7�
��G]|?ԣ��2A���)�0��[����	2��wj�{ŉ�"�ji�cl�˝;�ig]���_`�] ��7�[%����\4H�$J�@�^����ur�A�Gi�������&z�"y���"����X���9���I[}����/����Z�鞐/�Y"�Y�u�K� �E[#�k(����H��'k�����s���{�n�d}@KgΎ���ʧ��������ȃ�9/r�d���{[T�5l?'J�{_�=�VV�:(0C؝B����w�^W�~�m��;}%Qv%�qU�g��(��iμl
�4G�)P'K��Fj��W�9�~ƀ��U��� ����*g�%q�����������v�t1���5�#��_��=U�}��l�`Ƹ�y��b}3��ܠ�E:y��H�+Z��؝
	�����J�0xOO>��9�����zY���#�&O��� ��I����4��S���9�׭�߷�O��A��< '��@*�Ѣ:!VW��BF��[��Y�l���2�7py��_�$hVoR�g�<W0*x�Ʒ���}�eq�$|q��Y��+�d#�˙ȷAx�q%����P�+̢d$Y�xo^A,qTQe�nJp$w�����#
c��e��"wM}�ѩ5DN�q����7Ӡ�<�_(e@)� �Z�fk�(��b�qz(d�PL�ћg�(�z,�9݂�7H6y~���G�[�H%�C�E��f�ʷc��-��
y�f��6��[:��'��X�+y����U��h;/�m��ɭ[-^��rTHX�P��l+�T'�=��z-�F�yZ�Clǅ�<	w������6�!|�Pܠ�AJb�/['r|zR�  ;v���r� ��}�4��k2	t�2��yL�`�M!�V]w�.10���AX� ��쬳���P��qet}E��y3~����Z����%����{	N��o;�8J�#����O,�ݞ[f�^mѷ�q��Q�oP���G�9��p�1$�$Y����&�E�d\�#(gp~9�V��Cݮ�Ys~�oG���Ɏ�ƿ��~r]���8�m7���6�ުʭۧ�z=~Bmm��7����[]ޛ�J`��dۋ�qX�.���"��Rg)8گG.�]M��Z	/sA��5��+�)�H㘹��(��!�M2vGд���58���,�_ �����2l��%�P��%�297��*1P
�24{�sإ�,C�4�&A1r�eW�������3�~��^v:�"׏^����X<re�g�~v�}��DS�-gWe�4�g�[z`B��E�e�E!wޓ`^�ӆ6���I���M����O�|����1}����.P�mDB�d�k�LY��Q̗�Q��A���J�|�5���?��!����Ə���A�I_�3!�s���,�h��
x=�P�����g��l2C�G&h_g����#�*����'��� ��٫71��� ���M��Pv߾��[~'ى�M�v��fzr�o8H��R5 ��^��?���(~���/�S�͎�H�YlN��pS�:��u�t��A	H<kS�K���n�t9�t^��ć�������<љ�/US8y$���]T���I��9�U��@��WP����d���*�+2C��ppwVIbV��� �8�3�
�G��X�2�| ���Xǻ��Lj�cq�ܜ�t�=S��i���|�fR����X��T�1KB��,E�0��ákU�����Ev�l�w	�g-x�
DU������&�B_������®�z	�p���S-����c�0�%�m��Ē���
ti��/�
�t7w�`D>�Uә��t��:��}���sqk����꼇�7�T^]=x��1�f;$����c�_�[S�Ƙ���FG��L2� 8�#�Uy]S����Ci�ES>O�4?�sU�i�&�Њ�?��"�R	�6�m�>�)�|4�./W���M\�q(�5����=P�§3�|q�X��#:�B�EA�<̒x,e��x�k�e��]�}�I���'_y,�5��W��wzx�Q�u�����`X��C�e�{9ih���U9��U��w��1�������E�0ba:��_�0�*�lf ߙ�S�y���Ð ��I?�˝3���Z�ԱG?�-����fO�WA�8Y�L��S,^F����j� ���<K��t�� �I=K;��t��<:D�.ϋj��C�V�p-���X[���@�C�a���O�����2��亂e���[7r��ҽ�r`@�Z�FX`�m�m���~��9�6�6,�U���Ky_�!�k<[F�kkl���i�#j�m��Rbs:G����R��]�!40˚�f�(lZ�q8T�휈*��v�b{��J���>��^�3�+B�/�Y�e��l��
�0I �r�T�����RQcWZ��/�""݄Vi�B��8��k�����RkѶV�eV0�� *g�3��̚�/��&��W'y@�'r$N���i��X���To\��(bR9�U>۠�&wt׭GB:V��nU��O��㗤 ��]jk݂z�0k��_U?�G'��g&�^\LT(X��_}��~lpV��ܧm��m	�%���%#^��iw-��5䣑+_��������j���ݢ�H�XjM�<x�GE鎅���I)��cʸ���o�i������]F���������&K�P�Њ'��ݞ�u�D�9t�Q�J�tS �i�(��0@�s*������\}�������x�fA��H��E0jWtk��
�r���b@#�Y��L4m7 �7����`�*�ؒ�J��_��+ ���O��P�%Ƀ�b�pw����7�9�=���M�j$2�/��fma��S��	�����F��-:3�s�ŐZE�?ب0���zH�"9��*��%�2U6DP�^���G2%�vgPȏ�ׅ\�B(GP�-���/���,��"ǻ?��*���2�����h�S��Bt�)I�P�b�TE��	\zQ�aF��ھ�EGp�mE<�,KN�Ж��(�,N�zs�Q̆�XH�,Z�gWꋶGm�r������J��F��y�/��\X�d\�����$u*4Ik]Vմ��)�۰gE�Qzgqu�Wh��a��8	N7�N{2B�G%2w�p�_MJ-nO�GW�������f@����ʅ���_Lj�$I���R)p��.��EiBM=B����]u-n�R�p���"��[���E��Y���(em� ��K��mx6zb�& �o�I5_�SN��u��?�
��1>�AC�|�B��Q� �j P���2���\�4�p又{�l2%�L���d�d��C��_G�D.	�ړd�0.k\�'q�E�*�G���Ƿ?���v{qP}�Y�pL��¦���|f��
��N�@�u�i��w,P�☘�{��!
��X`'�>�K�ݔ�|�U��d�?�je�J�f"�"��j�e����̎�������=%r��q��0���\=;(H��-��<	�'�����n,Ž	���Un4�E����6�Λ�����3CzN�4�6�����F�`D_����=��z)e��$�4���3�pε�]:�b˘K�$�}5���7��YE�z<�[ ��b�,��s��Ჾ�-���u\ԁ�OFh�s|(� �186�q'�;_���{��5�LYG�6���n'N�DA��̩��e	�W��e�Fqw	�TkL�$�����e������[�����#�5�]��K<�b�y(:q���䡏�E�SVU���S%��_�E��Յ�:4��m�"�P@�٢̓\�J�ȲV��t�ed�'d����>Z�O�6R�E�B�6e����4��٦�Y�M�dv��,茅z���o�::�d��p�<`�a���b�-Q̼2�5�����^0�~4.��3� 63yqJ�i�k� wpLo�"|;&a�������I����o���F��JT�Ӥ([T+?Mo���=�~P�#`���uF�A��|�Ք�d�-��(-:|kwF6l�vo=�;�x�Dw�����>���X�?F�����W/ ��y�q�׸��߰�1��l<�� c�@u �����S�4��Ml.�^�5��CJ�>��HLޤl��q��3C]��˷���ڡ�e���F��it����������f9�ڡ{mw�aXL�Om�k�& q0��9[�Zo��\�=�3�vDN���MEUZ�d*���g\���O�=Fw%!`�R�sOĜ����%H,��	���q�������Q9T�Q�-��ߣ �A��F��l=��ׁk�?wӳ�@��pQ�3�o�B��p�S ��/`����eK��5�t4\൴�ā �����l���ߙ�����7=&1�¬D{&�9�x����A�)�[Qx
�*�7X{������r7���J"?��a�~oMu�K�mA��3q�!�E�o�	p� ��pr���ws]�z������L�u�|��x'*��4K�`K;�7�4?c�s�5v��1.F��T�/Q|˗3 �X�;�Oc��	������@�9�L�k�G�����IW3��
�����7���05��loh��"�_Tb��.';J-�P靾�!��}���O�G'f}�h�!�Ze;w�����Gp��Ы��s�`�����>����������c�(�*��O6o�S�I֡�^����a�\�+!�Rz\����2N�bk![S�(6�eZ�����Z�un6�G>m$r����]ј����K�^||��q��p��!�>�*�ط��}i���G��'�CF���4Z����1zC J�6|7�g�I�t��M$��⸠_� V�ϊr!�l������l����X���Aj�Ij���O�#�ܦ����lFD��!<�)���1�83�f�!״��L��)����N�
�3�A&���h�md-���^r�h����`Ι]�cn[A�Դ�0�V���(�F
��X�S[�ܠ�!m���@���+�
DTw�6�,!n�.���P	t h ���U�:%�n��6����63��i�x)�	���&j%�x���F�t/J�� F�Eq��}��&��ɪ���|��({4��4&K�<���v�RTݔ��}W9��°ۙ��1�j��˽���~&��`i*��M�4W�������T�,���r��bT5'���[���!0H�������y��ӻ;IiP��ɷ�W�7,Fk*�x���A�~���0�9�6����P��<���f��,�b��񵘝ġo��E��Lܤ���V���Hj�oEPX--�7�\r�? :)�e)�qg�&��m�z�d�� � �z����\�~������^i%��]�"�)�xPI�Km�������s�t����l�/?�Do�l§j借�����0����,�d+>���`Q�#k��օ�?��>���N$�<eCҝ�nq�H=`l0���|������k��Yp;�$�|F&�sK,B3����P��zewy|�^i����g�NKb��.W�.Ć���.� x'��I���0[�"I�w�Rf@̆�J^���42=��	
���w�<��=d?ժ�3����#��]d[E�L���X,\�����>t�Ƹ*�	�zݺ�@����	G���s�^v�J�PV�����p8#�8FM�]����N;JM��%��Gs{%�8�W��ǚݨ`�9;��� �f�(��"k���2� ���2K����03!�^{N���k�5|���+���p��,�7&����t�u�8���8!`p�B˙'� �4Y;0̼4�'`�����~ B	Enp�dqt�q
}�K��Ő���T+T	u��  I��������37z�x��i�e�m��ញ:j1�p�5��Ie�m�<�˅��\�9H�����{���/	��%�$��))+��9.�ۯ �**N�
�xu4���:��߮MfP澖�sv��SL��'���[}vE�+�n���uβ�+�TF0�����2Y�m9�F�N:�(a�t3��|����P7U�7Na7��S��rr5ֹ4/).X�lK3��r{>��3m6*}Tڲ���,{���%��:�)��"���{�"a<UL=����rܙ���k��м��?a���\�Ͽ`Y �e����|&�j4o�P����#(���:0���+.��e�P��hީtX��.��̗�c��_5�*^.}���f���O�?�e�?Rx ��sw�s��S�Z']�%�9�RV�n�̀��I����9�zŜ:�8_.\�П���ky|����+��<��y��~x���6#�X"���[���*������py3e@�8��Q�R���KHd��IM͇�)�+�!!�$�on�i"Ý�I8#�xxƟ��Ľ�������x��lo�\|�u���|�AS�=�wIŊ�3�z�w��^���όw�({�.3=HC��7��Q/�!x��U�*�,�穰���t�1�FY�,p$P�%���0�)��Ӿ�.y?�[���Ǒ�8v���3�W�a��s���1)�*����D�avY3gza�O����B}�q֒�*���'<$wM�n&@e
~�i �@���?�䣿~�N�@��!]�>A��~.�Y�Cn���てr�4���;q�TW���8oX��yL���7��'\Woj�����M�����C0Om��4aZ�y��g��j�)�Q�&�1��!c�K�{P�AWy����n��̡'�{8��l��ܻ����˓�� �#VaQμjNFpj�+��~��ak�?x��=�����-Fx:���3�$�6��l��U�����@�8-���Ű���2�����/���j�z�p˥Z��J��B��5���v�^Kr�W� �=��U�������DT,�'U��[s���뮰�-W��C�"����\��U�n,�ߩ糧�
�)W��HŋYÎ9f��3��ڧw�K6O�igF���m~�r���/�E���_ɵ��� ��ۅ���L�%�w�T/?��u:�h�ueQ��aA��Ru(���!�dj�`�Ī���㿾�=��,�E����^�l&w��� ص9M�=���"�N�_Wp�g�s���L��$8S�z�HI�iʓ�AT�X^R��9�~%�P$pHf����1bg��]7�(�wZ�q�,2PԪ��o��1���x���������/$!&u+ky�������<�Q�u��8D9���2m�����قn#F��#�[	z�|���������\�I�m�� �qmOT�uy��y
#�n<��~a{̰y*+�t�
{�/��Q	�ui0g������Q�D1]���@M�A5��������3C���!k*�C��&���OjD��Ku�y�J�S�]o�/ZԦ�aϿ,����X��O���,`�L�E�)w�I�s�;�=7����ۍH�-R�Q��E)�s�I�H|!��(�"��MSW8�,����(���u�x�����B*��Z�ӥ]��>���S�go�8#��dՏ�Fp�G��~Ѯ�v�2O/�|��4�dՒo	��P w]_NW#��Ψ�-�q�i����Q����gn����m���XsN�G���n���˩j�:����ij�0U�d�JV�R�@�"��A��*�J�&�Nno�=N�KA���iI� ��@O��'�qn�_-s?�;�C��!ө���]I��&�cF����11�2���y]8�K�:`H��m8���Α}�ȅK�~˪��w���8)���<���y�)#��r���;��L���H��i�˃�F3q�P��l��"�Hߚ�/	�w˂0���`�S.�8)�J�{�W���C�a,rp�ɵAF�X9������n��|�W2tJ)��|��R݃)���x@���5�[Q���
�4"hE�:T_:x�ry�D�CT�B�I���u(�(����ｼI�~�,L�io� ;A�X�U&���Ϲ�ę�|���YKw��~C���e	-B�QGk{�	Ci��s�{c�mk�}��T
�[��v�ar>0��?{R���P�4�R��x酓���G� �Y���_�u3�8���W�6E��bU�7���=�R��p��F�/��9��&O��35���5TH�^�z4�������|�Y_��&M�~#�������V7OK�a)���h�=%���g٢փh(v72]�w�	�=x�y��%,��@Yj�!�*h|��,��.z��~m���2�
)�E�ђ򠓰�K���V��`�O���F�!�b�y��9(�!7c�r�b�YrnGǩt��8�cd1���i��<G����-_��`�aW�FY��V�M�w�5��P>���A�T#`���N������sK��Cl�ڝT��C�F���!�SF������,� !΍i������ܘv�`�\1�������$6!���N�m�Ϛ�j�X�ZVl`�1݅�B��U��/��e=R��Q?�_YR?w">f	̮,��,+���}X1���55���ݾ��tH$o�8�3�[��K����^o�~
�r[S���by�#mi�-�.�N|:�2��xe;;�W���:�S��qw�rY���Y��YHL����MB��-%O�xWڰ�_h��K�<���v����i>��a��]h�j���#����D�X��`ƒ�g�����&�q���Ю�,�Qb��y��Z7ṗ<Nn���$.��M,dt�Uux��Ն�}IRqQuu�m�C�� �����^�YJpVڟ߁�1>��p䩐�~�/*���d�O�=���r�l2�I�!�ކ�=!���W��4R�ߗ��6�Jy@榶�.9a�L Qy�)���s|r�Z�G�o�FlNZ�;��<_��`��~V���92��s�l�}���p�������Q�pw�u��'P�~
��~��}4́F�G�~b��_6M���߆��.����h�[�C�*���/��4�j�5� HT���}i��weX�D�J:)�gpZwR�c�r�Ԝ��r� M��H�5��3NJ^�����7?n�����-,��1D�X����-r�ϐA� �*�ťyCV���`=^Ţ�yߟ{޷v#3�+��&DK'Q��w�C�c^��%��Ԡ}F�U�_��mr�-��_�}H�S�|�fOeV��	*�
�`U8���k�d��)�7%�88���Y` ��D��U.S� G�O) �`(Z�5-F���Er�Ĺ��K"�f�u}���xFsk�Tk�`AT�w�<���Ej��ø_��B�6���m_�Q����<d��e��i�d`�g+�
�H@K��0�q����=��Z�3A-����$KX H*����66]3;�|40�����x�\�Xd93����k<>̣�����30��h���K&ˎ��w��w���(��ґ����{�d[@��)O��ƍu^yXܛ����H�=`*� J�L�@���:�K֥�g	��7@�Pb��bVb�(
]�z�31��f<�2!h�u�tTy�=MS�����^��������x.ؤv<�M���l��B�6;ۨz�2��2����5H�������UZH�'���U�T��ʠ�䂤2Oِ�c���L�ƚ�~U���\�5����o��K�~�9��� `K
3�k);8tV{y�ht�I6uj���UBj��0����M�[q]sS�^���'���-�!"nwt��n|N~�B��c>M{��-
'c铽iK��噚�TD~qn�rŻ�	!~���N�	�O�y
����˙���J�y��K�f�dJw��x.�^x�2���bn�:�v�~E,�L���ԟ�>��G�^�,�j�I�C�1�,�h
Ǚړ`�̀��n�!����}�<��&3�F���=�(oA�ۋ�Y1f�;����jj�����Ƿ+��-�ݞ�<
�on�1�P]���޻6o�����}K���"�	5f�1�±����&|l��J�3]��Mݮu���8��}9�M���#���#b���7�	 !|�9�>�n�ȫyM��j�*黲41�ةf��(��k8�����] ����Zu�m��rh#kd�^�(7lp�v���o8��\Ӹc�:�)rNG��b�ij!�IH�
�"��
cu�X�W���[�s�jC�j��o��u�&/��j)"�Mr��0r���9��e��.7�����a"h@���4���v��(��I�����?#�Ң%!c�T�/����{��V~*Qe��� �>m;O5�k�;�����tVG�2�bJ� C���{�]����Ї���6��׻�;����!=�X�W"J���1������_�4�;�t'�bҞ���
B	�.�zr�?�	���wY��p���r�Z�K�_�xOAkG<��݉��|�P]����}Mq�,�<��t����aw.��d��{��9x��	B�@��K�J\���;un^{���_��i��*�8�����.�G5<,�����q�a*��Jo&-d��$���ʹ�"<!�'��Q-�Q0+D�������A��o��`��G�C�,�Y� ���>;�4�����dG<�0��Up.���epM��?�x�S�8�HQ�D[�<��K�zj�wu�yg{��o����}�Y�@��;[���%$մ��U$�\�Vc�t\�]�vUX�2B�~�K��(�T�$>��]k�C��)�v�~o�~�Z	R�����Ѽ���J:��6��������es3j����x��c]����y������0��*u�7�"���`����]��D ��ل�QXi-�^��U�A<
��(=I��n�$��e;4'�е9���9lG�a�ѢҰ�j��Έw����z�^kqȝ��`1;�^>ǀ8�������ɳ��
\Z1Q@�n~mi^! 7� ��F�������U���3���Wj���l��'��{t�9�C�p,\���M����-����H�ڨ5F�\�4=�V���H�����|�un1):l���yڔǓA����0f��j8����r�Q���-�ћ�؝P�g` xAXx
`|L�q2W����R�@�m���!!������Wf�aFN����eIΊҮ�1�4􁳟�S:��C�գ�?X�Cy�����]�%r�p x�7���^cxKL�d�z�B��% $IH:4%X|�����r�$~wz�5lb��P�N��������&2\,Y\�/�"�w������E,��ZJ�(���ГO��mA��6@���$�6%A��6+9:��S�r��pxTѺ�iΉ�JD.�G��F�e��f�����X��أ�����G%�A���]G��-�}>����m��ϛ���[ƛe{xa��=��_�=Z��4�?��T|}dl�)o�u����u\Jg]L]X��g��{��y�ѕ����n��Ad��.)P9h}s".�\I����4���f��=g)��ESZ �3r���:��"���������j^]��[Q��Ƣ�uV
�f��臭4�b?_'�B�����&�
J+���	@y�"�o�gSo� =<�8mѥ�4{7Pq+b�*��m�BM���W��P��]V(�Z�H��ޅUʑ��`��E��;P>�B�^Jȁ?x��6�©!31�zu���0�L�x��en������Ǎ�̶���.��£n�fB(�������!���vL#�sO�_�7�>(���$�N�ɸ�"��٬�eVN~i���B,0��iu:���U���9��HC�d #���`�z�NZ��]z���nc��Qi#k��*}���f[�Q~��i�&����e�a+;�+�1��B ��?
O"ߒcͤ�`��� ���XS�G�igy�\��=mr�6��G��:��K|�c���% �}w����E��oA�z����[Df�}�ߧ�Ǻ��,���ʭ[X����ë�c�����	=@&;#����E|���}�x4�c�(�-�	��~3�$�x�ho�h�F�e�
�����"1B����C�H�Y���  ɖge���L�cd*�]�����?�@+�d������a��D��3�2�2�[pR���IZY�7��/n6r�G]�"rF��:(�����\"�A�����|"ž/���Y������i��610��m��w��Ln�:B���.�bf��y�C�w��T?�|��H�I��K�4����`C*J�rc��LRfW����2��!�f{B'�
��R�n)(��q�HSg�T;�T6m�¼x���ͳ�k��拉��}���W�0R-�&p6O$oG@�'�4�����@.v�1+�}4I5$�������]Z�. �*Ne%Ԧ��_��:��؂ǝ�ej��-{Gl����/N�q�l��=>)#j��l�:u+���Oބ��1�WF^j(�3��Oj�!!p���'���Т��%m��N�`-T�u���j��Ĝ ����X�}�ʽ��@�r��B>�q���6�c��2�K:%�BO�-X�FI�:����}ſ��
�4̼]t�v
*T��)�m��m&X+I ~��)���	2��8!�w���9�e�!\�u���7YR$��W���i���P_��������g�`ͰX�U��l�z	�ڟ�/���1��r�:v�|��)�%ģ4����٪o��FAO�Qd���F^i���v^�aO���]K����,�ƞ�L�������V�0�0�d �V}�J�.����=�Y͎[���X��9!�M�4��w��
vO�M��(<�U\�����e$��oX
�}wO�%��\J8w@�p�ɒ�����k�.X����d�Uf�b��x���*wD��d�keޑ���~g=�	�<�:�/
1��p�7T~�0��H�W�/Wy=�$����'<��qݿfd$(#�Զ�v�b{#A����� ���?d�����*(�\�-�+�1�݈�E�3v-�{OO�8�����6��%�	4�:-F����3#w��\�%G�-?F g��_���%Q�݉f T��?]�>��W��Yy�zRC>��]o������4g�JB����	� _g $��A[8��j0՞2�hU|��s3���)�#�I�
����u.�{e�+�W�jʲ�E�T=+]<3j��?�U��R�����<V�o9���!�`����ӄ4d�7����7"m>$��L��q� �W��e��	O�q-ل�#O��.�ō���*�.��E�D|M�z9�HRfH�C7�5�v%l�f+"o)s9�f��+�>�CD�{��AHXG��c��mf�J�� �$~$�Ÿ౦�B�du����\���*0�����⥁�_ylg�x�ϫ�*_,=5�T�96\6ɞ���Ɋ�^�-�����F����O�݊K0�����a��Uh��Լk<�ݨUu:�k��_(��%�����>d%��B�hs��2u6fڗ4�-;�J�%"�|��bK���!ݹj��� О��"M�+�z�Z��fdC9�T(=64���0��E,��o9��eܟǭ���}J�y5�����۷B���M��$x2��JFh���ڹ�dV���Pr6�~��𘅙nr���'=���1���}���2�����(;3%�v[)��j���
���" �����"#p�]ŗ��R�u��S��q�>+�b*w8�y����{��P$p���j�cu����K�X�I���.)��9,Hi)5kP$dOՎ�2�ܟk�!E�۽�p�F��swd2cj��#ajQ5f��V�@A��ɩ�)y��Bw� ����ZF¦r�X���B�#lǃ�8���hEV�g>m3���6ї���&<�4�ΖHے���iYb�`�M(���5�2M�1Α��guӗbF��l�Ҷ`c���1�PMuuғ�}d��}cHP�%��cD���"��`�#m�
~4m���$QӇ�eL_e�ب=��<�
kS�m��Ɔ�hʋ��ϪN!�ɒ��π������C+�
���.��[[�GF��7����=�������0-�x�PKΞm#��qb�>�� Ig���%��*�M֮"�Ub����E�[FO������3	مE?_]v�ɾ�O筴8�s�<������49E�EN荁��x]�����f�,X���eF������d�m�$WZ��8���B�!Vp�G�"�S�:�b��M���� .�w��bع(K�k��g�	FV8�-ro.�Тa�����$����4�-�{VO�`\Ԫy������&Hd倷	�g �{l�*:�D�����K��8��J<�)��+~�{0�f[���᭸��}�����4A�}'�q�����K5u�&�+5K����JO')��H���r_y��T��cHel	Ý�y�Nʧ��c��I{�ﾕ�E�A)�ӈ
��f�#�l��X����6f�`��1�g�%��>�g^�|��e�O_x-2 ص����S4GBVI�Bh���u����t��a��j��:�����!9#7fN��|�.*,�&�j���"�0F�/��D:a�uQ�uf1�4�3L � ׭s���oM�8e^�Sp�������C`&W7�e���Nn
& �!;�E�����c������<_�YC*/���,ξ���t ��U��^OBS����/��f>))G�%z�G�6/��+L�UN�&^���o_��X��HEv�Pۯ9��hb����Y��)Q�Ah��Pv�xQ(Fۺ���Cg%��9������������,
�@ݿ�a�$�խ\&�����!2J��V�╍�lY�� �ב^y���:��+���D?sTS���3z��Ϸ��IE_j�OӤBb��`!&)�����T=D��Sބw�7@ ��ߝ���0� .ݝ�̻s^�V��YJV�jGs�IuC'�ɷq��ȵ$��d��]˥�I#X��>�ʛ�.�[���dp��K��k<8=*r�S�E&kq�0��^��SCZ�;C�J�r�?]P� ]V�s��h�4��ͥ��u���9�n�s���&A�i�J�
�3�W �r��n/t��U"H/�ǘ2�1�q�	�F�<�E�����7��%4���{$G1�'��	�Me`�,�Bux�/�A䜻u��y�ZJZ�A[t�n/Y���=4\����.2b�0_c��g�P[�+aV�Me���!@y|fd�@w�e�  �hQ�^��[�W�q���.�#ގI��-�% �{��T�ŊQF���8��Z�oԬU���9�qd����#��r����=��)v0�K���%������;a�;y�Z���7u6qi�G2�mR�z"T'A8�)��,V����m�"{�nO l&��=��mb#X��8�8/0E�_lY�֣�`Ca�E��U�v��~��~]W�%����;�F�>H:�vyr���&�v�V{����/�i<��ȬAJlO�T��x���������7�����ɍ���"���������c�L��u$�-�aETLP�.�<��@��վ�#v~�@���=�c�)n�vE�>ySH��_����E�y����ht�>�ꠐ$}�����S�%B����_��x+���������g�\G��È�ϼNa�fe����7��r4���eԤ_ʵ��h��u�K����"��l����I��	���F�ͼ'���/�JE����~ՑZa�d`��b������Xbx ��{H̡Py,OC��|f�7W1����g!�at`�qȐ�>j���*��*W�BR����x�^@@*�Q��󏦆�b����.�=;��Pʫ���SIp����Ԡ�h��iAE]?M�\�)z�^ �>�*�
��L6F޲G�];��,��]��*�f{%|������}:�
W� |kdYT>Wce߅��!f �;������jT;��+Y�,$�U� �Q�Cv���:��V�#�K&^�&K�9�i���J�E�@�A��*늧��Fe�b"�xx����/ۏ�۸i���&�D2�m1��,�-+�v � ��:���}��J�E����=��.��H!wTz�OG��x�88�� �����'��+��+nO��ppȏ�z8���D�(�K��ڏf#W��+&,���7��`�cH�܋��S�<�E$$dr���q��\�?��v���T�U�K�ף p�IR˽��u��J�cSƀ/j����%d�N��4ksK�s��4~�4�ڀ��٘�B�"���˴� Xm���]an0�}b5���\F��n�v�?�x9!gM�����U��ˀZ=�p���H�]���GSkΩO�Fv2Jq	H6 �jqwP��� �G����:�t�E38w��Z<��ċ��,�q��h�v�� �3h��U��hM#��*@� �h����Doͬ������~�^�ꔳ������c9���v�Mf��_�ƴ�zl���ɷ
BG����:�ܺ���������$���$�!3���0̆�;�T�|����Ϋ�`l�5�2L��8Ej�b��6��+ӈz� ��8=^G�Z�eR�y�W�i��FH�V���(�Ǧ%�~�sS�'|T�$Fң�֒��YVE�!��ߑ%�A�oȵ���H�(��\x�\Bv�;M?�jm�Yⱷ���/�L#/��N����r�z��3Z���Pa�JQ�8BMp�"J�1
�3�]jj��r4/��[�m|Z�ЃD��o�P�U8=MD:�,������������"����Uv�Q�D��6�j8��@)�:��d��3p:5��-$�?-)�n=�ԛ�RnJ봐�B��[� �%���b�o=����;y<gX��a��"���o�������͛"�������K꼋�'���ԜDu�5�5ͪ5�p$d���7Ea�B�ߗB�9N����@�x��s�j�lUf/".CR�2���/��'@�(��j���
p��d�]����S�o}�������>��6G �3U�ױ(���_՚8���c�C�Ѿ`A�� *K�j����Я�L�\��L������2 Y������]��e���P-�=ɺ�]ޛYM�nI/JO���k���J��[@+���>�~ǳ���c�;�Or��gd����QJ-�/)e���<���P���m�u:<E�ġ��?~�ij����#o��7���gG��ء��M�' ��)����[Z��Q��Z,�/M_�d����j�C��tf)z��'m��9�S�jy���(b���uX �\�'�Qv�uBe}��&�H&ˆ{�n
���"�����VS;�[�׎Ҽ�u�<�z c�|��CGiU��Z)0bm�w����Eq�ua̛�2_�hAF���p^��s���{Φ�m�g]ɠ�����fC��JF3#��@���ό[��HR�h�j�-�����×	��D�JR\�B��i6rWo�(�Bc+�'�l�N&�iC7�!���%4d�͗��T�����,�(Ԋl������	3d���!�ĄӍZ�g�]���`|B�IAVʩ������s�/��:~���oYN�c�*����f�Ӫ�HYq�*�TXBU��7�yK��^�EqY�ƻ�h��J���O|p��B~v4�Nkrt-�e�kx����Wv���^\-����2�6p�fl"��}G\oh7߄�"?�q��R	h�A2���U�܎很������-e���ȐPyQG�(���:��#7�����8dtm���'m�� ��K(������M=j@�h$��w��Dl��(0���r�kv ��عb��X�Fѐ���GVj?H?�D�$IÓ�D�wmU����� q�"�_]�jc[3�[�����%,3�T�	�۶� Q����žkS �t�ݝ���$E3��KYSN�9M'�uʍ��Sk�5�Km}-���zTS��
��jK��6����˥�f�S��|�:Xl���3���{'�ja,˷v�0wRO!��v�
���cJ�~�!��?�ů�13�i#+�$��͘��5�oۤ8�]�^H����~���'Ez��rt[��m%o�8�0lj�������Щ����q�$����t?
1��эM��-%S�xC`��<2����j�IXZ����u@Z�Q���3�:F���P��];���.yK�3�<�t�-�[�!�p�z端��Yn�a���ꃝ9�h��S�w⯈����G��pǘ��0؊��:�z�R�D~%Gs�^�HAG�w(�������s�<؉ѺyD*�Xֵ�\��d�IE��.��1�=QɂH���2
}��ן6ӟ��^����A��*�v�����L��i�4�g�z�ڛ�g�ͣ�zD򂬐v�(M�Jc��4�a�ek��/�Ewv/�DN�.^�����nX��S�#� -F��<GC��:>f���h��$_qrD�5Kf[h��dq%��L�-�����6��_Y̤"�dj���"�C��q9rGgǞ1?������{5������xz��X^_�BZg���[��!���o-�x�N��p���9"n�@�lR���D�0N�#���ڏ�M�֤���� ��q��IC(�*��2	����[��$u���D���
bH���=3�L����|.�|�mK]1||x0!0�rއ0�M�B�''Ʉ{�>�����G��-(68�ò�$�M��� (@k�=+�3x�[,?��Q�c���z��$s�g�N��H�>�8���2F��ކ�z�i�ֿ�ӕ+��f�UU��+֡�=ٌ*&���l�/���l�W�[�6ԤN2���i�4,B+G�GP�Ē�ޫZ"U���W���^cK��%��r�=/J��Oǈ<�,���?Y)���	n����&"w�K<�1��&�P~���U]�ɉ�ៈ����'�&��o����2��+&� �a�sۦx�D�M��,5;�Jf]v��Do�_�O/�O�Z��Ȯ�{:�e��n�5�+�"�x�{'g�� �M�<�b�C�|�G�J��O��Mp@48�(��1~�t�;�/�g���t�Yo�r�'֯��.B�k�5=�k��G4P�޹O���%�3�P�i7��ETG��6�#uQ��<���/0u�tPL�ѦD�_@�[T���݊z3���F����q�=ɺ�{G�*[]�������Y��YrW�9?Ë�W��?��>P���F������[�=ak͜���#|�H��Q��<>��<c��}l_v�
��_d�E��M�p�@;,KǇ�]DIsZ�}r�d�N�A��9]���ԯA%TI$�?�N����A�' ο�o�q+�<������o�n�ص����M:�>�Lf�'L���0Z�Q��b��}�/�Rׇ[�YzTLD'��GuF(Pxd���kUə�x\/e�	� /ht�9�y���3@��5)��g�)�`�tDH�_�p��;�G��ȱ�7�GE�s~��
����7U�F8�]̬���HLg�-_�B�c@��wʂ%�Ĵ]�qg�B'v��鸓s���/�������.�쾐�W���>�90�P�(Q=�2���j{�|(rˆ�(;�-�v3��ͼ{*+�=/HI؜ �$���	>�+:<����/ j��UldiD�����i�:����O�0[T���h�W�'��`��I�l��Pp0����	h�<�o�Y�3����Rʴ��h�N�-+|��I2ZڔK�xY�.��L�&oW�>��䜬�
o9�7^��5�����P�w����*���L���yA5K~�5m\ǩ8�q�0�=O1��TN2%#h��«�{"[���^���f�1�G�����x����<�<l���ؐ�:u����~Z �G�6��z�,啹:0�z����2.r�0ꋯ{S�X	P���@�KS%2�5𙋝	���[�O�α��3{�iJ�?9k�ʳt8�ؗDk}����I,
8�(��嫲�q�&�i����5`��֬	V	5��+HO(�r̡0���Okbó�&������YzϾ��9Ǩ^�W�0�Q�<�vO�ת0e�vPQ^yvC�]�m�ދlw ��Jh8)�%�۸��g�L�Y�X�&��{������!%�g��� :��w�|;�ޘ#�{=p�qm�ܝ��6�~�����\�_%��DW�@Ś��=Jׂ""6�p����Q �����f�����V��	j�t~ոh;f�