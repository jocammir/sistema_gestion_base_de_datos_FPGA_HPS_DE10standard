��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��Nڭ�	�����B�#Z���?�4�j��0�ΐz�A�y�[��I4�fB���_Ɛ���-����B���M'~��k,���'zf���]A�� -̭���ҧ���D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T��P�]��h�� �x��ɻ/�akB�����L%��s�A�ۆ�)�a7�$�HID	���� ��Ѫ�2O�ұ-�(Y����a���D[9�.��:k=%WX�o�>�s���g�>��'�{�ܥ��3���0V���>�hV3]܋y���"�fD�����t�Q�k��p|�m� �2�{�!!M1g�b�þ����M���:�֘Kk�I������3.R�����W�����s,��W����rm	I��/���Q6�aźm�.}fEM��u2�rz�>���}���Q^�"�#�'��̤��`�}�Z�M�:@��,k�<�#�]��4=m'*~��3�V��j:d����������<��#i�)ZE_FZ�������fs��I
��ű��i��e$	��0��;�fb���z�����7��\��Z����v�,=Ţ5=��-�.�CRd��D���MlD%�p�J[�Mif��p9�څ�K�r�9lu��~iw�7��ٹH�4���]��$���[��7O�%ƕ�p��~3�tO�F��7��A���\O=G���F�E3�1���h���U�\�Y�.o����D��Am��^���j��h���8�������4��M���o�}!nK�z�(l�0����F��*���]W�H�d��uP3�KW���x.��Q���B������j�W� �PnW`U%�]J���ݤ�㎩!�kN�B��.���W��>$��ލ�v� �?���I��m��߬�J�"+�h�V&�1m�C��orP��#�����,�놈վν���5���2��3 �N�!��53s ���D�p���M9�%А|�L������n�Tz�M��]
Դe��j�`�i?���em+D��j���jTt�C8wMݨ[}�i�ț�q5"@��G�Ә(4����r}$b��$��b�Q)y42]���9XB�av���~��?9�!c���њ4�f"Z}G�c�$���/*e��i�f��op#P\B<����5�[ׁ��Z�7~����u�J囥��㥒;��~"���� <���{�p-B����h�9J�}#ieI�>5��+�S
^K���G*��኎x'��E�N=Q�6H�HL��^�%�UH����݅����(����3�z�����;�x�)�;�l��<�*��Y.����o�N�c)4dϻ�#Zή����`5(�~�xl7��_��)��;b�ދ�O �~�|k���4q�����@¿�y(�SD�y��/OZ�����>YJ#���ϛ�M,nhb[����bd�t�8��\vV�c�|�G���F��
�����y�/��	��r}� �lh�\�C�T�=c���ط��e�Cu.�� 8�p�`+���x�puG6s��f�?�g��GJ�V=/����Ċz��Q�0��\@�y�Tz�۶u��g=�⾄t9�Es>�w���6H�g�$K��<Eu�(�k�^ʝ�n�k��[`|m��0y�<'ؒƑO��\��RR�ĭU��F#]DF��ogTo��o��rzL+�a�����1����!�[�S�i�h���
ڶ(���`��.�u�4*��0�d1���Z� %Խ�<�~(\
�]ۼP�ґ�1��z��&���������R�`�@��5Z-���Yt�4:�u�Z�aN5l(S����=�*)J]��[A��MǝM&�㼐	Ʀ�\��Ұ�j��Ԋ�Q������3��4P�a�'�B���!n%�yh�8����?���3���`q���(�@f/L&���M(ٽ��SZV�=gQS��J��G���O�=��Y��q�G\F�MN��b���<P�/uR�L�9�g��ȕ�$h�����|A�#i�E��X�lp.-!c{�FP,g`�3	��"�ir7k��b�C�����c2'���/Kbt
�Q��=,��m%Ũ�E9E��Ty~�{�2�+� ���1�Gߐ���/y��E>}^����^�@��M�(Fhy��
��:s����N�jە�W�F�<�	��K%^� ;'̻��/_M��R�m�a��M��ί�2���Q�u�3u��������i�ъ| ��'��΁Fe��Hv��x�@UpNH��/ʇd�Q8��2Jǧ)aE��3lj����*���2��r��z�[����,<~F��� �NP��e�S�.N���R��?.:НF.��|ǣD_�'��}��dfԪr���=gN�l2c���q0��+Kw��w�=JowdG�l�M�[���2�{�sUv-��;TF������?�i���,�"����l��J�1�iCğ"�����ɦ/:De�Â=?�{ݰ��m�[�U�So(�&+��S��={�0wv��A�Z�q1���Z�����mӁ:Cm����{>ܲ���y���8Xi��<��1�1�|�#�kX�[�vlׇ�nåՌh?�
3	ɠ�L��G��A��~�"��Ɔmf�ޯ�� d����D�A2�t]�J��d�q�U�yzm/|�\J�l�O���NB��ٴ�s���W7����,��k�������O��;Ծ��_��Q�P�_��[n��X��������3m�صy���F��^I�Vպ죔��ي�i �B �[\��(�Jb%Q�N��^�S�_p�5z�r؃�y�v�ʏ�ߍ2p��!֛t����?S�#z2F�;e���$��/������*�vu���-�4;���Z�*6��_���2L�؃���dyhpI�N�����>nⅆ�2��`��l$���*�mZe��a�y�W=��XZ�=��oRFU.��m=;���^X���s\/֞Wr�&���Ba�%�doi'��s!Bp�Kv�(H(�&�	�i�����B4�~Z��d��I0�
�۰��
(�"��d|��3Yq"�!::`��(��Q,�t2:{\5��)�C�O��X����a#5ƻ�h�3�*����,�zM�OOq�3ZR�3NO�=z�6&�>�@P�j ˂��3��u2<�����[��-"U��@sYh�x9ND-�D�&��$��<�p3*�\w���)M��.���4��&�Η�-ՀJ��u��@�~B��"���#Vb�A>@K�=6��poucxǭMJ�����Q-gi���X���}�u W �u>�7|WCcvNq�ޓ5�m��e���x���!ߐ���&����ԥ��)/���s��
LE�##F@Ā��wD�v��K�~�#)l�釺ě+B\̮���K��x��cӥ_5�(�r>*^-� �,B��o �9��bذ�q�|T�9���ZhhxT��Z��1+gf�Ź�2�BD(k�!;t���l�yiF�ұD��%)z�;<��0eݣy�&L;>-O�7�c@�L߮Bv䮌����ì�C*��{@%7�1'�R����j�ۇyd��@�ۺ���������!m��vsx���(��l�Q���m)��O�M�V?잴��Mzt�]%����9���D� ����P�A��$r��	��0�
���,�9�L�uJ��,��d6ZS��⯔0U���te=��ɞU�m~�2λ]ݍ)��G�yX)���p�>��ϏR�*�X�O4�eQ�;=ӧ(P�����8:��E_Y��j��85��v��{�P�F�t*�������=),�CJ�DI
d��=����`�L%C۠03=�ƍ�(ͼ@���+�y�P�5ډr
1�܊���E:y�ŀue�g�ğf��'����!��RЕHR�vT�	>����$|w/&%]v\K�.,�T�C.�X]��"�|aO>�:��4DүƅH�rщ���=H��D����}I{܄vE����
��"���@�W6�w��x�e����'�@�퉋���poP�y�Q{(C9�:�� f����]�	V?)ߠ7�Y�ĥ�LB/�؟!���z-��X�9#��������Q29�=1;J�Q*�SV�2+;	ʰ�#��6�M	��M�5�L�R���ѨJ��.�1�>����:csr;���Dm���*uI�k��6����?<�x�s8�Å�C7��+�?Ŭ;��2b�k�l��Y[:O�~���J?���.B�$�c\E(���C܁���*$+}�Lq"=G�M�R���|�����xIj�]��fHz��$(�+�i�T��'����"4wx�R�S۞"�({��<�9y��H��oA�Ku"��4Rk�]�A��I+�}0F����!�9�+��r1�p�ƀ� 3�k�V���|�+pv\r{��M��$A�{��]��ߟ�,ԧ�[���4\��ڤ�C5Tjɡ�����$8��	��n����%'�2	k���aw����%��I�V�����q����10���O��i�g2��W�v��Hx�]���B�ᄛ݅֌��̷	����C��k4�v
`t�>p[OK? �9eM�'W�-�[qђ�}>��EdL&��e�ɗL!8x"b��Pҕ��"�>���s�-+����9��L�=��*�gd�z�i��_Q�E[o�r:"�b	eK �p�Kb���^A6N��XǺS�:@����x��?�%X�*Q<��M� .��� �8��4��6e�{-����n�g�t�*��M{4�8�A�:�8�e�����H&����ֈ]I�<��2��*��*X�m�g��c��્:����	��RW)$���Y9�="Ch�Elf�(@`S/"n�. ؜,򂇒�`&vf?n�
D׌IXjj��,��A��r��5U�6��a���s�����N>\D߿�N�j��v�Nvn������=�]�#R'��<��Z1yd������i�-ءC��uù�d�Ls�$g���믹�澾"T��~�T�,��C��aƅ�${+�dZY�W��~c����܎���Ԫ ���o�ܬ[�Y�ݸ�LL��h[�Ü��ٗJ�����S��"�S�ףn�*��������"�>���;�^;�#jg �ϣ���[&1��GhX�,%�L(@cR�T-ÈC�sl�̍H; �O3�&�p�%f�����A2ڏ,�5�K��`˞������gBS�7<7��B��H�cj����S��a������AJ��U!~�%����9��t˼o�w���a�y��g�"C
2�������t�`��d� O��������{��0�����ˍ(�$!�z'+[�c�����5�C�!q�-P��<% � S�8�TI6ya6-��vn6_�I�=`�_�Ē��W(�	�jI�WL,D��g�8cb��k�F�j��x{�<�x]��K���Ơ�������{a��q�٬qR����U�����Z);q�ZSuZ����|j8�o|5-b�$�\�w�Ql�4��
to�QN��v� ��P|vC�\�xmm�-uI��Wǀw4�.�PO~�K8�]� O-ݽ��4R��b��p>)����Ty���χɍ�gr�	�	3�9� o����"��
@�Zr�!�$���|���r;�q���if2����j�T-��B�V�ka<�-�;11o�f�9�kγm@���$�ƚ"Z5��PX�<��`kG���ݷ�h ��pH���,'���?ֹ� �{3IL2�ƻEڋ3�QgYz6չ�HO�ƶ���ߕ'1��e^&q�P 2��)���\5�SF����֜�5��K���#��J /�`����R;�p//>��G��Qu�{�V�����P7��H��l�QF���[����O��������,OcIi�����{L�=�|Z���=a��Ɯ�9~V΃(eM�y��R�b�����dCt����6t>�z|�n]팋[u%���4�VXr*��Q�
�g1�q
�Jv���� ���3���\��w���(���CQ��.	@���[=d�{1�*�px��K�E�����m���T[x�=Z+ΐ�������~��rՒ9E~:���=�xNV��x�h o�����~w�N��7	�<�?(ohxV�����Z�_
$t�����X�4��b)�YmC_��눗��������1` w����E� -�2��N������Ԟ���T����P��-zg�t��V��j���(�jP�T�&���mwx�@�aul8��rF�$�[%O�̠�-]O�1}.a.r��cp� s��Uӑ��#��@C�4�p<B�k�ٰ�#�+����ti�){�;x�z����3*�;���[����#RgTX^N�5��9h�3���|I�E���fO��3��"}����<�h�-
!��:�Jz�Wfz*����N��J*�� ����!	1�w�Mi�	�?�����.����֖/e?���7�G}uw�<��u�#I�䣳��k�O�K���劝��Rv���i`66�����vY2�)�0�:�%��@=�NU�ȯ�)sn�dW�+�F�I�5�D�����k�w��eD���s�/|G�ڮ�G6��1������dr�u7��|/Ri����$��`�ᥤ���?'!��+�|�W)Xp��Y>��
���5�81�\�H �g�9��9.��G�	d3�x��_�5���p:)�>52��	?X�[���`��"���(�J������j}�D<������Q$`��D�y��?��l5�,ɳtV��}Væ�a�ݵ��Fp�^;�3���vݎ��}�	�d��)
@�����J��;�ۡS������36݊�8��w�cTt%��-�z�d*A��x��g��\��n�W��ɓ��5�]��K���@�=� -���{Jϰ&2�7��3�,�49:{��:b����7ףi�N���\�p�_�z��a`�͞� 
�������?�i,B4��Q�@E��f?/ȬDs4l
����L7ݻ�wR���pc���*��Y1|����kf��as`&�*��v����ei�FC4�!k���q�_gM�K+�?
���� Z��X(SϢ>��.�Wo�"E`�;���-B1;����W�� .��h��۲a�FF��HT3�� ��BO�����m��Z_ʈ��/O��"��ʍ5�J9u{r�<��I�k�ӭ4��6�Wt�J������ss���J��Ӳ���x-y_~��q�D���7�^?�uU�a�A���v���vU��mS�MT�>����&��W�e{zm{4���0	��=ҫp�W� R��KKPUw�&yj��JRt=qCҷG����M�C/�L#&OBط�;<v��PN�i�גt���w��FDn�e��$��@\R��!&�sӻr ��8���_��p9 ���#�N���-�,��z߫��
���cS��Tc��a��Yk��c�N��r���F�k[ i&��^_��W��()QxO��~Ch��O�?�і�~�	��<����*"�e-�!��$��a1T
n�g�$w�1=-�ez�J��q�+�����������Y��K?��;�ALV���i� DY�^��I��<㫃�`���16@��2K�;�� ���K7) �3���Щ2��� N__gK�0{�����je� ��I��څz8���L���n!׌e�*q�-q��M�j�H�4:�Z{�̙��t��C~��Ƥej%@U�<=��oR���(Hh����g�p;f=c�<J�E��7�FM�c�����QL�.վ*�ƞ�݂o��!��f����X��єp��,n<!���~�C3)h8'����q�mo��g�h A����3c�,�sO�iM��;,B�hFD�!D5�/�ێ0�����S�5�hO$}�
��y� >�ċv��6ec�k�6n[d�A|�Ā�i���p��I$ѢۆD���a��u�eU�=?��SP��޼��w��"�^?�6v �Ƕ�ė4���4+����9���o�@�p��6L�2Lо�p����7���ޞ ��@TH��h���l��� u������K1�Zp�18���I���B{1R~��2���1�Gܩ�Cm���,�T�7��vZߓS�Ó�Č���Md���6���G������DTLg�	!�σN`�iZ)h�<��GUM��rL���9	�b�Z��r���`�Sӽ}s	r�N���i�������.,�4��`�i��
4�P��h �i̮0!�Wa�ܚA�l=:Lzb���j�m��J���X���p�yH�v�¢d��ж�������X���y׌�n�����rɬ��-�w�Ǡ0��顄��W�/���'2ӫ!��Q�u��|)t���������o)������ؕc��9��&�]$	�@��t'%3(����>{e��qW��<�/�}��c�L����җ
� �ՇN�_=�8�J�bx�v�ϗSqc��Ξ�e��6��\�ա���}x�'������s�c�~^A��$H:��i���X�^�m��� ���-Y�,nR�~O����?�F�LW��&��Gg��{����QH�Lԙ��zv��p8)wc$��k^y�#͊s?�^ Ⱐ�����TI���p���b��t���q�"*�F�v�H��3��r3$1��s��v�~��Qܥ�x�F��	�=�]^j���gupi@2�93Rr7��c�M ���G��Y\b�䮖:HDC�#�� Yo��n�Og<X��]	��viE���lo�[�hf��3�d�sMV+�Xr?�Jk��B�s�� �c�F�.G�ۜ����B�!	����mh�efͿ����|�[�o�|�:c��6�t�P�Q5H�:��ET*z,g0���]Ӊ�$$�t�=NĲ��d��+�(ŵ?�͈���0��yV���Yp�-?t��]�O��������h�d�B��vfIIc��5��h��:nu Q=����/<X�F�a�L��'��x*@f�_�
��p.�B�P0t]H���*�F�򘔵s�����9�x��ӫF�?�u���z�ı�������))ٯ���bN����?u	
C�p����I�F�3}�d�x���0�jT�3ʮ�;�Z)K�z�� ��x�$�b�<��ɸ����𘗓�Sd�����Sh�?��|�czj�?���	�U>�4M����#T��yu�ֲ�ǚx/'�r5��M=0��*SQ�Wf(\�78GMUˡ�<˧��~K��Pyo"���Z3�v�s6!-{3�R%MЁe~��e�8"�H�'���g��-:��6�
[/��{̐=��5d�Ν*7Bi0�/��"H�qzs߅�O��&¬ô����
D�q���HD��|�]2%��[r�"�"��k5�VT����?�t"z&����f��ql���}
%���z�G�9 ;Z�JAG�w���붸�_p���E�ޛ�FL�۴*wv짐w�v��z���b�X%�SVt�����Ԋ�z>��4$��=����*Ja ���ǓUi�P�L�(�:
�%�]���;Ax��\�<(g���N�U�b#i�NT������H�QA����|���e���8P������״��A��D��WT�Nɳ�ޙqQ�Ը��i�c���Ч@6����KE}Aba�e�&O�W!�S3��v��U:� ��\���eZL����=��/Ĕ�P��.i�"�%Y&��W_x{;���d���i`��������/X���v0��heS�lI��6�6��m$�A.P񘠱���Eɋ���{)쉗�/�_�މyJ�r�F�LNҨ+�� �(�ͺ�۟I���p�}&��G���[Ƴh��?�,�"�˘ϐ|��n�w��"w �KP�āT���*�nrɛ9����qҦQֿ_ʷP�:����G�K(�i�SJ{`�k����ụ(����u�D֡��'��vc8QE�|u*+�l����@�r����Ex8������0X����4Y|�v#��k���Ԥû�� q� ��p!<�`����P�°V�yw�p�8/m�y8�=���L��:����Z0��k�_�|D�b��|�i�$�>$�?���W���2T�V0yPC�Ua�&�i�$Js^n�1$+����V5-���}mjj�I��Ԯt�0Qv�w�	m%��e�>J��4�C5�M�Dn�:�V�7v����V��.����:-��_'j��.[�D�V:��C[R�j(&�L�A��r獊x��0�� ��,3`}�%6gj��Y�k%�Ϸ��`��30B-�U���g����� ��p��D#�k�g��Z6�;t��!�/D.��aa+;#��G�O�%`����g}=��`f��;�
Х��!���~��|]#'$}�b��Xg�u��?J�K��,��u�I'z��`J��j�&C�X�+�<��d�LM�=���۷����k�πTq�z*xw�t��+��֑�y U�]^C�0��~���jJL�������s3��`�n|}�h��LE��:���SF� �I��bJ�r�1iN���j]}�����Dr� U��jwb�R�rU�B�[��tJM1,��-�YW|��WG�zg�y;��&S�*y�W��L���d��U���Ts�*JW���Ȉ���i�/�O���3N�S��R/Q���qK�����TJ*�w�p����$��ˬ=������UN(��1~�lpZ�HSu�ê�_ �I�̼�u�್d�h��9�<����Q uz�y��.��Q�4��KG`�������TB��5`г�yrm9��!�=~��Dx]q[sbn�,��O5t��zĄ����MB�5jN ����Pl������U"uȻ�t[7�Aw���8�$|b��_�)�M�Xd�sm��y>���}���Ź��jd������c�����i) 
Լp�k_�d��`D1o>���۠�uw�ھ�W�QΧ��abEIԇ�cs[�CVv����]��
�% �M7��Y	r'���u��5]w`XZ��d�ѹ%:��bu/��1��=W��apk���Q
�Q+o`ҩkٵe�>�V�C�=�l��QE�c�ˈ0I���Rf��mIv���
�������?��K2�9 ��'����.��yHi��a�1k[�ǅߘC�3���G	8Nkgon���+XN�S�,&->�����y&�E���9;ϤV��-��d#9]a#k���Lj�� 貸ʯI��R���Z�<�G�5�Y����|٪��?�A�h�p(�0�s������j�z��$Y�5�r�3A~G6s�j�Pѳ�tY�^?��Mv���{8n���,�,�R�z���=�g�L^�j�emTv5e���ѱ�$�oda��u?����rb,+ɈWR��q
�Mg^H��Lpl�e����ǔ�b�x�F��ű��<V[`��6�=f���?~�r���:`4�1p�3���ߦ� �q��vP���=��u�,`�V�f��+l������ȍqE�t���0��(߶�Y�6mqWtZ mu$�i �U���Di��>���LD))kT�c<�J��p�1r'�?�����#�D c�"�Y�u`�9峑��㵰���;A�,�S���y8����z�\� ����z��&�ݔH��+�-�{{4��(�v��娄�IxB��Ǯ��%X5��yr�^��\^x���,�����	����I�.a�� ��	tu���>i��,���H!8]-AEͺV0��^[c�A��Z]Q~L2*�I�IE���E!Pŋ�
@N�M�k�Ş�����]�=��AK�7mx̍
hZ+���ѡ3j�'���b�`i
ݦA�7���4O4�o3��?��S�P��R����]���k܎��.z(YY�79%-�dԷ�k�uL���Dg�|�d$��w�I�$���)sC�\���~��M�#Ȁ�%Z� ?�뱀�X�+q�E�G�*_oP���[�w`Cg�J����J��Д!�ǜ8˚�Jz;|�o@�]���n�ҿ�u�D�ƽL� �c�ܐ���E��sx�D�S9Q8���s|^�3�}�N���2����L$�|�Eb{�-�������Q��Q��F����>$�0<]Es|�j5Кh��:o0(r��xVc�`\��z1F�������Fu �t�_f8��k�~O�*��df(�]S����#�.��Û� #�)vY3�S����(�-����m��ܢ�j�삔]��+�%�����c�j��b<SȜJ?��/,g���nd�z"����i W�⎽�_:������/��kﻷ�����$�G��^,P�u|Px�H�7�I���Mc���12	�j���|L��W�"���z��'�G�2��M���N�e�aF�R�ݩ��_� ���͟�	��*8J>6N��Z�����m"ݢ��5,S�Iqp�i}����r�L���Ty�`p��e|�=|�]#&.��'�-E*������~�J�}��S�O� b�l�=���i��S��-��rat�k�n�_Ȟ�r4�A �g���a�#�O��*�1��-�cO'!�S٥�����J�i>��/O�C6�ݎc1*tC11�(M�(TS�-��ت84��Fy�2��ܐ��� �=��ڈn��gb��#��%���6DN�ϜO��d�m�N�%��Ƕ�����	]ڶ�]Q��<����Z#�xs���$�s<y�](s)��/]�g�=1�iZ�)k
�Y��7�3p��.r[�n��G�h�)R#�(.5�B� qi��%DA�ষy6@+�b���$d!��&�ػS����f���́�I�R��zx���%�ߜ�)�*3q =��5�
u�=ݡ<!�^�Ց������=m�z�پ-sĜb���9�P+*Ze��Yo%�r�ZJ�ma���"H�@Zl�0����ʑi՞	����g@��bE/l�@����&A\���{7f+�M���Jg-HU#S`Ű�즬��dp�*:%�Ґ*���7Y�'�2�<}�������V��ڷÄΓ�/0r�J�6,�FB�
?0w�yI��J�&U%��E3Ң���P>f�sȢv��QQ*�" A��-��Ti��~v���l�����{��n�BU,c��,Y����tG�7��`�����-�"�B���ʥ���Q����b�~������YR=,��z\'*����+��TEQJ���f�z���yE��?���r�;��قؼ�<�յ���8�$���_p�>��{��I��T��a��"rj#d#���&�8�o��!� L��sRzǬYD���<�&P��y�$��ؕ=�7��).�Ӷp�ω��P��ǳ��x+���vCd�	7^{ɭm�4+�Es�B�o�+�%�l�ol?���+�H�������.�Ѷ���N�`Ζb	�|�$�u�k��Z7�/�t�ޓ
��2h��A�l�H������o��O&�&�rG�ø�x����϶��K��j�<]y�"Gu�1��{�$,�s��Y2�.��w`�/dG��<O�i&!#m�Qb��8��Xl�mF|:>DL�a�d�[]������	tQ21��Y]�;W�9�/!}6.��;�QJ��|��.���`��X�X���般������\y�A"��������DcT�iM��#Ѻu۞D>d���N$��u����\ą����"��.��%&@�@�M@9cg�Y�~!�9J���rHA�b�=�&I��H��6V��s�j�O 8�.��	�� 0w��1WK�@c̽��`;p��r,�x�5�Gq�t�~5饲�H�����W�B��a�Ȁ�
��d�X���*���R��K�/2�g��8AY����a�D�����*�g/�C�������~uH틿���t���b^��k�����=���8��H�N�C)໫�kF���I��h��	]j4��T�˙��8��@W�:C��}1yC�����]�`�����r &���(.���c c>$����n��`$,����8�H�I[�.�7��`z�I8pR]��i�$� ���?��u��س�+n9z[JF4�4m98�eW�ā�^S�֒��$�ϱZ��iC��Ӛ�-�akS$//Y��G4Sio�uZ���\��{e�Q"=T&~Mf+k�@�We����>��!�օ7�*f����C3&a�b�u�<X�OН\�5�>�t����鄠]<��M�@�3'?|QX9���T��0��$_ ���´���[3>5cZ�;�	@:.k�qe<"�V3j���,fZ��`��Hb�ƕ���l������������F�	+���%�B?|��&��u�\�">���`����W5��1�Q���G�hږ)��?�\(�ˮ,�2v8��`��uν���)��aen���]кq�s�rG[(�+�����zʏ�-a`{�e0k��yK�����9T)mK�����$�N��Ƽ�s�1$�cb	�{��l�2�d@�A�J	�>�\Nyؘ��S}%�G���P�1�0v�V5)*�j�Sa>�w�� 6�LiYݞ`����7�B�8���D)+��s�Xm�����H�9�
��v��P�|q����K-�����R�Nf:-�X�m?�N��5�^�]��d�o�F�l=��ncw���o˫���� ��fb�\�kVy���JiR�曔����+tP>q/����e�JV$�1��������=����=M�h�66Fӵ��Sx�ePL5�)P+������U�1�@\���f)�l�o3�^Ʋy�K~s�
�&2J��т<N�.�7�<�b���Wo�0[��D���I]��O^eղ�i�)�@�˔I�����8oYx�s�F�[�,֔]?���J��ܴ�1a�N�a����1�p��Z����0����������;�I�S��B̨�LR@F�s�II#���)��'K�+]�؜�WF~1��̜O&#��:���V&P]1��gm3��K�۽��"��/Q "��M���$7y���{o;�iw��!V$�3B-�����+�dMX#�9�V��O� M�-�s(���V��Au�~�g�VG��x��/+S�ď-؋MU���y�H���!�<ᶃb1䍩�(:��f������T �Ca5��ƹv�Tt��%~\j)�.��]Rz�g9I��c����r�N�KgP��ß)�v��<�K|_��ε`��|nQ���e��ı�K�� ��]�`Q!��W��[�e�6��oc������nGJ�����t%�)�4E\P�" r���B�)�3m��JbQC����-�x
jaZg�8�����%�`f��b7�:��MF�����3��.�jB+��ʴ�j��4:�i��|�l̻
�����JB�ԣl<@F-��#�2�����|ǭ��3�/�߶��<����&�:��ĕܒ�Ӵ`��/z>��y0�y���GTDB)ڕ��A�l��i�l��