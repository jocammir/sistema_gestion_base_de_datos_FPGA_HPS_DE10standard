��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�G��?M`^ NmK0���C	�i��E��t= �5������1�m"N�I<�<�*�	FW���O��H�S�E����ߴ���oo1� 2��I�U�Ź�暰��	������S�U�I�����S�,��o~���G{xG�` �B��=��5M�7����~�Q�s��n���OJ8?pZG\
g,���P̐�tb���}�7L�,X
��?᫺D
����o�,矔����H��A�#�d}��k�7}�%��ƃ�\��4���R�^$H��-e&#�K?6�^��x)	]s�O��3
�+9�qWs�@ ��PV4��@�.�.R�����>�=�Y%=Ă?�W���@�-���N�7�-����U�K���W2�y��c�}r�%��GQ�]k��1�j��ǿsL�y�c���n��D��H&���uf����l�+a[���f럃�t��E
pd���w46,��N��R��sD!3�W���W�K��u����٨�;�?�߽hi&V�yE�π���`Q�a�b c�/r��=��I��
��Nd!r L�h�#����B�㾍-�ɠO�`��..h�ѽ���)��P)?gU�`?0�_�J���r<H���u�1?5���|7�8\i�q��Q/���e���ǭ�'��V�u�r���Rɫ�*E�o�d�&� g�cb5�Q�/Ǳ��{ط*�_Q.◢H=�*K�x�弹=��E����6~����:�ם!=2�	�x:�ȢN�:��fi��*k��M���8�%�s���[��.	KqQ+��C���J}X�	���p�b��S�	X/�^*�bJY��^��*��Ax��pmE�ؑ�����	{�̀+�ǵ#U�MT��}�i��}�
�����N8���cXw]H98�S�	� �/�'��O�ޮ�a^�����b�\i�\ �2_�1�'�,0f��Vb7O�[�{�I�X�ɽ!��{Ω< *�	f!�U۰�{!��YI8�z�n	���.Џ!�Y���MG���$ �-�`0�	�'�����s���)'����Z1MW��[�VD���Q� �!�mO�T�Sn�K�~�>K#fb���Dh�R�!?&@��;BɆ^]�Z�y�128�Tِ�\���ֈ��3"�w��J40��43>AҲp���3L��F��h	e9W3T��D��?�x=�����/��5���C�l]��<ܫ��潍Z��£�/��|r��D���CS���۟�XV<+��R/���sk� ���Q�
/��q,�� ��^��ei�[�{%�nZ3����T1Xx*V�8|�%�_y��3_�4ee�uͽ~3�$���[��2����e����*B����ЅR�rc�O9��}�e�՗��;���s�W�t�?���l��5��I�i�k��v�#&˫��>�z78ˆ<�	k��y��c�e�a��Zs.���We�]Q��'�K�����@��DBη(STx�DJ�>�g��6g̽���:��d��q:��).�E%(�̮`�"�ƻq�9�&���Z[c;sU��=���]�T��N�?a�*K�v��x��U� ����6�L?t|S!�gF�K�|��us厀��s�$�L�B?�'�/�`�e9}(�@�cU>V���o����~9<c�SJ�O͇���r,�������/��$͈�0R���:;����K)�/�|���%�+~/��l�>%�n��E�@m�e��&���h�3\����:�L�8G.��W�O�٣{t�oo#(oDb~�}>�ɏ,E�&��@��p�f�H.0�[�Em�b# �~�x7� ᗶ��?�o��nd�6�����b���?������gg������^��ȵ�ϳt=2�Q�a�Y�MΠ�K��S��Y�r�(=�uh3��V-M�K�B�_��mV����+�A��#�dѣH�	��uƂ	�Ui��p}��`�"�@l�9�"k�ne* RO5�{kMt�:s*�-y��I���A�er��}���?�{K#U:���6���=�}֍��K���ڲ�!�Ḵ{C�%3����Il�K�����[$P
�Ҕ�-����޽{��2k�o�9<����s<���-_�]�lS/���Ē�ɖ6lЫV���.�C�X]�D��-�ch3���ʪ����I